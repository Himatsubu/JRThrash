/*
TimeStamp:	2017/1/18		15:13
*/


module subunder(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy,	
	input  signed  [13:0] i_fld_u_0_addr_0,	
	input          [31:0] i_fld_u_0_datain_0,	
	output         [31:0] o_fld_u_0_dataout_0,	
	input                 i_fld_u_0_r_w_0,	
	input  signed  [13:0] i_fld_result_1_addr_0,	
	input          [31:0] i_fld_result_1_datain_0,	
	output         [31:0] o_fld_result_1_dataout_0,	
	input                 i_fld_result_1_r_w_0,

	//ここから追加部分
	//under2up
	output         [31:0] r_ip_fifo_under2up_in_0,
	output         [31:0] r_ip_fifo_under2up_s_we_0,
	output         [31:0] r_ip_fifo_under2up_s_re_0,
	input          [31:0] w_ip_fifo_under2up_resut_0,

	//up2under
	output         [31:0] r_ip_fifo_up2under_in_0,
	output         [31:0] r_ip_fifo_up2under_s_we_0,
	output         [31:0] r_ip_fifo_up2under_s_re_0,
	input          [31:0] w_ip_fifo_up2under_result_0
		
);

	reg         [31:0] r_ip_AddFloat_portA_0;
	reg         [31:0] r_ip_AddFloat_portB_0;
	wire        [31:0] w_ip_AddFloat_result_0;
	reg         [31:0] r_ip_MultFloat_multiplicand_0;
	reg         [31:0] r_ip_MultFloat_multiplier_0;
	wire        [31:0] w_ip_MultFloat_product_0;
	reg  signed [31:0] r_ip_FixedToFloat_fixed_0;
	wire        [31:0] w_ip_FixedToFloat_floating_0;
	reg         [31:0] r_ip_fifo_under2up_in_0;
	reg  signed [31:0] r_ip_fifo_under2up_s_we_0;
	reg  signed [31:0] r_ip_fifo_under2up_s_re_0;
	wire        [31:0] w_ip_fifo_under2up_result_0;
	reg                r_ip_fifo_under2up_newData_0;
	reg         [31:0] r_ip_fifo_up2under_in_0;
	reg  signed [31:0] r_ip_fifo_up2under_s_we_0;
	reg  signed [31:0] r_ip_fifo_up2under_s_re_0;
	wire        [31:0] w_ip_fifo_up2under_result_0;
	reg                r_ip_fifo_up2under_newData_0;
	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 5:0] r_sys_run_phase;
	reg         [ 1:0] r_sys_run_stage;
	reg         [ 8:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 1:0] w_sys_run_stage_p1;
	wire        [ 8:0] w_sys_run_step_p1;
	wire signed [13:0] w_fld_u_0_addr_0;
	wire        [31:0] w_fld_u_0_datain_0;
	wire        [31:0] w_fld_u_0_dataout_0;
	wire               w_fld_u_0_r_w_0;
	wire               w_fld_u_0_ce_0;
	reg  signed [13:0] r_fld_u_0_addr_1;
	reg         [31:0] r_fld_u_0_datain_1;
	wire        [31:0] w_fld_u_0_dataout_1;
	reg                r_fld_u_0_r_w_1;
	wire               w_fld_u_0_ce_1;
	wire signed [13:0] w_fld_result_1_addr_0;
	wire        [31:0] w_fld_result_1_datain_0;
	wire        [31:0] w_fld_result_1_dataout_0;
	wire               w_fld_result_1_r_w_0;
	wire               w_fld_result_1_ce_0;
	reg  signed [13:0] r_fld_result_1_addr_1;
	reg         [31:0] r_fld_result_1_datain_1;
	wire        [31:0] w_fld_result_1_dataout_1;
	reg                r_fld_result_1_r_w_1;
	wire               w_fld_result_1_ce_1;
	reg         [31:0] r_fld_r1_2;
	reg         [31:0] r_fld_r2_3;
	reg         [31:0] r_fld_dx_4;
	reg         [31:0] r_fld_dy_5;
	reg         [31:0] r_fld_dt_6;
	reg  signed [31:0] r_run_k_7;
	reg  signed [31:0] r_run_j_8;
	reg  signed [31:0] r_run_s_under2up_re_9;
	reg  signed [31:0] r_run_s_under2up_we_10;
	reg  signed [31:0] r_run_s_up2under_re_11;
	reg  signed [31:0] r_run_s_up2under_we_12;
	reg  signed [31:0] r_run_copy0_j_19;
	reg  signed [31:0] r_run_copy1_j_20;
	reg  signed [31:0] r_run_copy2_j_21;
	reg  signed [31:0] r_run_copy3_j_22;
	reg  signed [31:0] r_run_copy4_j_23;
	reg  signed [31:0] r_run_copy5_j_24;
	reg  signed [31:0] r_run_copy6_j_25;
	reg  signed [31:0] r_run_copy7_j_26;
	reg  signed [31:0] r_run_copy0_j_27;
	reg  signed [31:0] r_sys_tmp0_int;
	reg  signed [31:0] r_sys_tmp1_int;
	reg  signed [31:0] r_sys_tmp2_int;
	reg  signed [31:0] r_sys_tmp3_int;
	reg  signed [31:0] r_sys_tmp4_int;
	reg  signed [31:0] r_sys_tmp5_int;
	reg  signed [31:0] r_sys_tmp6_int;
	reg  signed [31:0] r_sys_tmp7_int;
	reg  signed [31:0] r_sys_tmp8_int;
	reg  signed [31:0] r_sys_tmp9_int;
	reg  signed [31:0] r_sys_tmp10_int;
	reg  signed [31:0] r_sys_tmp11_int;
	reg  signed [31:0] r_sys_tmp12_int;
	reg  signed [31:0] r_sys_tmp13_int;
	reg  signed [31:0] r_sys_tmp14_int;
	reg  signed [31:0] r_sys_tmp15_int;
	reg  signed [31:0] r_sys_tmp16_int;
	reg  signed [31:0] r_sys_tmp17_int;
	reg  signed [31:0] r_sys_tmp18_int;
	reg  signed [31:0] r_sys_tmp19_int;
	reg  signed [31:0] r_sys_tmp20_int;
	reg  signed [31:0] r_sys_tmp21_int;
	reg  signed [31:0] r_sys_tmp22_int;
	reg  signed [31:0] r_sys_tmp23_int;
	reg  signed [31:0] r_sys_tmp24_int;
	reg  signed [31:0] r_sys_tmp25_int;
	reg  signed [31:0] r_sys_tmp26_int;
	reg  signed [31:0] r_sys_tmp27_int;
	reg  signed [31:0] r_sys_tmp28_int;
	reg  signed [31:0] r_sys_tmp29_int;
	reg  signed [31:0] r_sys_tmp30_int;
	reg  signed [31:0] r_sys_tmp31_int;
	reg  signed [31:0] r_sys_tmp32_int;
	reg  signed [31:0] r_sys_tmp33_int;
	reg  signed [31:0] r_sys_tmp34_int;
	reg  signed [31:0] r_sys_tmp35_int;
	reg  signed [31:0] r_sys_tmp36_int;
	reg  signed [31:0] r_sys_tmp37_int;
	reg  signed [31:0] r_sys_tmp38_int;
	reg  signed [31:0] r_sys_tmp39_int;
	reg  signed [31:0] r_sys_tmp40_int;
	reg  signed [31:0] r_sys_tmp41_int;
	reg  signed [31:0] r_sys_tmp42_int;
	reg  signed [31:0] r_sys_tmp43_int;
	reg  signed [31:0] r_sys_tmp44_int;
	reg  signed [31:0] r_sys_tmp45_int;
	reg  signed [31:0] r_sys_tmp46_int;
	reg  signed [31:0] r_sys_tmp47_int;
	reg  signed [31:0] r_sys_tmp48_int;
	reg  signed [31:0] r_sys_tmp49_int;
	reg  signed [31:0] r_sys_tmp50_int;
	reg  signed [31:0] r_sys_tmp51_int;
	reg  signed [31:0] r_sys_tmp52_int;
	reg  signed [31:0] r_sys_tmp53_int;
	reg  signed [31:0] r_sys_tmp54_int;
	reg  signed [31:0] r_sys_tmp55_int;
	reg  signed [31:0] r_sys_tmp56_int;
	reg  signed [31:0] r_sys_tmp57_int;
	reg  signed [31:0] r_sys_tmp58_int;
	reg  signed [31:0] r_sys_tmp59_int;
	reg  signed [31:0] r_sys_tmp60_int;
	reg  signed [31:0] r_sys_tmp61_int;
	reg  signed [31:0] r_sys_tmp62_int;
	reg  signed [31:0] r_sys_tmp63_int;
	reg  signed [31:0] r_sys_tmp64_int;
	reg  signed [31:0] r_sys_tmp65_int;
	reg  signed [31:0] r_sys_tmp66_int;
	reg  signed [31:0] r_sys_tmp67_int;
	reg  signed [31:0] r_sys_tmp68_int;
	reg  signed [31:0] r_sys_tmp69_int;
	reg  signed [31:0] r_sys_tmp70_int;
	reg  signed [31:0] r_sys_tmp71_int;
	reg  signed [31:0] r_sys_tmp72_int;
	reg  signed [31:0] r_sys_tmp73_int;
	reg  signed [31:0] r_sys_tmp74_int;
	reg  signed [31:0] r_sys_tmp75_int;
	reg  signed [31:0] r_sys_tmp76_int;
	reg  signed [31:0] r_sys_tmp77_int;
	reg  signed [31:0] r_sys_tmp78_int;
	reg  signed [31:0] r_sys_tmp79_int;
	reg  signed [31:0] r_sys_tmp80_int;
	reg  signed [31:0] r_sys_tmp81_int;
	reg  signed [31:0] r_sys_tmp82_int;
	reg  signed [31:0] r_sys_tmp83_int;
	reg  signed [31:0] r_sys_tmp84_int;
	reg  signed [31:0] r_sys_tmp85_int;
	reg  signed [31:0] r_sys_tmp86_int;
	reg  signed [31:0] r_sys_tmp87_int;
	reg  signed [31:0] r_sys_tmp88_int;
	reg  signed [31:0] r_sys_tmp89_int;
	reg  signed [31:0] r_sys_tmp90_int;
	reg  signed [31:0] r_sys_tmp91_int;
	reg  signed [31:0] r_sys_tmp92_int;
	reg  signed [31:0] r_sys_tmp93_int;
	reg  signed [31:0] r_sys_tmp94_int;
	reg  signed [31:0] r_sys_tmp95_int;
	reg  signed [31:0] r_sys_tmp96_int;
	reg  signed [31:0] r_sys_tmp97_int;
	reg  signed [31:0] r_sys_tmp98_int;
	reg  signed [31:0] r_sys_tmp99_int;
	reg  signed [31:0] r_sys_tmp100_int;
	reg  signed [31:0] r_sys_tmp101_int;
	reg  signed [31:0] r_sys_tmp102_int;
	reg  signed [31:0] r_sys_tmp103_int;
	reg  signed [31:0] r_sys_tmp104_int;
	reg  signed [31:0] r_sys_tmp105_int;
	reg  signed [31:0] r_sys_tmp106_int;
	reg  signed [31:0] r_sys_tmp107_int;
	reg  signed [31:0] r_sys_tmp108_int;
	reg  signed [31:0] r_sys_tmp109_int;
	reg  signed [31:0] r_sys_tmp110_int;
	reg  signed [31:0] r_sys_tmp111_int;
	reg  signed [31:0] r_sys_tmp112_int;
	reg  signed [31:0] r_sys_tmp113_int;
	reg  signed [31:0] r_sys_tmp114_int;
	reg  signed [31:0] r_sys_tmp115_int;
	reg  signed [31:0] r_sys_tmp116_int;
	reg  signed [31:0] r_sys_tmp117_int;
	reg  signed [31:0] r_sys_tmp118_int;
	reg  signed [31:0] r_sys_tmp119_int;
	reg  signed [31:0] r_sys_tmp120_int;
	reg  signed [31:0] r_sys_tmp121_int;
	reg  signed [31:0] r_sys_tmp122_int;
	reg  signed [31:0] r_sys_tmp123_int;
	reg  signed [31:0] r_sys_tmp124_int;
	reg  signed [31:0] r_sys_tmp125_int;
	reg  signed [31:0] r_sys_tmp126_int;
	reg  signed [31:0] r_sys_tmp127_int;
	reg  signed [31:0] r_sys_tmp128_int;
	reg  signed [31:0] r_sys_tmp129_int;
	reg  signed [31:0] r_sys_tmp130_int;
	reg  signed [31:0] r_sys_tmp131_int;
	reg  signed [31:0] r_sys_tmp132_int;
	reg  signed [31:0] r_sys_tmp133_int;
	reg  signed [31:0] r_sys_tmp134_int;
	reg  signed [31:0] r_sys_tmp135_int;
	reg  signed [31:0] r_sys_tmp136_int;
	reg  signed [31:0] r_sys_tmp137_int;
	reg  signed [31:0] r_sys_tmp138_int;
	reg  signed [31:0] r_sys_tmp139_int;
	reg  signed [31:0] r_sys_tmp140_int;
	reg  signed [31:0] r_sys_tmp141_int;
	reg  signed [31:0] r_sys_tmp142_int;
	reg  signed [31:0] r_sys_tmp143_int;
	reg  signed [31:0] r_sys_tmp144_int;
	reg  signed [31:0] r_sys_tmp145_int;
	reg  signed [31:0] r_sys_tmp146_int;
	reg  signed [31:0] r_sys_tmp147_int;
	reg  signed [31:0] r_sys_tmp148_int;
	reg  signed [31:0] r_sys_tmp149_int;
	reg  signed [31:0] r_sys_tmp150_int;
	reg  signed [31:0] r_sys_tmp151_int;
	reg  signed [31:0] r_sys_tmp152_int;
	reg  signed [31:0] r_sys_tmp153_int;
	reg  signed [31:0] r_sys_tmp154_int;
	reg  signed [31:0] r_sys_tmp155_int;
	reg  signed [31:0] r_sys_tmp156_int;
	reg  signed [31:0] r_sys_tmp157_int;
	reg  signed [31:0] r_sys_tmp158_int;
	reg  signed [31:0] r_sys_tmp159_int;
	reg  signed [31:0] r_sys_tmp160_int;
	reg  signed [31:0] r_sys_tmp161_int;
	reg  signed [31:0] r_sys_tmp162_int;
	reg  signed [31:0] r_sys_tmp163_int;
	reg  signed [31:0] r_sys_tmp164_int;
	reg  signed [31:0] r_sys_tmp165_int;
	reg  signed [31:0] r_sys_tmp166_int;
	reg  signed [31:0] r_sys_tmp167_int;
	reg  signed [31:0] r_sys_tmp168_int;
	reg  signed [31:0] r_sys_tmp169_int;
	reg  signed [31:0] r_sys_tmp170_int;
	reg  signed [31:0] r_sys_tmp171_int;
	reg  signed [31:0] r_sys_tmp172_int;
	reg  signed [31:0] r_sys_tmp173_int;
	reg  signed [31:0] r_sys_tmp174_int;
	reg  signed [31:0] r_sys_tmp175_int;
	reg  signed [31:0] r_sys_tmp176_int;
	reg  signed [31:0] r_sys_tmp177_int;
	reg  signed [31:0] r_sys_tmp178_int;
	reg  signed [31:0] r_sys_tmp179_int;
	reg  signed [31:0] r_sys_tmp180_int;
	reg  signed [31:0] r_sys_tmp181_int;
	reg  signed [31:0] r_sys_tmp182_int;
	reg  signed [31:0] r_sys_tmp183_int;
	reg  signed [31:0] r_sys_tmp184_int;
	reg  signed [31:0] r_sys_tmp185_int;
	reg  signed [31:0] r_sys_tmp186_int;
	reg  signed [31:0] r_sys_tmp187_int;
	reg  signed [31:0] r_sys_tmp188_int;
	reg  signed [31:0] r_sys_tmp189_int;
	reg  signed [31:0] r_sys_tmp190_int;
	reg  signed [31:0] r_sys_tmp191_int;
	reg  signed [31:0] r_sys_tmp192_int;
	reg  signed [31:0] r_sys_tmp193_int;
	reg  signed [31:0] r_sys_tmp194_int;
	reg  signed [31:0] r_sys_tmp195_int;
	reg  signed [31:0] r_sys_tmp196_int;
	reg  signed [31:0] r_sys_tmp197_int;
	reg  signed [31:0] r_sys_tmp198_int;
	reg  signed [31:0] r_sys_tmp199_int;
	reg  signed [31:0] r_sys_tmp200_int;
	reg  signed [31:0] r_sys_tmp201_int;
	reg  signed [31:0] r_sys_tmp202_int;
	reg  signed [31:0] r_sys_tmp203_int;
	reg  signed [31:0] r_sys_tmp204_int;
	reg  signed [31:0] r_sys_tmp205_int;
	reg  signed [31:0] r_sys_tmp206_int;
	reg  signed [31:0] r_sys_tmp207_int;
	reg  signed [31:0] r_sys_tmp208_int;
	reg  signed [31:0] r_sys_tmp209_int;
	reg  signed [31:0] r_sys_tmp210_int;
	reg  signed [31:0] r_sys_tmp211_int;
	reg  signed [31:0] r_sys_tmp212_int;
	reg  signed [31:0] r_sys_tmp213_int;
	reg  signed [31:0] r_sys_tmp214_int;
	reg  signed [31:0] r_sys_tmp215_int;
	reg  signed [31:0] r_sys_tmp216_int;
	reg  signed [31:0] r_sys_tmp217_int;
	reg  signed [31:0] r_sys_tmp218_int;
	reg  signed [31:0] r_sys_tmp219_int;
	reg  signed [31:0] r_sys_tmp220_int;
	reg  signed [31:0] r_sys_tmp221_int;
	reg  signed [31:0] r_sys_tmp222_int;
	reg  signed [31:0] r_sys_tmp223_int;
	reg  signed [31:0] r_sys_tmp224_int;
	reg  signed [31:0] r_sys_tmp225_int;
	reg  signed [31:0] r_sys_tmp226_int;
	reg  signed [31:0] r_sys_tmp227_int;
	reg  signed [31:0] r_sys_tmp228_int;
	reg  signed [31:0] r_sys_tmp229_int;
	reg  signed [31:0] r_sys_tmp230_int;
	reg  signed [31:0] r_sys_tmp231_int;
	reg  signed [31:0] r_sys_tmp232_int;
	reg  signed [31:0] r_sys_tmp233_int;
	reg  signed [31:0] r_sys_tmp234_int;
	reg  signed [31:0] r_sys_tmp235_int;
	reg  signed [31:0] r_sys_tmp236_int;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg         [31:0] r_sys_tmp4_float;
	reg         [31:0] r_sys_tmp5_float;
	reg         [31:0] r_sys_tmp6_float;
	reg         [31:0] r_sys_tmp7_float;
	reg         [31:0] r_sys_tmp8_float;
	reg         [31:0] r_sys_tmp9_float;
	reg         [31:0] r_sys_tmp10_float;
	reg         [31:0] r_sys_tmp11_float;
	reg         [31:0] r_sys_tmp12_float;
	reg         [31:0] r_sys_tmp13_float;
	reg         [31:0] r_sys_tmp14_float;
	reg         [31:0] r_sys_tmp15_float;
	reg         [31:0] r_sys_tmp16_float;
	reg         [31:0] r_sys_tmp17_float;
	reg         [31:0] r_sys_tmp18_float;
	reg         [31:0] r_sys_tmp19_float;
	reg         [31:0] r_sys_tmp20_float;
	reg         [31:0] r_sys_tmp21_float;
	reg         [31:0] r_sys_tmp22_float;
	reg         [31:0] r_sys_tmp23_float;
	reg         [31:0] r_sys_tmp24_float;
	reg         [31:0] r_sys_tmp25_float;
	reg         [31:0] r_sys_tmp26_float;
	reg         [31:0] r_sys_tmp27_float;
	reg         [31:0] r_sys_tmp28_float;
	reg         [31:0] r_sys_tmp29_float;
	reg         [31:0] r_sys_tmp30_float;
	reg         [31:0] r_sys_tmp31_float;
	reg         [31:0] r_sys_tmp32_float;
	reg         [31:0] r_sys_tmp33_float;
	reg         [31:0] r_sys_tmp34_float;
	reg         [31:0] r_sys_tmp35_float;
	reg         [31:0] r_sys_tmp36_float;
	reg         [31:0] r_sys_tmp37_float;
	reg         [31:0] r_sys_tmp38_float;
	reg         [31:0] r_sys_tmp39_float;
	reg         [31:0] r_sys_tmp40_float;
	reg         [31:0] r_sys_tmp41_float;
	reg         [31:0] r_sys_tmp42_float;
	reg         [31:0] r_sys_tmp43_float;
	reg         [31:0] r_sys_tmp44_float;
	reg         [31:0] r_sys_tmp45_float;
	reg         [31:0] r_sys_tmp46_float;
	reg         [31:0] r_sys_tmp47_float;
	reg         [31:0] r_sys_tmp48_float;
	reg         [31:0] r_sys_tmp49_float;
	reg         [31:0] r_sys_tmp50_float;
	reg         [31:0] r_sys_tmp51_float;
	reg         [31:0] r_sys_tmp52_float;
	reg         [31:0] r_sys_tmp53_float;
	reg         [31:0] r_sys_tmp54_float;
	reg         [31:0] r_sys_tmp55_float;
	reg         [31:0] r_sys_tmp56_float;
	reg         [31:0] r_sys_tmp57_float;
	reg         [31:0] r_sys_tmp58_float;
	reg         [31:0] r_sys_tmp59_float;
	reg         [31:0] r_sys_tmp60_float;
	reg         [31:0] r_sys_tmp61_float;
	reg         [31:0] r_sys_tmp62_float;
	reg         [31:0] r_sys_tmp63_float;
	reg         [31:0] r_sys_tmp64_float;
	reg         [31:0] r_sys_tmp65_float;
	reg         [31:0] r_sys_tmp66_float;
	reg         [31:0] r_sys_tmp67_float;
	reg         [31:0] r_sys_tmp68_float;
	reg         [31:0] r_sys_tmp69_float;
	reg         [31:0] r_sys_tmp70_float;
	reg         [31:0] r_sys_tmp71_float;
	reg         [31:0] r_sys_tmp72_float;
	reg         [31:0] r_sys_tmp73_float;
	reg         [31:0] r_sys_tmp74_float;
	reg         [31:0] r_sys_tmp75_float;
	reg         [31:0] r_sys_tmp76_float;
	reg         [31:0] r_sys_tmp77_float;
	reg         [31:0] r_sys_tmp78_float;
	reg         [31:0] r_sys_tmp79_float;
	reg         [31:0] r_sys_tmp80_float;
	reg         [31:0] r_sys_tmp81_float;
	reg         [31:0] r_sys_tmp82_float;
	reg         [31:0] r_sys_tmp83_float;
	reg         [31:0] r_sys_tmp84_float;
	reg         [31:0] r_sys_tmp85_float;
	reg         [31:0] r_sys_tmp86_float;
	reg         [31:0] r_sys_tmp87_float;
	reg         [31:0] r_sys_tmp88_float;
	reg         [31:0] r_sys_tmp89_float;
	reg         [31:0] r_sys_tmp90_float;
	reg         [31:0] r_sys_tmp91_float;
	reg         [31:0] r_sys_tmp92_float;
	reg         [31:0] r_sys_tmp93_float;
	reg         [31:0] r_sys_tmp94_float;
	reg         [31:0] r_sys_tmp95_float;
	reg         [31:0] r_sys_tmp96_float;
	reg         [31:0] r_sys_tmp97_float;
	wire        [31:0] w_sys_tmp1;
	wire        [31:0] w_sys_tmp3;
	wire        [31:0] w_sys_tmp4;
	wire signed [31:0] w_sys_tmp6;
	wire               w_sys_tmp7;
	wire               w_sys_tmp8;
	wire signed [31:0] w_sys_tmp9;
	wire signed [31:0] w_sys_tmp10;
	wire signed [31:0] w_sys_tmp11;
	wire               w_sys_tmp12;
	wire               w_sys_tmp13;
	wire signed [31:0] w_sys_tmp14;
	wire signed [31:0] w_sys_tmp17;
	wire signed [31:0] w_sys_tmp18;
	wire        [31:0] w_sys_tmp19;
	wire signed [31:0] w_sys_tmp20;
	wire signed [31:0] w_sys_tmp21;
	wire        [31:0] w_sys_tmp23;
	wire signed [31:0] w_sys_tmp25;
	wire signed [31:0] w_sys_tmp26;
	wire        [31:0] w_sys_tmp29;
	wire        [31:0] w_sys_tmp30;
	wire signed [31:0] w_sys_tmp31;
	wire signed [31:0] w_sys_tmp33;
	wire signed [31:0] w_sys_tmp34;
	wire signed [31:0] w_sys_tmp38;
	wire signed [31:0] w_sys_tmp39;
	wire signed [31:0] w_sys_tmp44;
	wire signed [31:0] w_sys_tmp46;
	wire signed [31:0] w_sys_tmp47;
	wire        [31:0] w_sys_tmp50;
	wire signed [31:0] w_sys_tmp51;
	wire signed [31:0] w_sys_tmp52;
	wire signed [31:0] w_sys_tmp53;
	wire signed [31:0] w_sys_tmp54;
	wire signed [31:0] w_sys_tmp55;
	wire signed [31:0] w_sys_tmp56;
	wire signed [31:0] w_sys_tmp57;
	wire signed [31:0] w_sys_tmp58;
	wire signed [31:0] w_sys_tmp59;
	wire signed [31:0] w_sys_tmp61;
	wire signed [31:0] w_sys_tmp62;
	wire signed [31:0] w_sys_tmp64;
	wire signed [31:0] w_sys_tmp65;
	wire signed [31:0] w_sys_tmp68;
	wire signed [31:0] w_sys_tmp69;
	wire signed [31:0] w_sys_tmp72;
	wire signed [31:0] w_sys_tmp73;
	wire signed [31:0] w_sys_tmp74;
	wire signed [31:0] w_sys_tmp79;
	wire signed [31:0] w_sys_tmp80;
	wire signed [31:0] w_sys_tmp82;
	wire signed [31:0] w_sys_tmp83;
	wire signed [31:0] w_sys_tmp84;
	wire signed [31:0] w_sys_tmp87;
	wire signed [31:0] w_sys_tmp88;
	wire signed [31:0] w_sys_tmp89;
	wire signed [31:0] w_sys_tmp94;
	wire signed [31:0] w_sys_tmp95;
	wire signed [31:0] w_sys_tmp97;
	wire signed [31:0] w_sys_tmp98;
	wire signed [31:0] w_sys_tmp99;
	wire signed [31:0] w_sys_tmp102;
	wire signed [31:0] w_sys_tmp1707;
	wire               w_sys_tmp1708;
	wire               w_sys_tmp1709;
	wire signed [31:0] w_sys_tmp1710;
	wire signed [31:0] w_sys_tmp1711;
	wire signed [31:0] w_sys_tmp1712;
	wire               w_sys_tmp1713;
	wire               w_sys_tmp1714;
	wire signed [31:0] w_sys_tmp1715;
	wire signed [31:0] w_sys_tmp1718;
	wire signed [31:0] w_sys_tmp1719;
	wire        [31:0] w_sys_tmp1720;
	wire signed [31:0] w_sys_tmp1721;
	wire signed [31:0] w_sys_tmp1722;
	wire signed [31:0] w_sys_tmp1724;
	wire signed [31:0] w_sys_tmp1725;
	wire signed [31:0] w_sys_tmp1727;
	wire signed [31:0] w_sys_tmp1728;
	wire signed [31:0] w_sys_tmp1731;
	wire signed [31:0] w_sys_tmp1732;
	wire               w_sys_tmp2036;
	wire signed [31:0] w_sys_tmp2037;
	wire        [31:0] w_sys_tmp2039;
	wire        [31:0] w_sys_tmp2040;
	wire signed [31:0] w_sys_tmp2041;
	wire signed [31:0] w_sys_tmp2042;
	wire signed [31:0] w_sys_tmp2043;
	wire               w_sys_tmp2044;
	wire signed [31:0] w_sys_tmp2045;
	wire signed [31:0] w_sys_tmp2048;
	wire        [31:0] w_sys_tmp2049;
	wire        [31:0] w_sys_tmp2050;
	wire signed [31:0] w_sys_tmp2051;
	wire        [31:0] w_sys_tmp2052;
	wire        [31:0] w_sys_tmp2053;
	wire        [31:0] w_sys_tmp2054;
	wire        [31:0] w_sys_tmp2055;
	wire        [31:0] w_sys_tmp2056;
	wire signed [31:0] w_sys_tmp2057;
	wire signed [31:0] w_sys_tmp2058;
	wire signed [31:0] w_sys_tmp2059;
	wire signed [31:0] w_sys_tmp2060;
	wire signed [31:0] w_sys_tmp2061;
	wire signed [31:0] w_sys_tmp2062;
	wire signed [31:0] w_sys_tmp2063;
	wire signed [31:0] w_sys_tmp2064;
	wire signed [31:0] w_sys_tmp2065;
	wire signed [31:0] w_sys_tmp2066;
	wire signed [31:0] w_sys_tmp2067;
	wire signed [31:0] w_sys_tmp2068;
	wire signed [31:0] w_sys_tmp2069;
	wire signed [31:0] w_sys_tmp2070;
	wire signed [31:0] w_sys_tmp2071;
	wire signed [31:0] w_sys_tmp2072;
	wire signed [31:0] w_sys_tmp2343;
	wire signed [31:0] w_sys_tmp2344;
	wire signed [31:0] w_sys_tmp2345;
	wire signed [31:0] w_sys_tmp2406;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 2'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 9'h1);
	assign o_fld_u_0_dataout_0 = w_fld_u_0_dataout_0;
	assign w_fld_u_0_addr_0 = i_fld_u_0_addr_0;
	assign w_fld_u_0_datain_0 = i_fld_u_0_datain_0;
	assign w_fld_u_0_r_w_0 = i_fld_u_0_r_w_0;
	assign w_fld_u_0_ce_0 = w_sys_ce;
	assign w_fld_u_0_ce_1 = w_sys_ce;
	assign o_fld_result_1_dataout_0 = w_fld_result_1_dataout_0;
	assign w_fld_result_1_addr_0 = i_fld_result_1_addr_0;
	assign w_fld_result_1_datain_0 = i_fld_result_1_datain_0;
	assign w_fld_result_1_r_w_0 = i_fld_result_1_r_w_0;
	assign w_fld_result_1_ce_0 = w_sys_ce;
	assign w_fld_result_1_ce_1 = w_sys_ce;
	assign w_sys_tmp1 = 32'h3c000000;
	assign w_sys_tmp3 = 32'h3ba3d70a;
	assign w_sys_tmp4 = 32'h42a3d70a;
	assign w_sys_tmp6 = 32'sh00000002;
	assign w_sys_tmp7 = ( !w_sys_tmp8 );
	assign w_sys_tmp8 = (w_sys_tmp9 < r_run_k_7);
	assign w_sys_tmp9 = 32'sh00000080;
	assign w_sys_tmp10 = (r_run_k_7 + w_sys_intOne);
	assign w_sys_tmp11 = 32'sh00000002;
	assign w_sys_tmp12 = ( !w_sys_tmp13 );
	assign w_sys_tmp13 = (w_sys_tmp14 < r_run_j_8);
	assign w_sys_tmp14 = 32'sh00000041;
	assign w_sys_tmp17 = (r_run_j_8 * w_sys_tmp18);
	assign w_sys_tmp18 = 32'sh00000081;
	assign w_sys_tmp19 = w_ip_AddFloat_result_0;
	assign w_sys_tmp20 = (w_sys_tmp21 + r_run_k_7);
	assign w_sys_tmp21 = (r_run_copy7_j_26 * w_sys_tmp18);
	assign w_sys_tmp23 = w_ip_MultFloat_product_0;
	assign w_sys_tmp25 = (w_sys_tmp26 * w_sys_tmp18);
	assign w_sys_tmp26 = (r_run_copy6_j_25 + w_sys_intOne);
	assign w_sys_tmp29 = 32'h40000000;
	assign w_sys_tmp30 = w_fld_u_0_dataout_1;
	assign w_sys_tmp31 = (r_run_copy5_j_24 * w_sys_tmp18);
	assign w_sys_tmp33 = (w_sys_tmp34 * w_sys_tmp18);
	assign w_sys_tmp34 = (r_run_copy4_j_23 - w_sys_intOne);
	assign w_sys_tmp38 = (w_sys_tmp39 + r_run_k_7);
	assign w_sys_tmp39 = (r_run_copy3_j_22 * w_sys_tmp18);
	assign w_sys_tmp44 = (r_run_copy2_j_21 * w_sys_tmp18);
	assign w_sys_tmp46 = (w_sys_tmp47 + r_run_k_7);
	assign w_sys_tmp47 = (r_run_copy1_j_20 * w_sys_tmp18);
	assign w_sys_tmp50 = 32'h42c80000;
	assign w_sys_tmp51 = (r_run_copy0_j_19 + w_sys_tmp52);
	assign w_sys_tmp52 = 32'sh0000003e;
	assign w_sys_tmp53 = (r_run_k_7 - w_sys_intOne);
	assign w_sys_tmp54 = (r_run_copy0_j_19 + w_sys_intOne);
	assign w_sys_tmp55 = (r_run_copy1_j_20 + w_sys_intOne);
	assign w_sys_tmp56 = (r_run_copy2_j_21 + w_sys_intOne);
	assign w_sys_tmp57 = (r_run_copy3_j_22 + w_sys_intOne);
	assign w_sys_tmp58 = (r_run_copy4_j_23 + w_sys_intOne);
	assign w_sys_tmp59 = (r_run_copy5_j_24 + w_sys_intOne);
	assign w_sys_tmp61 = (r_run_copy7_j_26 + w_sys_intOne);
	assign w_sys_tmp62 = (r_run_j_8 + w_sys_intOne);
	assign w_sys_tmp64 = (w_sys_tmp65 * w_sys_tmp18);
	assign w_sys_tmp65 = w_sys_tmp62;
	assign w_sys_tmp68 = (w_sys_tmp69 * w_sys_tmp18);
	assign w_sys_tmp69 = w_sys_tmp61;
	assign w_sys_tmp72 = (w_sys_tmp73 * w_sys_tmp18);
	assign w_sys_tmp73 = (w_sys_tmp74 + w_sys_intOne);
	assign w_sys_tmp74 = w_sys_tmp26;
	assign w_sys_tmp79 = (w_sys_tmp80 * w_sys_tmp18);
	assign w_sys_tmp80 = w_sys_tmp59;
	assign w_sys_tmp82 = (w_sys_tmp83 * w_sys_tmp18);
	assign w_sys_tmp83 = (w_sys_tmp84 - w_sys_intOne);
	assign w_sys_tmp84 = w_sys_tmp58;
	assign w_sys_tmp87 = (w_sys_tmp88 + r_run_k_7);
	assign w_sys_tmp88 = (w_sys_tmp89 * w_sys_tmp18);
	assign w_sys_tmp89 = w_sys_tmp57;
	assign w_sys_tmp94 = (w_sys_tmp95 * w_sys_tmp18);
	assign w_sys_tmp95 = w_sys_tmp56;
	assign w_sys_tmp97 = (w_sys_tmp98 + r_run_k_7);
	assign w_sys_tmp98 = (w_sys_tmp99 * w_sys_tmp18);
	assign w_sys_tmp99 = w_sys_tmp55;
	assign w_sys_tmp102 = w_sys_tmp54;
	assign w_sys_tmp1707 = 32'sh00000002;
	assign w_sys_tmp1708 = ( !w_sys_tmp1709 );
	assign w_sys_tmp1709 = (w_sys_tmp1710 < r_run_k_7);
	assign w_sys_tmp1710 = 32'sh00000080;
	assign w_sys_tmp1711 = (r_run_k_7 + w_sys_intOne);
	assign w_sys_tmp1712 = 32'sh00000002;
	assign w_sys_tmp1713 = ( !w_sys_tmp1714 );
	assign w_sys_tmp1714 = (w_sys_tmp1715 < r_run_j_8);
	assign w_sys_tmp1715 = 32'sh00000041;
	assign w_sys_tmp1718 = (r_run_j_8 * w_sys_tmp1719);
	assign w_sys_tmp1719 = 32'sh00000081;
	assign w_sys_tmp1720 = w_fld_result_1_dataout_1;
	assign w_sys_tmp1721 = (w_sys_tmp1722 + r_run_k_7);
	assign w_sys_tmp1722 = (r_run_copy0_j_27 * w_sys_tmp1719);
	assign w_sys_tmp1724 = (r_run_copy0_j_27 + w_sys_intOne);
	assign w_sys_tmp1725 = (r_run_j_8 + w_sys_intOne);
	assign w_sys_tmp1727 = (w_sys_tmp1728 * w_sys_tmp1719);
	assign w_sys_tmp1728 = w_sys_tmp1725;
	assign w_sys_tmp1731 = (w_sys_tmp1732 * w_sys_tmp1719);
	assign w_sys_tmp1732 = w_sys_tmp1724;
	assign w_sys_tmp2036 = (r_run_k_7 < w_sys_tmp2037);
	assign w_sys_tmp2037 = 32'sh00000081;
	assign w_sys_tmp2039 = w_ip_fifo_under2up_result_0;
	assign w_sys_tmp2040 = w_fld_u_0_dataout_1;
	assign w_sys_tmp2041 = (w_sys_tmp2042 + r_run_k_7);
	assign w_sys_tmp2042 = 32'sh00002040;
	assign w_sys_tmp2043 = (r_run_k_7 + w_sys_intOne);
	assign w_sys_tmp2044 = (r_run_k_7 < w_sys_tmp2045);
	assign w_sys_tmp2045 = 32'sh00000081;
	assign w_sys_tmp2048 = 32'sh000020c1;
	assign w_sys_tmp2049 = w_ip_fifo_up2under_result_0;
	assign w_sys_tmp2050 = 32'h0;
	assign w_sys_tmp2051 = (r_run_k_7 + w_sys_intOne);
	assign w_sys_tmp2052 = 32'h0;
	assign w_sys_tmp2053 = 32'h0;
	assign w_sys_tmp2054 = 32'h0;
	assign w_sys_tmp2055 = 32'h0;
	assign w_sys_tmp2056 = 32'h0;
	assign w_sys_tmp2057 = (w_sys_tmp17 + r_run_k_7);
	assign w_sys_tmp2058 = (w_sys_tmp25 + r_run_k_7);
	assign w_sys_tmp2059 = (w_sys_tmp31 + r_run_k_7);
	assign w_sys_tmp2060 = (w_sys_tmp33 + r_run_k_7);
	assign w_sys_tmp2061 = (w_sys_tmp38 + w_sys_intOne);
	assign w_sys_tmp2062 = (w_sys_tmp44 + r_run_k_7);
	assign w_sys_tmp2063 = (w_sys_tmp46 - w_sys_intOne);
	assign w_sys_tmp2064 = (w_sys_tmp64 + r_run_k_7);
	assign w_sys_tmp2065 = (w_sys_tmp68 + r_run_k_7);
	assign w_sys_tmp2066 = (w_sys_tmp72 + r_run_k_7);
	assign w_sys_tmp2067 = (w_sys_tmp79 + r_run_k_7);
	assign w_sys_tmp2068 = (w_sys_tmp82 + r_run_k_7);
	assign w_sys_tmp2069 = (w_sys_tmp87 + w_sys_intOne);
	assign w_sys_tmp2070 = (w_sys_tmp94 + r_run_k_7);
	assign w_sys_tmp2071 = (w_sys_tmp97 - w_sys_intOne);
	assign w_sys_tmp2072 = (w_sys_tmp102 + w_sys_tmp52);
	assign w_sys_tmp2343 = (w_sys_tmp1718 + r_run_k_7);
	assign w_sys_tmp2344 = (w_sys_tmp1727 + r_run_k_7);
	assign w_sys_tmp2345 = (w_sys_tmp1731 + r_run_k_7);
	assign w_sys_tmp2406 = (w_sys_tmp2048 + r_run_k_7);


	DualPortRAM #(.DWIDTH(32), .AWIDTH(14), .WORDS(8643) )
		dpram_u_0(
			.clk (clock),
			.ce_0 (w_fld_u_0_ce_0),
			.addr_0 (w_fld_u_0_addr_0),
			.datain_0 (w_fld_u_0_datain_0),
			.dataout_0 (w_fld_u_0_dataout_0),
			.r_w_0 (w_fld_u_0_r_w_0),
			.ce_1 (w_fld_u_0_ce_1),
			.addr_1 (r_fld_u_0_addr_1),
			.datain_1 (r_fld_u_0_datain_1),
			.dataout_1 (w_fld_u_0_dataout_1),
			.r_w_1 (r_fld_u_0_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(14), .WORDS(8643) )
		dpram_result_1(
			.clk (clock),
			.ce_0 (w_fld_result_1_ce_0),
			.addr_0 (w_fld_result_1_addr_0),
			.datain_0 (w_fld_result_1_datain_0),
			.dataout_0 (w_fld_result_1_dataout_0),
			.r_w_0 (w_fld_result_1_r_w_0),
			.ce_1 (w_fld_result_1_ce_1),
			.addr_1 (r_fld_result_1_addr_1),
			.datain_1 (r_fld_result_1_datain_1),
			.dataout_1 (w_fld_result_1_dataout_1),
			.r_w_1 (r_fld_result_1_r_w_1)
		);

	AddFloat
		AddFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_AddFloat_portA_0),
			.b (r_ip_AddFloat_portB_0),
			.result (w_ip_AddFloat_result_0)
		);

	MultFloat
		MultFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_MultFloat_multiplicand_0),
			.b (r_ip_MultFloat_multiplier_0),
			.result (w_ip_MultFloat_product_0)
		);

	FixedToFloat
		FixedToFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_FixedToFloat_fixed_0),
			.result (w_ip_FixedToFloat_floating_0)
		);
/*
	fifo_under2up
		fifo_under2up_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.operation_nd (r_ip_fifo_under2up_newData_0),
			.in (r_ip_fifo_under2up_in_0),	// in 32bit
			.s_we (r_ip_fifo_under2up_s_we_0),	// in 32bit
			.s_re (r_ip_fifo_under2up_s_re_0),	// in 32bit
			.p (w_ip_fifo_under2up_result_0)	// out 32bit
		);

	fifo_up2under
		fifo_up2under_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.operation_nd (r_ip_fifo_up2under_newData_0),
			.in (r_ip_fifo_up2under_in_0),	// in 32bit
			.s_we (r_ip_fifo_up2under_s_we_0),	// in 32bit
			.s_re (r_ip_fifo_up2under_s_re_0),	// in 32bit
			.p (w_ip_fifo_up2under_result_0)	// out 32bit
		);
*/
	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h8a) || (r_sys_run_step==9'h91) || (r_sys_run_step==9'h98) || (r_sys_run_step==9'hbf) || (r_sys_run_step==9'hf9)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp86_float;

									end
									else
									if((r_sys_run_step==9'h13) || (r_sys_run_step==9'h3a) || (r_sys_run_step==9'h55) || (r_sys_run_step==9'h72) || (r_sys_run_step==9'ha4) || (r_sys_run_step==9'haa) || (r_sys_run_step==9'he9)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp87_float;

									end
									else
									if((r_sys_run_step==9'ha5) || (r_sys_run_step==9'hec)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp48_float;

									end
									else
									if((r_sys_run_step==9'h40) || (r_sys_run_step==9'hf8) || (r_sys_run_step==9'h10c) || (r_sys_run_step==9'h11c)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp75_float;

									end
									else
									if((r_sys_run_step==9'h5c) || (r_sys_run_step==9'h110) || (r_sys_run_step==9'h11f) || (r_sys_run_step==9'h123)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp72_float;

									end
									else
									if((r_sys_run_step==9'h1a) || (r_sys_run_step==9'h41) || (r_sys_run_step==9'h5f) || (r_sys_run_step==9'h79) || (r_sys_run_step==9'hae) || (r_sys_run_step==9'hb4) || (r_sys_run_step==9'hcd) || (r_sys_run_step==9'h103)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp93_float;

									end
									else
									if((r_sys_run_step==9'h84) || (r_sys_run_step==9'hb5) || (r_sys_run_step==9'he3) || (r_sys_run_step==9'he8) || (r_sys_run_step==9'hfd) || (r_sys_run_step==9'h113) || (r_sys_run_step==9'h120)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp77_float;

									end
									else
									if((r_sys_run_step==9'hc3) || (r_sys_run_step==9'he6)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp55_float;

									end
									else
									if((r_sys_run_step==9'ha6) || (r_sys_run_step==9'had) || (r_sys_run_step==9'hee)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp49_float;

									end
									else
									if((r_sys_run_step==9'hd3)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp52_float;

									end
									else
									if((r_sys_run_step==9'hb9) || (r_sys_run_step==9'hba) || (r_sys_run_step==9'hdd)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp69_float;

									end
									else
									if((r_sys_run_step==9'hb0)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp51_float;

									end
									else
									if((r_sys_run_step==9'h63) || (r_sys_run_step==9'h89) || (r_sys_run_step==9'h116)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp65_float;

									end
									else
									if((r_sys_run_step==9'h8d) || (r_sys_run_step==9'hbe)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp53_float;

									end
									else
									if((r_sys_run_step==9'h21) || (r_sys_run_step==9'h28) || (r_sys_run_step==9'h52) || (r_sys_run_step==9'h59) || (r_sys_run_step==9'h60) || (r_sys_run_step==9'h67) || (r_sys_run_step==9'h80) || (r_sys_run_step==9'hb7) || (r_sys_run_step==9'hde)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp92_float;

									end
									else
									if((r_sys_run_step==9'h7b) || (r_sys_run_step==9'hab) || (r_sys_run_step==9'hac) || (r_sys_run_step==9'hda) || (r_sys_run_step==9'hfc) || (r_sys_run_step==9'h111) || (r_sys_run_step==9'h11d)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp71_float;

									end
									else
									if((r_sys_run_step==9'h51) || (r_sys_run_step==9'hc8) || (r_sys_run_step==9'hf1) || (r_sys_run_step==9'h10b) || (r_sys_run_step==9'h11a)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp70_float;

									end
									else
									if((r_sys_run_step==9'h17) || (r_sys_run_step==9'h2e) || (r_sys_run_step==9'h48) || (r_sys_run_step==9'h68) || (r_sys_run_step==9'h6e) || (r_sys_run_step==9'h87) || (r_sys_run_step==9'hc0) || (r_sys_run_step==9'hc6) || (r_sys_run_step==9'hfe)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp91_float;

									end
									else
									if((r_sys_run_step==9'hf7)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp39_float;

									end
									else
									if((r_sys_run_step==9'h1e) || (r_sys_run_step==9'h35) || (r_sys_run_step==9'h4f) || (r_sys_run_step==9'h74) || (r_sys_run_step==9'h8e) || (r_sys_run_step==9'hca) || (r_sys_run_step==9'hd0)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp95_float;

									end
									else
									if((r_sys_run_step==9'hd8)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp74_float;

									end
									else
									if((r_sys_run_step==9'hb1) || (r_sys_run_step==9'hbb) || (r_sys_run_step==9'hc2) || (r_sys_run_step==9'hc9) || (r_sys_run_step==9'he5)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp79_float;

									end
									else
									if((r_sys_run_step==9'h9) || (r_sys_run_step==9'h24) || (r_sys_run_step==9'h33) || (r_sys_run_step==9'h4e) || (r_sys_run_step==9'h5d) || (r_sys_run_step==9'h86) || (r_sys_run_step==9'h95) || (r_sys_run_step==9'hd5) || (r_sys_run_step==9'hdb) || (r_sys_run_step==9'h10d)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp90_float;

									end
									else
									if((r_sys_run_step==9'hc) || (r_sys_run_step==9'h25) || (r_sys_run_step==9'h3c) || (r_sys_run_step==9'h56) || (r_sys_run_step==9'h7d) || (r_sys_run_step==9'h83) || (r_sys_run_step==9'h9c) || (r_sys_run_step==9'hdc) || (r_sys_run_step==9'he2)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp94_float;

									end
									else
									if((r_sys_run_step==9'h71) || (r_sys_run_step==9'ha2) || (r_sys_run_step==9'h106)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp45_float;

									end
									else
									if((r_sys_run_step==9'h7f) || (r_sys_run_step==9'heb) || (r_sys_run_step==9'h102)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp43_float;

									end
									else
									if((r_sys_run_step==9'he) || (r_sys_run_step==9'h11) || (r_sys_run_step==9'h15) || (r_sys_run_step==9'h18) || (r_sys_run_step==9'h1c) || (r_sys_run_step==9'h1f) || (r_sys_run_step==9'h23) || (r_sys_run_step==9'h26) || (r_sys_run_step==9'h2a) || (r_sys_run_step==9'h2d) || (r_sys_run_step==9'h31) || (r_sys_run_step==9'h34) || (r_sys_run_step==9'h38) || (r_sys_run_step==9'h3b) || (r_sys_run_step==9'h3f) || (r_sys_run_step==9'h42) || (r_sys_run_step==9'h46) || (r_sys_run_step==9'h49) || (r_sys_run_step==9'h4d) || (r_sys_run_step==9'h50) || (r_sys_run_step==9'h54) || (r_sys_run_step==9'h57) || (r_sys_run_step==9'h5b) || (r_sys_run_step==9'h5e) || (r_sys_run_step==9'h62) || (r_sys_run_step==9'h65) || (r_sys_run_step==9'h69) || (r_sys_run_step==9'h6c) || (r_sys_run_step==9'h70) || (r_sys_run_step==9'h73) || (r_sys_run_step==9'h77) || (r_sys_run_step==9'h7a) || (r_sys_run_step==9'h7e) || (r_sys_run_step==9'h81) || (r_sys_run_step==9'h85) || (r_sys_run_step==9'h88) || (r_sys_run_step==9'h8c) || (r_sys_run_step==9'h8f) || (r_sys_run_step==9'h93) || (r_sys_run_step==9'h96) || (r_sys_run_step==9'h9a) || (r_sys_run_step==9'h9d) || (r_sys_run_step==9'ha1) || (r_sys_run_step==9'ha8) || (r_sys_run_step==9'haf) || (r_sys_run_step==9'hb2) || (r_sys_run_step==9'hb6) || (r_sys_run_step==9'hbd) || (r_sys_run_step==9'hc4) || (r_sys_run_step==9'hc7) || (r_sys_run_step==9'hcb) || (r_sys_run_step==9'hce) || (r_sys_run_step==9'hd2) || (r_sys_run_step==9'hd9) || (r_sys_run_step==9'he0) || (r_sys_run_step==9'he7) || (r_sys_run_step==9'hea)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp19;

									end
									else
									if((r_sys_run_step==9'h10) || (r_sys_run_step==9'h29) || (r_sys_run_step==9'h2f) || (r_sys_run_step==9'h36) || (r_sys_run_step==9'h3d) || (r_sys_run_step==9'h44) || (r_sys_run_step==9'h6b) || (r_sys_run_step==9'h99) || (r_sys_run_step==9'h9f) || (r_sys_run_step==9'hb8) || (r_sys_run_step==9'hf3)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp96_float;

									end
									else
									if((r_sys_run_step==9'h66) || (r_sys_run_step==9'h97)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp62_float;

									end
									else
									if((r_sys_run_step==9'h76) || (r_sys_run_step==9'h9b) || (r_sys_run_step==9'h101) || (r_sys_run_step==9'h114)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp60_float;

									end
									else
									if((r_sys_run_step==9'h75) || (r_sys_run_step==9'h7c) || (r_sys_run_step==9'ha3) || (r_sys_run_step==9'he4)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp73_float;

									end
									else
									if((r_sys_run_step==9'h37) || (r_sys_run_step==9'ha7) || (r_sys_run_step==9'hcc) || (r_sys_run_step==9'h117) || (r_sys_run_step==9'h122)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp76_float;

									end
									else
									if((r_sys_run_step==9'h6d) || (r_sys_run_step==9'h92) || (r_sys_run_step==9'hf2) || (r_sys_run_step==9'h107) || (r_sys_run_step==9'h119) || (r_sys_run_step==9'h121) || (r_sys_run_step==9'h124)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp88_float;

									end
									else
									if((r_sys_run_step==9'hd7)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp59_float;

									end
									else
									if((r_sys_run_step==9'hc1)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp54_float;

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp56_float;

									end
									else
									if((r_sys_run_step==9'hd6) || (r_sys_run_step==9'hdf)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp58_float;

									end
									else
									if((r_sys_run_step==9'h1d) || (r_sys_run_step==9'h2c) || (r_sys_run_step==9'h45) || (r_sys_run_step==9'h4b) || (r_sys_run_step==9'h64) || (r_sys_run_step==9'h90) || (r_sys_run_step==9'hd4) || (r_sys_run_step==9'h108)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp97_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'ha1) || (r_sys_run_step==9'ha2) || (r_sys_run_step==9'hac) || (r_sys_run_step==9'hb6)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp86_float;

									end
									else
									if((r_sys_run_step==9'h1c) || (r_sys_run_step==9'h2a) || (r_sys_run_step==9'h34) || (r_sys_run_step==9'h62) || (r_sys_run_step==9'h6c)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp87_float;

									end
									else
									if((r_sys_run_step==9'h5d)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'hd4)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h23) || (r_sys_run_step==9'h31) || (r_sys_run_step==9'h3b) || (r_sys_run_step==9'h69) || (r_sys_run_step==9'h73) || (r_sys_run_step==9'hbd) || (r_sys_run_step==9'hc7)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp93_float;

									end
									else
									if((r_sys_run_step==9'ha7) || (r_sys_run_step==9'hd5) || (r_sys_run_step==9'hd6)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp81_float;

									end
									else
									if((r_sys_run_step==9'had)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'hc9)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h36)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h4f)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h60)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'hbb)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h48)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'ha6)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h8e)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h1d) || (r_sys_run_step==9'h29) || (r_sys_run_step==9'h2e) || (r_sys_run_step==9'h37) || (r_sys_run_step==9'h3c) || (r_sys_run_step==9'h45) || (r_sys_run_step==9'h47) || (r_sys_run_step==9'h51) || (r_sys_run_step==9'h55) || (r_sys_run_step==9'h63) || (r_sys_run_step==9'h66) || (r_sys_run_step==9'h68) || (r_sys_run_step==9'h76) || (r_sys_run_step==9'h84) || (r_sys_run_step==9'h8d) || (r_sys_run_step==9'h92) || (r_sys_run_step==9'h97) || (r_sys_run_step==9'h99) || (r_sys_run_step==9'h9b) || (r_sys_run_step==9'hab) || (r_sys_run_step==9'hb5) || (r_sys_run_step==9'hb9) || (r_sys_run_step==9'hbe) || (r_sys_run_step==9'hc0) || (r_sys_run_step==9'hc3) || (r_sys_run_step==9'hc8) || (r_sys_run_step==9'hca) || (r_sys_run_step==9'hcc) || (r_sys_run_step==9'hda) || (r_sys_run_step==9'hdc) || (r_sys_run_step==9'hdd) || (r_sys_run_step==9'he3) || (r_sys_run_step==9'he4) || (r_sys_run_step==9'he6) || (r_sys_run_step==9'he9) || (r_sys_run_step==9'heb) || (r_sys_run_step==9'hec) || (r_sys_run_step==9'hee) || (r_sys_run_step==9'hf1) || (r_sys_run_step==9'hf2) || (r_sys_run_step==9'hf3) || (r_sys_run_step==9'hf7) || (r_sys_run_step==9'hf8) || (r_sys_run_step==9'hf9) || (r_sys_run_step==9'hfc) || (r_sys_run_step==9'hfd) || (r_sys_run_step==9'hfe) || (r_sys_run_step==9'h101) || (r_sys_run_step==9'h102) || (r_sys_run_step==9'h103) || (r_sys_run_step==9'h106) || (r_sys_run_step==9'h107) || (r_sys_run_step==9'h108) || (r_sys_run_step==9'h10b) || (r_sys_run_step==9'h10c) || (r_sys_run_step==9'h10d) || (r_sys_run_step==9'h110) || (r_sys_run_step==9'h111) || (r_sys_run_step==9'h113) || (r_sys_run_step==9'h114) || (r_sys_run_step==9'h116) || (r_sys_run_step==9'h117) || (r_sys_run_step==9'h119) || (r_sys_run_step==9'h11a) || (r_sys_run_step==9'h11c) || (r_sys_run_step==9'h11d) || (9'h11f<=r_sys_run_step && r_sys_run_step<=9'h124)) begin
										r_ip_AddFloat_portB_0 <= w_sys_tmp23;

									end
									else
									if((r_sys_run_step==9'h64)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'hd2) || (r_sys_run_step==9'hdf)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp79_float;

									end
									else
									if((r_sys_run_step==9'hae)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp84_float;

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h9f)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h59)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h4d) || (r_sys_run_step==9'h5b) || (r_sys_run_step==9'h65) || (r_sys_run_step==9'ha8) || (r_sys_run_step==9'hb2)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp96_float;

									end
									else
									if((r_sys_run_step==9'h87)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h44)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h28)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h56)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'hb8)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'hd7)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h85) || (r_sys_run_step==9'h93) || (r_sys_run_step==9'h9d)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp73_float;

									end
									else
									if((r_sys_run_step==9'h7f) || (r_sys_run_step==9'hb0)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp83_float;

									end
									else
									if((r_sys_run_step==9'hb1)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'hd0)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h2c)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'hde)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h3a)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h26) || (r_sys_run_step==9'h54) || (r_sys_run_step==9'h5e) || (r_sys_run_step==9'h9a) || (r_sys_run_step==9'ha5) || (r_sys_run_step==9'haf) || (r_sys_run_step==9'hba) || (r_sys_run_step==9'hc4) || (r_sys_run_step==9'hce)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp97_float;

									end
									else
									if((r_sys_run_step==9'h33)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'hb4)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h67)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h75)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h83)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h91)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h90)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp78_float;

									end
									else
									if((r_sys_run_step==9'h80)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h8a)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h40)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp67_float;

									end
									else
									if((r_sys_run_step==9'he2)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h98)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h7b) || (r_sys_run_step==9'h7d)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp66_float;

									end
									else
									if((r_sys_run_step==9'hdb)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'hbf)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h70) || (r_sys_run_step==9'h7a) || (r_sys_run_step==9'hc1) || (r_sys_run_step==9'hcb) || (r_sys_run_step==9'hd8) || (r_sys_run_step==9'he7)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp92_float;

									end
									else
									if((r_sys_run_step==9'h7c)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h41)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h11) || (r_sys_run_step==9'h38) || (r_sys_run_step==9'h42) || (r_sys_run_step==9'h77) || (r_sys_run_step==9'h81)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp91_float;

									end
									else
									if((r_sys_run_step==9'h6b)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'he) || (r_sys_run_step==9'h18) || (r_sys_run_step==9'h3f) || (r_sys_run_step==9'h49) || (r_sys_run_step==9'h7e) || (r_sys_run_step==9'h88) || (r_sys_run_step==9'hd9) || (r_sys_run_step==9'he8)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp95_float;

									end
									else
									if((r_sys_run_step==9'he5)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h5c) || (r_sys_run_step==9'h71) || (r_sys_run_step==9'h74)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp74_float;

									end
									else
									if((r_sys_run_step==9'h79)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h2d) || (r_sys_run_step==9'h57) || (r_sys_run_step==9'h8f)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp90_float;

									end
									else
									if((r_sys_run_step==9'h95)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'hc2)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h15) || (r_sys_run_step==9'h1f) || (r_sys_run_step==9'h46) || (r_sys_run_step==9'h50) || (r_sys_run_step==9'h8c) || (r_sys_run_step==9'h96)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp94_float;

									end
									else
									if((r_sys_run_step==9'h35) || (r_sys_run_step==9'h89)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp82_float;

									end
									else
									if((r_sys_run_step==9'h5f)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp68_float;

									end
									else
									if((r_sys_run_step==9'haa)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h6d) || (r_sys_run_step==9'hd3)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp61_float;

									end
									else
									if((r_sys_run_step==9'hc6)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h21)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h6e)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'hcd)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h9c)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h24) || (r_sys_run_step==9'ha4)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp80_float;

									end
									else
									if((r_sys_run_step==9'h86) || (r_sys_run_step==9'hb7)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp63_float;

									end
									else
									if((r_sys_run_step==9'h72)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'he0) || (r_sys_run_step==9'hea)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp59_float;

									end
									else
									if((r_sys_run_step==9'ha3)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp23[31], w_sys_tmp23[30:0] };

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp44_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hd) || (r_sys_run_step==9'h17) || (r_sys_run_step==9'h2d) || (r_sys_run_step==9'h4f) || (r_sys_run_step==9'h7c) || (r_sys_run_step==9'hab) || (r_sys_run_step==9'hda) || (r_sys_run_step==9'hfa) || (r_sys_run_step==9'h10d) || (r_sys_run_step==9'h119)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp84_float;

									end
									else
									if((r_sys_run_step==9'h33) || (r_sys_run_step==9'h5d) || (r_sys_run_step==9'h8e) || (r_sys_run_step==9'hc2) || (r_sys_run_step==9'heb) || (r_sys_run_step==9'h104)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp68_float;

									end
									else
									if((r_sys_run_step==9'h1b) || (r_sys_run_step==9'h34) || (r_sys_run_step==9'h5c) || (r_sys_run_step==9'h88) || (r_sys_run_step==9'hb7) || (r_sys_run_step==9'he2) || (r_sys_run_step==9'hff) || (r_sys_run_step==9'h110) || (r_sys_run_step==9'h11d)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp82_float;

									end
									else
									if((r_sys_run_step==9'h87) || (r_sys_run_step==9'hb9) || (r_sys_run_step==9'he6)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp41_float;

									end
									else
									if((r_sys_run_step==9'h57) || (r_sys_run_step==9'h86) || (r_sys_run_step==9'hb8) || (r_sys_run_step==9'he5)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp47_float;

									end
									else
									if((r_sys_run_step==9'h47) || (r_sys_run_step==9'h73) || (r_sys_run_step==9'ha3) || (r_sys_run_step==9'hd4) || (r_sys_run_step==9'hf6)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp57_float;

									end
									else
									if((r_sys_run_step==9'h8) || (r_sys_run_step==9'h10) || (r_sys_run_step==9'h21) || (r_sys_run_step==9'h3e) || (r_sys_run_step==9'h65) || (r_sys_run_step==9'h92) || (r_sys_run_step==9'hc0) || (r_sys_run_step==9'he8) || (r_sys_run_step==9'h100) || (r_sys_run_step==9'h111) || (r_sys_run_step==9'h11b) || (r_sys_run_step==9'h11e) || (r_sys_run_step==9'h11f)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp89_float;

									end
									else
									if((r_sys_run_step==9'h1d) || (r_sys_run_step==9'h3b) || (r_sys_run_step==9'h61) || (r_sys_run_step==9'h8f) || (r_sys_run_step==9'hbf) || (r_sys_run_step==9'hea) || (r_sys_run_step==9'h101) || (r_sys_run_step==9'h113)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp78_float;

									end
									else
									if((r_sys_run_step==9'h6b) || (r_sys_run_step==9'h9b) || (r_sys_run_step==9'hcd) || (r_sys_run_step==9'hf7)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp61_float;

									end
									else
									if((r_sys_run_step==9'h32) || (r_sys_run_step==9'h3a) || (r_sys_run_step==9'h42) || (r_sys_run_step==9'h4c) || (r_sys_run_step==9'h56) || (r_sys_run_step==9'h5e) || (r_sys_run_step==9'h67) || (r_sys_run_step==9'h71) || (r_sys_run_step==9'h79) || (r_sys_run_step==9'h83) || (r_sys_run_step==9'h8d) || (r_sys_run_step==9'h96) || (r_sys_run_step==9'ha0) || (r_sys_run_step==9'haa) || (r_sys_run_step==9'hb4) || (r_sys_run_step==9'hbe) || (r_sys_run_step==9'hc7) || (r_sys_run_step==9'hd0) || (r_sys_run_step==9'hd8) || (r_sys_run_step==9'he1) || (r_sys_run_step==9'he7) || (r_sys_run_step==9'hed) || (r_sys_run_step==9'hf3) || (r_sys_run_step==9'hf8) || (r_sys_run_step==9'hfd) || (r_sys_run_step==9'h102) || (r_sys_run_step==9'h107) || (r_sys_run_step==9'h10c) || (r_sys_run_step==9'h10f) || (r_sys_run_step==9'h112) || (r_sys_run_step==9'h115) || (r_sys_run_step==9'h118)) begin
										r_ip_MultFloat_multiplicand_0 <= r_fld_r2_3;

									end
									else
									if((r_sys_run_step==9'h3d) || (r_sys_run_step==9'h68) || (r_sys_run_step==9'h98) || (r_sys_run_step==9'hc9) || (r_sys_run_step==9'hf0) || (r_sys_run_step==9'h10b)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp67_float;

									end
									else
									if((r_sys_run_step==9'h36) || (r_sys_run_step==9'h60) || (r_sys_run_step==9'h91) || (r_sys_run_step==9'hc3) || (r_sys_run_step==9'hec) || (r_sys_run_step==9'h106)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp64_float;

									end
									else
									if((r_sys_run_step==9'h28) || (r_sys_run_step==9'h4b) || (r_sys_run_step==9'h75) || (r_sys_run_step==9'ha4) || (r_sys_run_step==9'hd3) || (r_sys_run_step==9'hf5) || (r_sys_run_step==9'h10a) || (r_sys_run_step==9'h117)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp81_float;

									end
									else
									if((r_sys_run_step==9'h4e) || (r_sys_run_step==9'h7a) || (r_sys_run_step==9'hae) || (r_sys_run_step==9'hdc) || (r_sys_run_step==9'hfc)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp66_float;

									end
									else
									if((r_sys_run_step==9'h6a) || (r_sys_run_step==9'h99) || (r_sys_run_step==9'hcc) || (r_sys_run_step==9'hf1)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp46_float;

									end
									else
									if((r_sys_run_step==9'ha) || (r_sys_run_step==9'h13) || (r_sys_run_step==9'h26) || (r_sys_run_step==9'h45) || (r_sys_run_step==9'h6f) || (r_sys_run_step==9'h9c) || (r_sys_run_step==9'hca) || (r_sys_run_step==9'hef) || (r_sys_run_step==9'h105) || (r_sys_run_step==9'h114) || (r_sys_run_step==9'h11c)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp85_float;

									end
									else
									if((r_sys_run_step==9'h16) || (r_sys_run_step==9'h2c) || (r_sys_run_step==9'h53) || (r_sys_run_step==9'h7d) || (r_sys_run_step==9'had) || (r_sys_run_step==9'hdb) || (r_sys_run_step==9'hfb) || (r_sys_run_step==9'h10e) || (r_sys_run_step==9'h11a)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp83_float;

									end
									else
									if((r_sys_run_step==9'h22) || (r_sys_run_step==9'h44) || (r_sys_run_step==9'h72) || (r_sys_run_step==9'ha2) || (r_sys_run_step==9'hd1) || (r_sys_run_step==9'hf2) || (r_sys_run_step==9'h109) || (r_sys_run_step==9'h116)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp80_float;

									end
									else
									if((r_sys_run_step==9'h55) || (r_sys_run_step==9'h84) || (r_sys_run_step==9'hb5) || (r_sys_run_step==9'he3)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp63_float;

									end
									else
									if((r_sys_run_step==9'h4) || (r_sys_run_step==9'h7) || (r_sys_run_step==9'hb) || (r_sys_run_step==9'he) || (r_sys_run_step==9'h12) || (r_sys_run_step==9'h15) || (r_sys_run_step==9'h19) || (r_sys_run_step==9'h1c) || (r_sys_run_step==9'h20) || (r_sys_run_step==9'h23) || (r_sys_run_step==9'h27) || (r_sys_run_step==9'h2a) || (r_sys_run_step==9'h2e) || (r_sys_run_step==9'h31) || (r_sys_run_step==9'h35) || (r_sys_run_step==9'h38) || (r_sys_run_step==9'h3c) || (r_sys_run_step==9'h3f) || (r_sys_run_step==9'h43) || (r_sys_run_step==9'h46) || (r_sys_run_step==9'h4a) || (r_sys_run_step==9'h4d) || (r_sys_run_step==9'h51) || (r_sys_run_step==9'h54) || (r_sys_run_step==9'h58) || (r_sys_run_step==9'h5b) || (r_sys_run_step==9'h5f) || (r_sys_run_step==9'h62) || (r_sys_run_step==9'h66) || (r_sys_run_step==9'h69) || (r_sys_run_step==9'h6d) || (r_sys_run_step==9'h70) || (r_sys_run_step==9'h74) || (r_sys_run_step==9'h77) || (r_sys_run_step==9'h7b) || (r_sys_run_step==9'h7e) || (r_sys_run_step==9'h82) || (r_sys_run_step==9'h85) || (r_sys_run_step==9'h89) || (r_sys_run_step==9'h8c) || (r_sys_run_step==9'h90) || (r_sys_run_step==9'h93) || (r_sys_run_step==9'h97) || (r_sys_run_step==9'h9a) || (r_sys_run_step==9'h9e) || (r_sys_run_step==9'ha1) || (r_sys_run_step==9'ha5) || (r_sys_run_step==9'ha8) || (r_sys_run_step==9'hac) || (r_sys_run_step==9'haf) || (r_sys_run_step==9'hb3) || (r_sys_run_step==9'hb6) || (r_sys_run_step==9'hba) || (r_sys_run_step==9'hbd) || (r_sys_run_step==9'hc1) || (r_sys_run_step==9'hc4) || (r_sys_run_step==9'hc8) || (r_sys_run_step==9'hcb) || (r_sys_run_step==9'hcf) || (r_sys_run_step==9'hd2) || (r_sys_run_step==9'hd6) || (r_sys_run_step==9'hd9) || (r_sys_run_step==9'hdd) || (r_sys_run_step==9'he0)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp29;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h3) || (r_sys_run_step==9'h5) || (r_sys_run_step==9'h6) || (r_sys_run_step==9'h9) || (r_sys_run_step==9'hc) || (r_sys_run_step==9'hf) || (r_sys_run_step==9'h11) || (r_sys_run_step==9'h14) || (r_sys_run_step==9'h1a) || (r_sys_run_step==9'h1f) || (r_sys_run_step==9'h25) || (r_sys_run_step==9'h2b) || (r_sys_run_step==9'h30) || (r_sys_run_step==9'h39) || (r_sys_run_step==9'h41) || (r_sys_run_step==9'h49) || (r_sys_run_step==9'h52) || (r_sys_run_step==9'h5a) || (r_sys_run_step==9'h64) || (r_sys_run_step==9'h6e) || (r_sys_run_step==9'h78) || (r_sys_run_step==9'h81) || (r_sys_run_step==9'h8b) || (r_sys_run_step==9'h95) || (r_sys_run_step==9'h9f) || (r_sys_run_step==9'ha9) || (r_sys_run_step==9'hb2) || (r_sys_run_step==9'hbc) || (r_sys_run_step==9'hc6)) begin
										r_ip_MultFloat_multiplicand_0 <= r_fld_dt_6;

									end
									else
									if((r_sys_run_step==9'h7f) || (r_sys_run_step==9'hb0) || (r_sys_run_step==9'hde)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp44_float;

									end
									else
									if((r_sys_run_step==9'h18) || (r_sys_run_step==9'h1e) || (r_sys_run_step==9'h24) || (r_sys_run_step==9'h29) || (r_sys_run_step==9'h2f) || (r_sys_run_step==9'h37) || (r_sys_run_step==9'h40) || (r_sys_run_step==9'h48) || (r_sys_run_step==9'h50) || (r_sys_run_step==9'h59) || (r_sys_run_step==9'h63) || (r_sys_run_step==9'h6c) || (r_sys_run_step==9'h76) || (r_sys_run_step==9'h80) || (r_sys_run_step==9'h8a) || (r_sys_run_step==9'h94) || (r_sys_run_step==9'h9d) || (r_sys_run_step==9'ha7) || (r_sys_run_step==9'hb1) || (r_sys_run_step==9'hbb) || (r_sys_run_step==9'hc5) || (r_sys_run_step==9'hce) || (r_sys_run_step==9'hd7) || (r_sys_run_step==9'hdf) || (r_sys_run_step==9'he4) || (r_sys_run_step==9'he9) || (r_sys_run_step==9'hee) || (r_sys_run_step==9'hf4) || (r_sys_run_step==9'hf9) || (r_sys_run_step==9'hfe) || (r_sys_run_step==9'h103) || (r_sys_run_step==9'h108)) begin
										r_ip_MultFloat_multiplicand_0 <= r_fld_r1_2;

									end
									else
									if((r_sys_run_step==9'ha6) || (r_sys_run_step==9'hd5)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp74_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hde)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp23_float;

									end
									else
									if((r_sys_run_step==9'h45) || (r_sys_run_step==9'h11e)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp35_float;

									end
									else
									if((r_sys_run_step==9'h17) || (r_sys_run_step==9'h7f)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp86_float;

									end
									else
									if((r_sys_run_step==9'h11f)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==9'h4) || (r_sys_run_step==9'h7) || (r_sys_run_step==9'hb) || (r_sys_run_step==9'he) || (r_sys_run_step==9'h12) || (r_sys_run_step==9'h15) || (r_sys_run_step==9'h19) || (r_sys_run_step==9'h1c) || (r_sys_run_step==9'h20) || (r_sys_run_step==9'h23) || (r_sys_run_step==9'h27) || (r_sys_run_step==9'h2a) || (r_sys_run_step==9'h2e) || (r_sys_run_step==9'h31) || (r_sys_run_step==9'h35) || (r_sys_run_step==9'h38) || (r_sys_run_step==9'h3c) || (r_sys_run_step==9'h3f) || (r_sys_run_step==9'h43) || (r_sys_run_step==9'h46) || (r_sys_run_step==9'h4a) || (r_sys_run_step==9'h4d) || (r_sys_run_step==9'h51) || (r_sys_run_step==9'h54) || (r_sys_run_step==9'h58) || (r_sys_run_step==9'h5b) || (r_sys_run_step==9'h5f) || (r_sys_run_step==9'h62) || (r_sys_run_step==9'h66) || (r_sys_run_step==9'h69) || (r_sys_run_step==9'h6d) || (r_sys_run_step==9'h70) || (r_sys_run_step==9'h74) || (r_sys_run_step==9'h77) || (r_sys_run_step==9'h7b) || (r_sys_run_step==9'h7e) || (r_sys_run_step==9'h82) || (r_sys_run_step==9'h85) || (r_sys_run_step==9'h89) || (r_sys_run_step==9'h8c) || (r_sys_run_step==9'h90) || (r_sys_run_step==9'h93) || (r_sys_run_step==9'h97) || (r_sys_run_step==9'h9a) || (r_sys_run_step==9'h9e) || (r_sys_run_step==9'ha1) || (r_sys_run_step==9'ha5) || (r_sys_run_step==9'ha8) || (r_sys_run_step==9'hac) || (r_sys_run_step==9'haf) || (r_sys_run_step==9'hb3) || (r_sys_run_step==9'hb6) || (r_sys_run_step==9'hba) || (r_sys_run_step==9'hbd) || (r_sys_run_step==9'hc1) || (r_sys_run_step==9'hc4) || (r_sys_run_step==9'hc8) || (r_sys_run_step==9'hcb) || (r_sys_run_step==9'hcf) || (r_sys_run_step==9'hd2) || (r_sys_run_step==9'hd6) || (r_sys_run_step==9'hd9) || (r_sys_run_step==9'hdd) || (r_sys_run_step==9'he0)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp30;

									end
									else
									if((r_sys_run_step==9'h29) || (r_sys_run_step==9'h67) || (r_sys_run_step==9'h76) || (r_sys_run_step==9'hb4) || (r_sys_run_step==9'hdf)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp75_float;

									end
									else
									if((r_sys_run_step==9'hf7)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==9'h99)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp49_float;

									end
									else
									if((r_sys_run_step==9'hf0)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==9'h5d) || (r_sys_run_step==9'ha0) || (r_sys_run_step==9'h10c)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp52_float;

									end
									else
									if((r_sys_run_step==9'h40) || (r_sys_run_step==9'ha7) || (r_sys_run_step==9'hd7) || (r_sys_run_step==9'hf9)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp65_float;

									end
									else
									if((r_sys_run_step==9'hb0)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp29_float;

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp71_float;

									end
									else
									if((r_sys_run_step==9'h6b)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp34_float;

									end
									else
									if((r_sys_run_step==9'he3)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp21_float;

									end
									else
									if((r_sys_run_step==9'hfc)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==9'h106)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==9'hb7) || (r_sys_run_step==9'hf8)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp40_float;

									end
									else
									if((r_sys_run_step==9'h2d) || (r_sys_run_step==9'he6)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp38_float;

									end
									else
									if((r_sys_run_step==9'h1d) || (r_sys_run_step==9'h9c)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp79_float;

									end
									else
									if((r_sys_run_step==9'hdb)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp22_float;

									end
									else
									if((r_sys_run_step==9'h101)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==9'h111)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==9'h37) || (r_sys_run_step==9'hbb) || (r_sys_run_step==9'he4) || (r_sys_run_step==9'h112)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp62_float;

									end
									else
									if((r_sys_run_step==9'h92) || (r_sys_run_step==9'hc5) || (r_sys_run_step==9'h102)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp42_float;

									end
									else
									if((r_sys_run_step==9'hd3)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp24_float;

									end
									else
									if((r_sys_run_step==9'h50) || (r_sys_run_step==9'he1)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp60_float;

									end
									else
									if((r_sys_run_step==9'h11a)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==9'ha6)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp30_float;

									end
									else
									if((r_sys_run_step==9'h68)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp73_float;

									end
									else
									if((r_sys_run_step==9'h36) || (r_sys_run_step==9'h3e) || (r_sys_run_step==9'h47) || (r_sys_run_step==9'h4f) || (r_sys_run_step==9'h57) || (r_sys_run_step==9'h60) || (r_sys_run_step==9'h6a) || (r_sys_run_step==9'h73) || (r_sys_run_step==9'h7d) || (r_sys_run_step==9'h87) || (r_sys_run_step==9'h91) || (r_sys_run_step==9'h9b) || (r_sys_run_step==9'ha4) || (r_sys_run_step==9'hae) || (r_sys_run_step==9'hb8) || (r_sys_run_step==9'hc2) || (r_sys_run_step==9'hcc) || (r_sys_run_step==9'hd4) || (r_sys_run_step==9'hdc) || (r_sys_run_step==9'he5) || (r_sys_run_step==9'heb) || (r_sys_run_step==9'hf1) || (r_sys_run_step==9'hf6) || (r_sys_run_step==9'hfb) || (r_sys_run_step==9'h100) || (r_sys_run_step==9'h105) || (r_sys_run_step==9'h10a) || (r_sys_run_step==9'h10d) || (r_sys_run_step==9'h110) || (r_sys_run_step==9'h113) || (r_sys_run_step==9'h116) || (r_sys_run_step==9'h119)) begin
										r_ip_MultFloat_multiplier_0 <= r_fld_dy_5;

									end
									else
									if((r_sys_run_step==9'h11d)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==9'h18) || (r_sys_run_step==9'h1e) || (r_sys_run_step==9'h24) || (r_sys_run_step==9'h42) || (r_sys_run_step==9'h48) || (r_sys_run_step==9'hd8)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp88_float;

									end
									else
									if((r_sys_run_step==9'hc0)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp26_float;

									end
									else
									if((r_sys_run_step==9'h114)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==9'h11c)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==9'hfa)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp14_float;

									end
									else
									if((r_sys_run_step==9'h22) || (r_sys_run_step==9'had) || (r_sys_run_step==9'he9)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp54_float;

									end
									else
									if((r_sys_run_step==9'h71) || (r_sys_run_step==9'haa) || (r_sys_run_step==9'hed) || (r_sys_run_step==9'h115)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp56_float;

									end
									else
									if((r_sys_run_step==9'h8f) || (r_sys_run_step==9'hb1) || (r_sys_run_step==9'h103)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp58_float;

									end
									else
									if((r_sys_run_step==9'ha3) || (r_sys_run_step==9'hce)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp48_float;

									end
									else
									if((r_sys_run_step==9'hec)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp20_float;

									end
									else
									if((r_sys_run_step==9'h7c)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp32_float;

									end
									else
									if((r_sys_run_step==9'h3a) || (r_sys_run_step==9'h8d) || (r_sys_run_step==9'hd0) || (r_sys_run_step==9'hf4)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp72_float;

									end
									else
									if((r_sys_run_step==9'h32) || (r_sys_run_step==9'h56)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp77_float;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h3) || (r_sys_run_step==9'h5) || (r_sys_run_step==9'h6) || (r_sys_run_step==9'h9) || (r_sys_run_step==9'hc) || (r_sys_run_step==9'hf) || (r_sys_run_step==9'h11) || (r_sys_run_step==9'h14) || (r_sys_run_step==9'h1a) || (r_sys_run_step==9'h1f) || (r_sys_run_step==9'h25) || (r_sys_run_step==9'h2b) || (r_sys_run_step==9'h30) || (r_sys_run_step==9'h39) || (r_sys_run_step==9'h41) || (r_sys_run_step==9'h49) || (r_sys_run_step==9'h52) || (r_sys_run_step==9'h5a) || (r_sys_run_step==9'h64) || (r_sys_run_step==9'h6e) || (r_sys_run_step==9'h78) || (r_sys_run_step==9'h81) || (r_sys_run_step==9'h8b) || (r_sys_run_step==9'h95) || (r_sys_run_step==9'h9f) || (r_sys_run_step==9'ha9) || (r_sys_run_step==9'hb2) || (r_sys_run_step==9'hbc) || (r_sys_run_step==9'hc6)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp50;

									end
									else
									if((r_sys_run_step==9'hf2)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp18_float;

									end
									else
									if((r_sys_run_step==9'h83) || (r_sys_run_step==9'h9d) || (r_sys_run_step==9'h108)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp55_float;

									end
									else
									if((r_sys_run_step==9'h4e) || (r_sys_run_step==9'h79) || (r_sys_run_step==9'h94) || (r_sys_run_step==9'h10f)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp69_float;

									end
									else
									if((r_sys_run_step==9'h72) || (r_sys_run_step==9'h8a) || (r_sys_run_step==9'hf3)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp51_float;

									end
									else
									if((r_sys_run_step==9'h3d) || (r_sys_run_step==9'h10e)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp36_float;

									end
									else
									if((r_sys_run_step==9'h86) || (r_sys_run_step==9'hc7) || (r_sys_run_step==9'hee) || (r_sys_run_step==9'h118)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp50_float;

									end
									else
									if((r_sys_run_step==9'h104)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==9'h61) || (r_sys_run_step==9'hfd)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp53_float;

									end
									else
									if((r_sys_run_step==9'h59) || (r_sys_run_step==9'h63) || (r_sys_run_step==9'h96)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp70_float;

									end
									else
									if((r_sys_run_step==9'hc3)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp27_float;

									end
									else
									if((r_sys_run_step==9'hcd)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp39_float;

									end
									else
									if((r_sys_run_step==9'h11b)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==9'h10b)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==9'h55) || (r_sys_run_step==9'hfe)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp74_float;

									end
									else
									if((r_sys_run_step==9'h88)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp31_float;

									end
									else
									if((r_sys_run_step==9'hd5)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp25_float;

									end
									else
									if((r_sys_run_step==9'he7)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp45_float;

									end
									else
									if((r_sys_run_step==9'hb9)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp28_float;

									end
									else
									if((r_sys_run_step==9'hbe)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp43_float;

									end
									else
									if((r_sys_run_step==9'hff)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==9'hea)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp19_float;

									end
									else
									if((r_sys_run_step==9'h34) || (r_sys_run_step==9'hf5)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp37_float;

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp19;

									end
									else
									if((r_sys_run_step==9'h109)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==9'h8) || (r_sys_run_step==9'ha) || (r_sys_run_step==9'hd) || (r_sys_run_step==9'h10) || (r_sys_run_step==9'h13) || (r_sys_run_step==9'h16) || (r_sys_run_step==9'h1b) || (r_sys_run_step==9'h21) || (r_sys_run_step==9'h26) || (r_sys_run_step==9'h2c) || (r_sys_run_step==9'h33) || (r_sys_run_step==9'h3b) || (r_sys_run_step==9'h44) || (r_sys_run_step==9'h4b) || (r_sys_run_step==9'h53) || (r_sys_run_step==9'h5c) || (r_sys_run_step==9'h65) || (r_sys_run_step==9'h6f) || (r_sys_run_step==9'h7a) || (r_sys_run_step==9'h84) || (r_sys_run_step==9'h8e) || (r_sys_run_step==9'h98) || (r_sys_run_step==9'ha2) || (r_sys_run_step==9'hab) || (r_sys_run_step==9'hb5) || (r_sys_run_step==9'hbf) || (r_sys_run_step==9'hc9) || (r_sys_run_step==9'hd1) || (r_sys_run_step==9'hda) || (r_sys_run_step==9'he2) || (r_sys_run_step==9'he8) || (r_sys_run_step==9'hef)) begin
										r_ip_MultFloat_multiplier_0 <= r_fld_dx_4;

									end
									else
									if((r_sys_run_step==9'h117)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==9'h5e) || (r_sys_run_step==9'h6c) || (r_sys_run_step==9'h80) || (r_sys_run_step==9'h107)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp76_float;

									end
									else
									if((r_sys_run_step==9'h28) || (r_sys_run_step==9'hca)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp59_float;

									end
									else
									if((r_sys_run_step==9'h75)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp33_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h31)) begin
										r_ip_FixedToFloat_fixed_0 <= r_sys_tmp15_int;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_ip_FixedToFloat_fixed_0 <= w_sys_tmp51;

									end
									else
									if((9'h1<=r_sys_run_step && r_sys_run_step<=9'h9) || (r_sys_run_step==9'hb) || (r_sys_run_step==9'hf) || (r_sys_run_step==9'h17) || (r_sys_run_step==9'h27)) begin
										r_ip_FixedToFloat_fixed_0 <= r_sys_tmp236_int;

									end
									else
									if((r_sys_run_step==9'h11) || (r_sys_run_step==9'h1b) || (r_sys_run_step==9'h2f)) begin
										r_ip_FixedToFloat_fixed_0 <= r_sys_tmp232_int;

									end
									else
									if((r_sys_run_step==9'h29)) begin
										r_ip_FixedToFloat_fixed_0 <= r_sys_tmp45_int;

									end
									else
									if((r_sys_run_step==9'h35)) begin
										r_ip_FixedToFloat_fixed_0 <= r_sys_tmp0_int;

									end
									else
									if((r_sys_run_step==9'h19) || (r_sys_run_step==9'h2b)) begin
										r_ip_FixedToFloat_fixed_0 <= r_sys_tmp204_int;

									end
									else
									if((r_sys_run_step==9'h2d)) begin
										r_ip_FixedToFloat_fixed_0 <= r_sys_tmp30_int;

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_ip_FixedToFloat_fixed_0 <= r_sys_tmp60_int;

									end
									else
									if((r_sys_run_step==9'h15) || (r_sys_run_step==9'h23)) begin
										r_ip_FixedToFloat_fixed_0 <= r_sys_tmp205_int;

									end
									else
									if((r_sys_run_step==9'ha) || (r_sys_run_step==9'hc) || (r_sys_run_step==9'he) || (r_sys_run_step==9'h10) || (r_sys_run_step==9'h12) || (r_sys_run_step==9'h14) || (r_sys_run_step==9'h16) || (r_sys_run_step==9'h18) || (r_sys_run_step==9'h1a) || (r_sys_run_step==9'h1c) || (r_sys_run_step==9'h1e) || (r_sys_run_step==9'h20) || (r_sys_run_step==9'h22) || (r_sys_run_step==9'h24) || (r_sys_run_step==9'h26) || (r_sys_run_step==9'h28) || (r_sys_run_step==9'h2a) || (r_sys_run_step==9'h2c) || (r_sys_run_step==9'h2e) || (r_sys_run_step==9'h30) || (r_sys_run_step==9'h32) || (r_sys_run_step==9'h34) || (9'h36<=r_sys_run_step && r_sys_run_step<=9'h3f)) begin
										r_ip_FixedToFloat_fixed_0 <= w_sys_tmp53;

									end
									else
									if((r_sys_run_step==9'h21)) begin
										r_ip_FixedToFloat_fixed_0 <= r_sys_tmp75_int;

									end
									else
									if((r_sys_run_step==9'h1d) || (r_sys_run_step==9'h33)) begin
										r_ip_FixedToFloat_fixed_0 <= r_sys_tmp203_int;

									end
									else
									if((r_sys_run_step==9'hd) || (r_sys_run_step==9'h13) || (r_sys_run_step==9'h1f)) begin
										r_ip_FixedToFloat_fixed_0 <= r_sys_tmp233_int;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_ip_fifo_under2up_in_0 <= w_sys_tmp2040;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_ip_fifo_under2up_s_we_0 <= w_sys_intOne;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_ip_fifo_under2up_s_re_0 <= r_sys_tmp4_int;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_ip_fifo_under2up_newData_0 <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_ip_fifo_up2under_in_0 <= w_sys_tmp2050;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_ip_fifo_up2under_s_we_0 <= r_run_s_up2under_we_12;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_ip_fifo_up2under_s_re_0 <= r_run_s_up2under_we_12;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_ip_fifo_up2under_newData_0 <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h26: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 6'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_phase <= 6'h2;
						end

						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'h4;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7) ? 6'h9 : 6'hf);

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'ha;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp12) ? 6'hd : 6'h6);

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h129)) begin
										r_sys_run_phase <= 6'ha;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'h10;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1708) ? 6'h14 : 6'h1a);

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'h10;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'h15;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1713) ? 6'h18 : 6'h11);

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h21)) begin
										r_sys_run_phase <= 6'h15;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'h1b;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2036) ? 6'h1e : 6'h20);

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_phase <= 6'h1b;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'h21;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2044) ? 6'h24 : 6'h26);

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_phase <= 6'h21;

									end
								end

							endcase
						end

						6'h26: begin
							r_sys_run_phase <= 6'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h129)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h21)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 9'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h128)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==9'h129)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h21)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h20)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						6'h26: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_addr_1 <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h87)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp92_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hc5)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp28_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h1e) || (r_sys_run_step==9'hdb)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp206_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hb1)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp51_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp141_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h57)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp144_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hac)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp54_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h6c)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp120_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h3a)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp173_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h31)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp178_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h9b)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp71_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp191_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h2a)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp183_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp154_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h7c)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp105_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hce)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp18_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hd6)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp11_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h49)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp155_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h55)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp142_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h76)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp111_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp169_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hd8)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp8_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hd) || (r_sys_run_step==9'h68)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp230_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h9d)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp73_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hb8)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp42_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h42)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp163_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h1c) || (r_sys_run_step==9'hcb)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp207_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h6b)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp124_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h6e)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp119_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h7b)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp107_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h95)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp79_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h66)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp125_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hb) || (r_sys_run_step==9'h58)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp229_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h96)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp77_int[13:0] );

									end
									else
									if((r_sys_run_step==9'ha0)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp68_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hbb)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp39_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h2) || (r_sys_run_step==9'h17) || (r_sys_run_step==9'haa)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp235_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hc) || (r_sys_run_step==9'h60)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp224_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h41)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp162_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hb7)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp41_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h64)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp131_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h14) || (r_sys_run_step==9'h99)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp215_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h8f)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp85_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h23)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp194_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hb0)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp50_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp153_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp149_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h22)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp195_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hbc)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp38_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h67)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp127_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h8a)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp91_int[13:0] );

									end
									else
									if((r_sys_run_step==9'he) || (r_sys_run_step==9'h69)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp220_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hbf)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp35_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h35)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp176_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hae)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp53_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h82)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp100_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h26)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp190_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h92)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp83_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h9f)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp70_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hcf)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp19_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h8b)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp90_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hdd)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp4_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h20)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp197_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h30)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp181_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h34)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp175_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h94)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp78_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hbd)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp33_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h53)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp146_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h33)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp180_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h44)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp161_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hb9)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp43_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h1d) || (r_sys_run_step==9'hd3)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp208_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h4f)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp150_int[13:0] );

									end
									else
									if((r_sys_run_step==9'ha6)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp63_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp170_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h2c)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp185_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp172_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h2d)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp186_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h5) || (r_sys_run_step==9'h2f)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp222_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h46)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp157_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h85)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp95_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h10) || (r_sys_run_step==9'h79)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp217_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h56)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp143_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h15) || (r_sys_run_step==9'h9a)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp213_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h11) || (r_sys_run_step==9'h81)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp218_int[13:0] );

									end
									else
									if((r_sys_run_step==9'ha5)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp62_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h62)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp129_int[13:0] );

									end
									else
									if((r_sys_run_step==9'haf)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp49_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h2e)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp182_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h36)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp174_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hc6)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp25_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hd4)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp14_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp159_int[13:0] );

									end
									else
									if((r_sys_run_step==9'ha1)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp67_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hb3)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp47_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h8e)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp84_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h90)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp86_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hda)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp7_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h61)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp132_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp192_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hc9)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp24_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h74)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp114_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h72)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp117_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hc0)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp36_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h4d)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp152_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h4a)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp156_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h1) || (r_sys_run_step==9'hf) || (r_sys_run_step==9'h71)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp234_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hc8)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp23_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h75)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp112_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h18) || (r_sys_run_step==9'hb2)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp214_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hb4)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp48_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hb5)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp46_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h45)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp160_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h86)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp96_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hc7)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp29_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h8) || (r_sys_run_step==9'h40)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp226_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h7f)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp103_int[13:0] );

									end
									else
									if((r_sys_run_step==9'ha) || (r_sys_run_step==9'h50)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp225_int[13:0] );

									end
									else
									if((r_sys_run_step==9'ha7)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp61_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h6) || (r_sys_run_step==9'h37)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp221_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h9e)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp69_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hb6)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp40_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h6a)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp123_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h5c)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp135_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h3f)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp166_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h43)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp164_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h8c)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp88_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h12) || (r_sys_run_step==9'h89)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp219_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h63)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp130_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h93)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp82_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h51)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp147_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hd2)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp13_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b) || (r_sys_run_step==9'hca)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp209_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h84)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp97_int[13:0] );

									end
									else
									if((r_sys_run_step==9'had)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp55_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hcc)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp21_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h5f)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp133_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hd1)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp16_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h19) || (r_sys_run_step==9'hba)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp210_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp168_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h7e)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp102_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h7) || (r_sys_run_step==9'h38)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp227_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hc4)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp27_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hab)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp57_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hcd)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp22_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h65)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp126_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h88)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp93_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hd0)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp17_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h77)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp109_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp20[13:0] );

									end
									else
									if((r_sys_run_step==9'hdc)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp3_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h3e)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp167_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hd9)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp6_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hbe)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp34_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a) || (r_sys_run_step==9'hc2)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp211_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h5e)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp137_int[13:0] );

									end
									else
									if((r_sys_run_step==9'ha3)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp64_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hd7)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp9_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hc3)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp31_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h80)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp99_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h83)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp98_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h29)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp188_int[13:0] );

									end
									else
									if((r_sys_run_step==9'ha9)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp56_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h70)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp116_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h9) || (r_sys_run_step==9'h48)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp228_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hd5)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp10_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp148_int[13:0] );

									end
									else
									if((r_sys_run_step==9'ha4)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp65_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h4) || (r_sys_run_step==9'h27)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp231_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h5b)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp134_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h3) || (r_sys_run_step==9'h1f)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp223_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h9c)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp72_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h6f)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp118_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hc1)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp32_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h78)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp110_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h16) || (r_sys_run_step==9'ha2)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp212_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hdf)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp1_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h13) || (r_sys_run_step==9'h91)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp216_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h59)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp140_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h2b)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp184_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h7d)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp104_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h28)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp189_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h5d)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp136_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h73)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp113_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h98)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp76_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h6d)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp121_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hde)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp2_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h32)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp179_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h97)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp80_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h7a)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp106_int[13:0] );

									end
									else
									if((r_sys_run_step==9'ha8)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp59_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h5a)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp139_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h21)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp196_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h8d)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp89_int[13:0] );

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h2) || (r_sys_run_step==9'h5) || (r_sys_run_step==9'h8) || (r_sys_run_step==9'hb) || (r_sys_run_step==9'he) || (r_sys_run_step==9'h11) || (r_sys_run_step==9'h14) || (r_sys_run_step==9'h17) || (r_sys_run_step==9'h1a) || (r_sys_run_step==9'h1d) || (r_sys_run_step==9'h20)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp1_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h4) || (r_sys_run_step==9'h7) || (r_sys_run_step==9'ha) || (r_sys_run_step==9'hd) || (r_sys_run_step==9'h10) || (r_sys_run_step==9'h13) || (r_sys_run_step==9'h16) || (r_sys_run_step==9'h19) || (r_sys_run_step==9'h1c) || (r_sys_run_step==9'h1f)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp0_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h3) || (r_sys_run_step==9'h6) || (r_sys_run_step==9'h9) || (r_sys_run_step==9'hc) || (r_sys_run_step==9'hf) || (r_sys_run_step==9'h12) || (r_sys_run_step==9'h15) || (r_sys_run_step==9'h18) || (r_sys_run_step==9'h1b) || (r_sys_run_step==9'h1e) || (r_sys_run_step==9'h21)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp2_int[13:0] );

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2041[13:0] );

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp5_int[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h21)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp1720;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp2049;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'hdf)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h21)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h26: begin
							r_fld_u_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_result_1_addr_1 <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hfc)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp115_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h128)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp12_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hf6)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp122_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h10b)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp94_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h110)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp87_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hba)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp171_int[13:0] );

									end
									else
									if((r_sys_run_step==9'ha7)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp187_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h80)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp200_int[13:0] );

									end
									else
									if((r_sys_run_step==9'he8)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp138_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h118)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp74_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h125)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp37_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h106)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp101_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h126)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp26_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h101)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp108_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hd8)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp151_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hb0)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp177_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h129)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp5_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hcd)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp158_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h9c)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp193_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hdf)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp145_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h76)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp201_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h124)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp44_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h11e)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp58_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h92)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp198_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h121)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp52_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hf0)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp128_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h11b)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp66_int[13:0] );

									end
									else
									if((r_sys_run_step==9'hc3)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp165_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h89)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp199_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h115)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp81_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h6b)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp202_int[13:0] );

									end
									else
									if((r_sys_run_step==9'h127)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp20_int[13:0] );

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_fld_result_1_addr_1 <= $signed( w_sys_tmp1721[13:0] );

									end
									else
									if((9'h1<=r_sys_run_step && r_sys_run_step<=9'h1f)) begin
										r_fld_result_1_addr_1 <= $signed( r_sys_tmp3_int[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h6b) || (r_sys_run_step==9'h76) || (r_sys_run_step==9'h80) || (r_sys_run_step==9'h89) || (r_sys_run_step==9'h92) || (r_sys_run_step==9'h9c) || (r_sys_run_step==9'ha7) || (r_sys_run_step==9'hb0) || (r_sys_run_step==9'hba) || (r_sys_run_step==9'hc3) || (r_sys_run_step==9'hcd) || (r_sys_run_step==9'hd8) || (r_sys_run_step==9'hdf) || (r_sys_run_step==9'he8) || (r_sys_run_step==9'hf0) || (r_sys_run_step==9'hf6) || (r_sys_run_step==9'hfc) || (r_sys_run_step==9'h101) || (r_sys_run_step==9'h106) || (r_sys_run_step==9'h10b) || (r_sys_run_step==9'h110) || (r_sys_run_step==9'h115) || (r_sys_run_step==9'h118) || (r_sys_run_step==9'h11b) || (r_sys_run_step==9'h11e) || (r_sys_run_step==9'h121) || (9'h124<=r_sys_run_step && r_sys_run_step<=9'h129)) begin
										r_fld_result_1_datain_1 <= w_sys_tmp19;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_result_1_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h6b) || (r_sys_run_step==9'h76) || (r_sys_run_step==9'h80) || (r_sys_run_step==9'h89) || (r_sys_run_step==9'h92) || (r_sys_run_step==9'h9c) || (r_sys_run_step==9'ha7) || (r_sys_run_step==9'hb0) || (r_sys_run_step==9'hba) || (r_sys_run_step==9'hc3) || (r_sys_run_step==9'hcd) || (r_sys_run_step==9'hd8) || (r_sys_run_step==9'hdf) || (r_sys_run_step==9'he8) || (r_sys_run_step==9'hf0) || (r_sys_run_step==9'hf6) || (r_sys_run_step==9'hfc) || (r_sys_run_step==9'h101) || (r_sys_run_step==9'h106) || (r_sys_run_step==9'h10b) || (r_sys_run_step==9'h110) || (r_sys_run_step==9'h115) || (r_sys_run_step==9'h118) || (r_sys_run_step==9'h11b) || (r_sys_run_step==9'h11e) || (r_sys_run_step==9'h121) || (9'h124<=r_sys_run_step && r_sys_run_step<=9'h129)) begin
										r_fld_result_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1f)) begin
										r_fld_result_1_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h26: begin
							r_fld_result_1_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_r1_2 <= w_sys_tmp2052;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_fld_r1_2 <= w_sys_tmp4;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_r2_3 <= w_sys_tmp2053;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_fld_r2_3 <= w_sys_tmp4;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_dx_4 <= w_sys_tmp2054;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_fld_dx_4 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_dy_5 <= w_sys_tmp2055;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_fld_dy_5 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_dt_6 <= w_sys_tmp2056;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_fld_dt_6 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_7 <= w_sys_tmp6;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_7 <= w_sys_tmp10;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_7 <= w_sys_tmp1707;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_7 <= w_sys_tmp1711;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_7 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_7 <= w_sys_tmp2043;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_7 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_7 <= w_sys_tmp2051;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_j_8 <= w_sys_tmp11;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1f)) begin
										r_run_j_8 <= w_sys_tmp62;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_j_8 <= w_sys_tmp1712;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1f)) begin
										r_run_j_8 <= w_sys_tmp1725;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_s_under2up_re_9 <= w_sys_intZero;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_s_under2up_re_9 <= w_sys_intZero;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_s_under2up_we_10 <= w_sys_intZero;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_s_under2up_we_10 <= w_sys_intOne;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_s_up2under_re_11 <= w_sys_intZero;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_s_up2under_re_11 <= w_sys_intOne;

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_run_s_up2under_re_11 <= w_sys_intZero;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_s_up2under_we_12 <= w_sys_intZero;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy0_j_19 <= r_run_j_8;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1f)) begin
										r_run_copy0_j_19 <= w_sys_tmp54;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy1_j_20 <= r_run_j_8;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1f)) begin
										r_run_copy1_j_20 <= w_sys_tmp55;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy2_j_21 <= r_run_j_8;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1f)) begin
										r_run_copy2_j_21 <= w_sys_tmp56;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy3_j_22 <= r_run_j_8;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1f)) begin
										r_run_copy3_j_22 <= w_sys_tmp57;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy4_j_23 <= r_run_j_8;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1f)) begin
										r_run_copy4_j_23 <= w_sys_tmp58;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy5_j_24 <= r_run_j_8;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1f)) begin
										r_run_copy5_j_24 <= w_sys_tmp59;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy6_j_25 <= r_run_j_8;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1f)) begin
										r_run_copy6_j_25 <= w_sys_tmp26;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy7_j_26 <= r_run_j_8;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1f)) begin
										r_run_copy7_j_26 <= w_sys_tmp61;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy0_j_27 <= r_run_j_8;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1f)) begin
										r_run_copy0_j_27 <= w_sys_tmp1724;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1e)) begin
										r_sys_tmp0_int <= w_sys_tmp2072;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1) || (r_sys_run_step==9'h4) || (r_sys_run_step==9'h7) || (r_sys_run_step==9'ha) || (r_sys_run_step==9'hd) || (r_sys_run_step==9'h10) || (r_sys_run_step==9'h13) || (r_sys_run_step==9'h16) || (r_sys_run_step==9'h19) || (r_sys_run_step==9'h1c)) begin
										r_sys_tmp0_int <= w_sys_tmp2344;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1e)) begin
										r_sys_tmp1_int <= w_sys_tmp2071;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_tmp1_int <= w_sys_tmp2343;

									end
									else
									if((r_sys_run_step==9'h2) || (r_sys_run_step==9'h5) || (r_sys_run_step==9'h8) || (r_sys_run_step==9'hb) || (r_sys_run_step==9'he) || (r_sys_run_step==9'h11) || (r_sys_run_step==9'h14) || (r_sys_run_step==9'h17) || (r_sys_run_step==9'h1a) || (r_sys_run_step==9'h1d)) begin
										r_sys_tmp1_int <= w_sys_tmp2344;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1e)) begin
										r_sys_tmp2_int <= w_sys_tmp2070;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0) || (r_sys_run_step==9'h3) || (r_sys_run_step==9'h6) || (r_sys_run_step==9'h9) || (r_sys_run_step==9'hc) || (r_sys_run_step==9'hf) || (r_sys_run_step==9'h12) || (r_sys_run_step==9'h15) || (r_sys_run_step==9'h18) || (r_sys_run_step==9'h1b) || (r_sys_run_step==9'h1e)) begin
										r_sys_tmp2_int <= w_sys_tmp2344;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1e)) begin
										r_sys_tmp3_int <= w_sys_tmp2068;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1e)) begin
										r_sys_tmp3_int <= w_sys_tmp2345;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1e)) begin
										r_sys_tmp4_int <= w_sys_tmp2069;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_tmp4_int <= r_run_s_under2up_re_9;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1e)) begin
										r_sys_tmp5_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_tmp5_int <= w_sys_tmp2406;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1e)) begin
										r_sys_tmp6_int <= w_sys_tmp2065;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1e)) begin
										r_sys_tmp7_int <= w_sys_tmp2066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1d)) begin
										r_sys_tmp8_int <= w_sys_tmp2071;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1d)) begin
										r_sys_tmp9_int <= w_sys_tmp2070;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1d)) begin
										r_sys_tmp10_int <= w_sys_tmp2068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1d)) begin
										r_sys_tmp11_int <= w_sys_tmp2069;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1d)) begin
										r_sys_tmp12_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1d)) begin
										r_sys_tmp13_int <= w_sys_tmp2065;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1d)) begin
										r_sys_tmp14_int <= w_sys_tmp2067;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1c)) begin
										r_sys_tmp15_int <= w_sys_tmp2072;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1c)) begin
										r_sys_tmp16_int <= w_sys_tmp2071;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1c)) begin
										r_sys_tmp17_int <= w_sys_tmp2070;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1c)) begin
										r_sys_tmp18_int <= w_sys_tmp2068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1c)) begin
										r_sys_tmp19_int <= w_sys_tmp2069;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1c)) begin
										r_sys_tmp20_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1c)) begin
										r_sys_tmp21_int <= w_sys_tmp2066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1c)) begin
										r_sys_tmp22_int <= w_sys_tmp2067;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sys_tmp23_int <= w_sys_tmp2069;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sys_tmp24_int <= w_sys_tmp2070;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sys_tmp25_int <= w_sys_tmp2067;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sys_tmp26_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sys_tmp27_int <= w_sys_tmp2065;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sys_tmp28_int <= w_sys_tmp2066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sys_tmp29_int <= w_sys_tmp2068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1a)) begin
										r_sys_tmp30_int <= w_sys_tmp2072;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1a)) begin
										r_sys_tmp31_int <= w_sys_tmp2071;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1a)) begin
										r_sys_tmp32_int <= w_sys_tmp2069;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1a)) begin
										r_sys_tmp33_int <= w_sys_tmp2065;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1a)) begin
										r_sys_tmp34_int <= w_sys_tmp2066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1a)) begin
										r_sys_tmp35_int <= w_sys_tmp2067;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1a)) begin
										r_sys_tmp36_int <= w_sys_tmp2068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1a)) begin
										r_sys_tmp37_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h19)) begin
										r_sys_tmp38_int <= w_sys_tmp2071;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h19)) begin
										r_sys_tmp39_int <= w_sys_tmp2070;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h19)) begin
										r_sys_tmp40_int <= w_sys_tmp2065;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h19)) begin
										r_sys_tmp41_int <= w_sys_tmp2066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h19)) begin
										r_sys_tmp42_int <= w_sys_tmp2067;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h19)) begin
										r_sys_tmp43_int <= w_sys_tmp2068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h19)) begin
										r_sys_tmp44_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_tmp45_int <= w_sys_tmp2072;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_tmp46_int <= w_sys_tmp2071;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_tmp47_int <= w_sys_tmp2069;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_tmp48_int <= w_sys_tmp2070;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_tmp49_int <= w_sys_tmp2065;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_tmp50_int <= w_sys_tmp2066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_tmp51_int <= w_sys_tmp2067;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_tmp52_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h17)) begin
										r_sys_tmp53_int <= w_sys_tmp2071;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h17)) begin
										r_sys_tmp54_int <= w_sys_tmp2069;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h17)) begin
										r_sys_tmp55_int <= w_sys_tmp2070;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h17)) begin
										r_sys_tmp56_int <= w_sys_tmp2066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h17)) begin
										r_sys_tmp57_int <= w_sys_tmp2068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h17)) begin
										r_sys_tmp58_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h17)) begin
										r_sys_tmp59_int <= w_sys_tmp2065;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h16)) begin
										r_sys_tmp60_int <= w_sys_tmp2072;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h16)) begin
										r_sys_tmp61_int <= w_sys_tmp2071;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h16)) begin
										r_sys_tmp62_int <= w_sys_tmp2069;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h16)) begin
										r_sys_tmp63_int <= w_sys_tmp2070;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h16)) begin
										r_sys_tmp64_int <= w_sys_tmp2067;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h16)) begin
										r_sys_tmp65_int <= w_sys_tmp2068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h16)) begin
										r_sys_tmp66_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h16)) begin
										r_sys_tmp67_int <= w_sys_tmp2065;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp68_int <= w_sys_tmp2071;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp69_int <= w_sys_tmp2069;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp70_int <= w_sys_tmp2070;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp71_int <= w_sys_tmp2066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp72_int <= w_sys_tmp2067;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp73_int <= w_sys_tmp2068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp74_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp75_int <= w_sys_tmp2072;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp76_int <= w_sys_tmp2070;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp77_int <= w_sys_tmp2068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp78_int <= w_sys_tmp2066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp79_int <= w_sys_tmp2067;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp80_int <= w_sys_tmp2069;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp81_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp82_int <= w_sys_tmp2065;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp83_int <= w_sys_tmp2071;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp84_int <= w_sys_tmp2067;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp85_int <= w_sys_tmp2068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp86_int <= w_sys_tmp2069;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp87_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp88_int <= w_sys_tmp2065;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp89_int <= w_sys_tmp2066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp90_int <= w_sys_tmp2071;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp91_int <= w_sys_tmp2070;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp92_int <= w_sys_tmp2067;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp93_int <= w_sys_tmp2068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp94_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp95_int <= w_sys_tmp2065;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp96_int <= w_sys_tmp2066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp97_int <= w_sys_tmp2071;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp98_int <= w_sys_tmp2070;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp99_int <= w_sys_tmp2067;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp100_int <= w_sys_tmp2069;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp101_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp102_int <= w_sys_tmp2065;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp103_int <= w_sys_tmp2066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp104_int <= w_sys_tmp2071;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp105_int <= w_sys_tmp2070;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp106_int <= w_sys_tmp2068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp107_int <= w_sys_tmp2069;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp108_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp109_int <= w_sys_tmp2065;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp110_int <= w_sys_tmp2066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp111_int <= w_sys_tmp2071;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp112_int <= w_sys_tmp2070;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp113_int <= w_sys_tmp2068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp114_int <= w_sys_tmp2069;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp115_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp116_int <= w_sys_tmp2065;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp117_int <= w_sys_tmp2067;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp118_int <= w_sys_tmp2071;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp119_int <= w_sys_tmp2070;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp120_int <= w_sys_tmp2068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp121_int <= w_sys_tmp2069;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp122_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp123_int <= w_sys_tmp2066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp124_int <= w_sys_tmp2067;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp125_int <= w_sys_tmp2069;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp126_int <= w_sys_tmp2068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp127_int <= w_sys_tmp2070;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp128_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp129_int <= w_sys_tmp2065;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp130_int <= w_sys_tmp2066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp131_int <= w_sys_tmp2067;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp132_int <= w_sys_tmp2071;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp133_int <= w_sys_tmp2069;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp134_int <= w_sys_tmp2065;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp135_int <= w_sys_tmp2066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp136_int <= w_sys_tmp2067;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp137_int <= w_sys_tmp2068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp138_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp139_int <= w_sys_tmp2071;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp140_int <= w_sys_tmp2070;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp141_int <= w_sys_tmp2065;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp142_int <= w_sys_tmp2066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp143_int <= w_sys_tmp2067;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp144_int <= w_sys_tmp2068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp145_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp146_int <= w_sys_tmp2071;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp147_int <= w_sys_tmp2069;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp148_int <= w_sys_tmp2070;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp149_int <= w_sys_tmp2066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp150_int <= w_sys_tmp2067;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp151_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp152_int <= w_sys_tmp2065;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp153_int <= w_sys_tmp2071;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp154_int <= w_sys_tmp2070;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp155_int <= w_sys_tmp2068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp156_int <= w_sys_tmp2069;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp157_int <= w_sys_tmp2065;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp158_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp159_int <= w_sys_tmp2066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp160_int <= w_sys_tmp2071;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp161_int <= w_sys_tmp2070;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp162_int <= w_sys_tmp2067;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp163_int <= w_sys_tmp2068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp164_int <= w_sys_tmp2069;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp165_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp166_int <= w_sys_tmp2065;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp167_int <= w_sys_tmp2071;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp168_int <= w_sys_tmp2070;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp169_int <= w_sys_tmp2068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp170_int <= w_sys_tmp2069;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp171_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp172_int <= w_sys_tmp2066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp173_int <= w_sys_tmp2067;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp174_int <= w_sys_tmp2070;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp175_int <= w_sys_tmp2068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp176_int <= w_sys_tmp2069;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp177_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp178_int <= w_sys_tmp2065;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp179_int <= w_sys_tmp2066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp180_int <= w_sys_tmp2067;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp181_int <= w_sys_tmp2071;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp182_int <= w_sys_tmp2069;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp183_int <= w_sys_tmp2065;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp184_int <= w_sys_tmp2066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp185_int <= w_sys_tmp2067;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp186_int <= w_sys_tmp2068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp187_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp188_int <= w_sys_tmp2071;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp189_int <= w_sys_tmp2070;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp190_int <= w_sys_tmp2068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp191_int <= w_sys_tmp2066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp192_int <= w_sys_tmp2067;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp193_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp194_int <= w_sys_tmp2065;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp195_int <= w_sys_tmp2071;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp196_int <= w_sys_tmp2070;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp197_int <= w_sys_tmp2069;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp198_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp199_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_tmp200_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_tmp201_int <= w_sys_tmp2064;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_tmp202_int <= w_sys_tmp2057;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h12) || (r_sys_run_step==9'h1d)) begin
										r_sys_tmp203_int <= w_sys_tmp2072;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h10) || (r_sys_run_step==9'h19)) begin
										r_sys_tmp204_int <= w_sys_tmp2072;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'he) || (r_sys_run_step==9'h15)) begin
										r_sys_tmp205_int <= w_sys_tmp2072;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h3) || (r_sys_run_step==9'h1e)) begin
										r_sys_tmp206_int <= w_sys_tmp2067;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h3) || (r_sys_run_step==9'h1c)) begin
										r_sys_tmp207_int <= w_sys_tmp2065;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h3) || (r_sys_run_step==9'h1d)) begin
										r_sys_tmp208_int <= w_sys_tmp2066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h2) || (r_sys_run_step==9'h1b)) begin
										r_sys_tmp209_int <= w_sys_tmp2071;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h2) || (r_sys_run_step==9'h19)) begin
										r_sys_tmp210_int <= w_sys_tmp2069;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h2) || (r_sys_run_step==9'h1a)) begin
										r_sys_tmp211_int <= w_sys_tmp2070;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h2) || (r_sys_run_step==9'h16)) begin
										r_sys_tmp212_int <= w_sys_tmp2066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h2) || (r_sys_run_step==9'h15)) begin
										r_sys_tmp213_int <= w_sys_tmp2065;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h2) || (r_sys_run_step==9'h18)) begin
										r_sys_tmp214_int <= w_sys_tmp2068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1) || (r_sys_run_step==9'h14)) begin
										r_sys_tmp215_int <= w_sys_tmp2071;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1) || (r_sys_run_step==9'h13)) begin
										r_sys_tmp216_int <= w_sys_tmp2070;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1) || (r_sys_run_step==9'h10)) begin
										r_sys_tmp217_int <= w_sys_tmp2067;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1) || (r_sys_run_step==9'h11)) begin
										r_sys_tmp218_int <= w_sys_tmp2068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1) || (r_sys_run_step==9'h12)) begin
										r_sys_tmp219_int <= w_sys_tmp2069;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1) || (r_sys_run_step==9'he)) begin
										r_sys_tmp220_int <= w_sys_tmp2065;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp221_int <= w_sys_tmp2071;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_tmp221_int <= w_sys_tmp2063;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp222_int <= w_sys_tmp2070;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_tmp222_int <= w_sys_tmp2062;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_tmp223_int <= w_sys_tmp2060;

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp223_int <= w_sys_tmp2068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0) || (r_sys_run_step==9'hc)) begin
										r_sys_tmp224_int <= w_sys_tmp2070;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0) || (r_sys_run_step==9'ha)) begin
										r_sys_tmp225_int <= w_sys_tmp2068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0) || (r_sys_run_step==9'h8)) begin
										r_sys_tmp226_int <= w_sys_tmp2066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0) || (r_sys_run_step==9'h7)) begin
										r_sys_tmp227_int <= w_sys_tmp2065;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0) || (r_sys_run_step==9'h9)) begin
										r_sys_tmp228_int <= w_sys_tmp2067;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0) || (r_sys_run_step==9'hb)) begin
										r_sys_tmp229_int <= w_sys_tmp2069;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0) || (r_sys_run_step==9'hd)) begin
										r_sys_tmp230_int <= w_sys_tmp2071;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp231_int <= w_sys_tmp2069;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_tmp231_int <= w_sys_tmp2061;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hc) || (r_sys_run_step==9'h11) || (r_sys_run_step==9'h1b)) begin
										r_sys_tmp232_int <= w_sys_tmp2072;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'ha) || (r_sys_run_step==9'hd) || (r_sys_run_step==9'h13)) begin
										r_sys_tmp233_int <= w_sys_tmp2072;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_tmp234_int <= w_sys_tmp2058;

									end
									else
									if((r_sys_run_step==9'h1) || (r_sys_run_step==9'hf)) begin
										r_sys_tmp234_int <= w_sys_tmp2066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h2) || (r_sys_run_step==9'h17)) begin
										r_sys_tmp235_int <= w_sys_tmp2067;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_tmp235_int <= w_sys_tmp2059;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h9) || (r_sys_run_step==9'hb) || (r_sys_run_step==9'hf) || (r_sys_run_step==9'h17)) begin
										r_sys_tmp236_int <= w_sys_tmp2072;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h46)) begin
										r_sys_tmp0_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h44)) begin
										r_sys_tmp1_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h43)) begin
										r_sys_tmp2_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h42)) begin
										r_sys_tmp3_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h41)) begin
										r_sys_tmp4_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h40)) begin
										r_sys_tmp5_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h3f)) begin
										r_sys_tmp6_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h3e)) begin
										r_sys_tmp7_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h3c)) begin
										r_sys_tmp8_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h3b)) begin
										r_sys_tmp9_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h3a)) begin
										r_sys_tmp10_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h39)) begin
										r_sys_tmp11_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h38)) begin
										r_sys_tmp12_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h37)) begin
										r_sys_tmp13_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h36)) begin
										r_sys_tmp14_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h35)) begin
										r_sys_tmp15_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h33)) begin
										r_sys_tmp16_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h32)) begin
										r_sys_tmp17_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h31)) begin
										r_sys_tmp18_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h30)) begin
										r_sys_tmp19_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h2f)) begin
										r_sys_tmp20_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h2e)) begin
										r_sys_tmp21_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h2c)) begin
										r_sys_tmp22_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h2b)) begin
										r_sys_tmp23_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h2a)) begin
										r_sys_tmp24_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h29)) begin
										r_sys_tmp25_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h26)) begin
										r_sys_tmp26_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h25)) begin
										r_sys_tmp27_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h23)) begin
										r_sys_tmp28_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h21)) begin
										r_sys_tmp29_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1f)) begin
										r_sys_tmp30_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h19)) begin
										r_sys_tmp31_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_tmp32_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp33_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp34_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'he) || (r_sys_run_step==9'h45)) begin
										r_sys_tmp35_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hd) || (r_sys_run_step==9'h3d)) begin
										r_sys_tmp36_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hc) || (r_sys_run_step==9'h34)) begin
										r_sys_tmp37_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hb) || (r_sys_run_step==9'h2d)) begin
										r_sys_tmp38_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hd1)) begin
										r_sys_tmp39_float <= w_ip_AddFloat_result_0;

									end
									else
									if((r_sys_run_step==9'h27)) begin
										r_sys_tmp39_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hb7)) begin
										r_sys_tmp40_float <= w_ip_AddFloat_result_0;

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_sys_tmp40_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h5a) || (r_sys_run_step==9'h8c) || (r_sys_run_step==9'hbd)) begin
										r_sys_tmp41_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h9f) || (r_sys_run_step==9'hc6)) begin
										r_sys_tmp42_float <= w_ip_AddFloat_result_0;

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_sys_tmp42_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h5a) || (r_sys_run_step==9'h7f) || (r_sys_run_step==9'hbe) || (r_sys_run_step==9'hee)) begin
										r_sys_tmp43_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h4d) || (r_sys_run_step==9'h54) || (r_sys_run_step==9'h82) || (r_sys_run_step==9'hb3)) begin
										r_sys_tmp44_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h45) || (r_sys_run_step==9'h72) || (r_sys_run_step==9'ha2) || (r_sys_run_step==9'heb)) begin
										r_sys_tmp45_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h42) || (r_sys_run_step==9'h6a) || (r_sys_run_step==9'h9e) || (r_sys_run_step==9'hcf)) begin
										r_sys_tmp46_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h32) || (r_sys_run_step==9'h58) || (r_sys_run_step==9'h8b) || (r_sys_run_step==9'hbc)) begin
										r_sys_tmp47_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'ha4) || (r_sys_run_step==9'ha6) || (r_sys_run_step==9'hcf)) begin
										r_sys_tmp48_float <= w_ip_AddFloat_result_0;

									end
									else
									if((r_sys_run_step==9'h20)) begin
										r_sys_tmp48_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'ha0) || (r_sys_run_step==9'ha7) || (r_sys_run_step==9'hb1)) begin
										r_sys_tmp49_float <= w_fld_u_0_dataout_1;

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_sys_tmp49_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h86) || (r_sys_run_step==9'hc9) || (r_sys_run_step==9'hef)) begin
										r_sys_tmp50_float <= w_ip_AddFloat_result_0;

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_sys_tmp50_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h75) || (r_sys_run_step==9'h8b) || (r_sys_run_step==9'hb1)) begin
										r_sys_tmp51_float <= w_ip_AddFloat_result_0;

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sys_tmp51_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h6a) || (r_sys_run_step==9'ha0) || (r_sys_run_step==9'hd3)) begin
										r_sys_tmp52_float <= w_ip_AddFloat_result_0;

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp52_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h61) || (r_sys_run_step==9'h8e) || (r_sys_run_step==9'hbf)) begin
										r_sys_tmp53_float <= w_ip_AddFloat_result_0;

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp53_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hc0) || (r_sys_run_step==9'hc2)) begin
										r_sys_tmp54_float <= w_ip_AddFloat_result_0;

									end
									else
									if((r_sys_run_step==9'h9) || (r_sys_run_step==9'h22)) begin
										r_sys_tmp54_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h55) || (r_sys_run_step==9'h83) || (r_sys_run_step==9'h9e) || (r_sys_run_step==9'hc5) || (r_sys_run_step==9'hec)) begin
										r_sys_tmp55_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h2e) || (r_sys_run_step==9'h47) || (r_sys_run_step==9'h71) || (r_sys_run_step==9'haa) || (r_sys_run_step==9'hed)) begin
										r_sys_tmp56_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h27) || (r_sys_run_step==9'h4a) || (r_sys_run_step==9'h74) || (r_sys_run_step==9'ha8) || (r_sys_run_step==9'hd8)) begin
										r_sys_tmp57_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h91) || (r_sys_run_step==9'hb3) || (r_sys_run_step==9'hdc) || (r_sys_run_step==9'he5)) begin
										r_sys_tmp58_float <= w_ip_AddFloat_result_0;

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sys_tmp58_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hd1) || (r_sys_run_step==9'hd7) || (r_sys_run_step==9'he1)) begin
										r_sys_tmp59_float <= w_fld_u_0_dataout_1;

									end
									else
									if((r_sys_run_step==9'ha) || (r_sys_run_step==9'h28)) begin
										r_sys_tmp59_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h4b) || (r_sys_run_step==9'h53) || (r_sys_run_step==9'h79) || (r_sys_run_step==9'h9b) || (r_sys_run_step==9'he2) || (r_sys_run_step==9'h103)) begin
										r_sys_tmp60_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h43) || (r_sys_run_step==9'h6c) || (r_sys_run_step==9'h6d) || (r_sys_run_step==9'ha0) || (r_sys_run_step==9'hd2) || (r_sys_run_step==9'hd9)) begin
										r_sys_tmp61_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h36) || (r_sys_run_step==9'h3c) || (r_sys_run_step==9'h68) || (r_sys_run_step==9'h98) || (r_sys_run_step==9'hbb) || (r_sys_run_step==9'he4)) begin
										r_sys_tmp62_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h31) || (r_sys_run_step==9'h57) || (r_sys_run_step==9'h85) || (r_sys_run_step==9'h86) || (r_sys_run_step==9'hb6) || (r_sys_run_step==9'hba)) begin
										r_sys_tmp63_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1c) || (r_sys_run_step==9'h39) || (r_sys_run_step==9'h62) || (r_sys_run_step==9'h96) || (r_sys_run_step==9'hc7) || (r_sys_run_step==9'hf0)) begin
										r_sys_tmp64_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h3d) || (r_sys_run_step==9'h41) || (r_sys_run_step==9'h64) || (r_sys_run_step==9'h8a) || (r_sys_run_step==9'had) || (r_sys_run_step==9'hd7) || (r_sys_run_step==9'h102)) begin
										r_sys_tmp65_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h2b) || (r_sys_run_step==9'h4e) || (r_sys_run_step==9'h7a) || (r_sys_run_step==9'h7b) || (r_sys_run_step==9'h81) || (r_sys_run_step==9'hb2) || (r_sys_run_step==9'he1)) begin
										r_sys_tmp66_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h20) || (r_sys_run_step==9'h3f) || (r_sys_run_step==9'h40) || (r_sys_run_step==9'h69) || (r_sys_run_step==9'h9a) || (r_sys_run_step==9'hce) || (r_sys_run_step==9'hf6)) begin
										r_sys_tmp67_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h19) || (r_sys_run_step==9'h38) || (r_sys_run_step==9'h5e) || (r_sys_run_step==9'h5f) || (r_sys_run_step==9'h94) || (r_sys_run_step==9'hc5) || (r_sys_run_step==9'hed)) begin
										r_sys_tmp68_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h4e) || (r_sys_run_step==9'h7c) || (r_sys_run_step==9'h95) || (r_sys_run_step==9'hb9) || (r_sys_run_step==9'hbc) || (r_sys_run_step==9'hdd)) begin
										r_sys_tmp69_float <= w_ip_AddFloat_result_0;

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp69_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h33) || (r_sys_run_step==9'h52) || (r_sys_run_step==9'h59) || (r_sys_run_step==9'h63) || (r_sys_run_step==9'h97) || (r_sys_run_step==9'hc8) || (r_sys_run_step==9'hf1) || (r_sys_run_step==9'h10d)) begin
										r_sys_tmp70_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h2b) || (r_sys_run_step==9'h4c) || (r_sys_run_step==9'h7b) || (r_sys_run_step==9'hab) || (r_sys_run_step==9'hac) || (r_sys_run_step==9'hdb) || (r_sys_run_step==9'hfe) || (r_sys_run_step==9'h112)) begin
										r_sys_tmp71_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1d) || (r_sys_run_step==9'h3a) || (r_sys_run_step==9'h5c) || (r_sys_run_step==9'h8d) || (r_sys_run_step==9'hd0) || (r_sys_run_step==9'hf7) || (r_sys_run_step==9'h111) || (r_sys_run_step==9'h11f)) begin
										r_sys_tmp72_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h6f) || (r_sys_run_step==9'h76) || (r_sys_run_step==9'h7c) || (r_sys_run_step==9'h8a) || (r_sys_run_step==9'h94) || (r_sys_run_step==9'h9d) || (r_sys_run_step==9'ha3)) begin
										r_sys_tmp73_float <= w_fld_u_0_dataout_1;

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp73_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hd5) || (r_sys_run_step==9'hde)) begin
										r_sys_tmp74_float <= w_ip_AddFloat_result_0;

									end
									else
									if((r_sys_run_step==9'h5b) || (r_sys_run_step==9'h70) || (r_sys_run_step==9'h71) || (r_sys_run_step==9'h78) || (r_sys_run_step==9'ha9)) begin
										r_sys_tmp74_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp74_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h28) || (r_sys_run_step==9'h29) || (r_sys_run_step==9'h40) || (r_sys_run_step==9'h67) || (r_sys_run_step==9'h78) || (r_sys_run_step==9'hb4) || (r_sys_run_step==9'he1) || (r_sys_run_step==9'hf8) || (r_sys_run_step==9'h10c)) begin
										r_sys_tmp75_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h22) || (r_sys_run_step==9'h39) || (r_sys_run_step==9'h60) || (r_sys_run_step==9'h6e) || (r_sys_run_step==9'h82) || (r_sys_run_step==9'ha9) || (r_sys_run_step==9'hcc) || (r_sys_run_step==9'h108) || (r_sys_run_step==9'h11c)) begin
										r_sys_tmp76_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h16) || (r_sys_run_step==9'h32) || (r_sys_run_step==9'h56) || (r_sys_run_step==9'h84) || (r_sys_run_step==9'hb5) || (r_sys_run_step==9'he3) || (r_sys_run_step==9'he9) || (r_sys_run_step==9'hfd) || (r_sys_run_step==9'h116)) begin
										r_sys_tmp77_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hf) || (r_sys_run_step==9'h1f) || (r_sys_run_step==9'h3b) || (r_sys_run_step==9'h61) || (r_sys_run_step==9'h8f) || (r_sys_run_step==9'h90) || (r_sys_run_step==9'hc4) || (r_sys_run_step==9'hea) || (r_sys_run_step==9'h104)) begin
										r_sys_tmp78_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hab) || (r_sys_run_step==9'hb5) || (r_sys_run_step==9'hbc) || (r_sys_run_step==9'hc3) || (r_sys_run_step==9'hc9) || (r_sys_run_step==9'hd3) || (r_sys_run_step==9'hdf)) begin
										r_sys_tmp79_float <= w_fld_u_0_dataout_1;

									end
									else
									if((r_sys_run_step==9'h8) || (r_sys_run_step==9'h1d)) begin
										r_sys_tmp79_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h12) || (r_sys_run_step==9'h23) || (r_sys_run_step==9'h24) || (r_sys_run_step==9'h49) || (r_sys_run_step==9'h73) || (r_sys_run_step==9'ha2) || (r_sys_run_step==9'ha4) || (r_sys_run_step==9'hd1) || (r_sys_run_step==9'hf4) || (r_sys_run_step==9'h109)) begin
										r_sys_tmp80_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h15) || (r_sys_run_step==9'h2a) || (r_sys_run_step==9'h4c) || (r_sys_run_step==9'h77) || (r_sys_run_step==9'ha5) || (r_sys_run_step==9'ha7) || (r_sys_run_step==9'hd3) || (r_sys_run_step==9'hd5) || (r_sys_run_step==9'hd6) || (r_sys_run_step==9'hf5) || (r_sys_run_step==9'h10a)) begin
										r_sys_tmp81_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'he) || (r_sys_run_step==9'h1b) || (r_sys_run_step==9'h34) || (r_sys_run_step==9'h35) || (r_sys_run_step==9'h5c) || (r_sys_run_step==9'h88) || (r_sys_run_step==9'h89) || (r_sys_run_step==9'hb7) || (r_sys_run_step==9'he7) || (r_sys_run_step==9'hff) || (r_sys_run_step==9'h118)) begin
										r_sys_tmp82_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hb) || (r_sys_run_step==9'h16) || (r_sys_run_step==9'h30) || (r_sys_run_step==9'h53) || (r_sys_run_step==9'h7e) || (r_sys_run_step==9'h7f) || (r_sys_run_step==9'haf) || (r_sys_run_step==9'hb0) || (r_sys_run_step==9'he0) || (r_sys_run_step==9'hfb) || (r_sys_run_step==9'h10f)) begin
										r_sys_tmp83_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h7) || (r_sys_run_step==9'hd) || (r_sys_run_step==9'h18) || (r_sys_run_step==9'h2d) || (r_sys_run_step==9'h50) || (r_sys_run_step==9'h7d) || (r_sys_run_step==9'hac) || (r_sys_run_step==9'hae) || (r_sys_run_step==9'hdf) || (r_sys_run_step==9'hfa) || (r_sys_run_step==9'h10e)) begin
										r_sys_tmp84_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h6) || (r_sys_run_step==9'ha) || (r_sys_run_step==9'h14) || (r_sys_run_step==9'h26) || (r_sys_run_step==9'h46) || (r_sys_run_step==9'h6f) || (r_sys_run_step==9'h9d) || (r_sys_run_step==9'hcb) || (r_sys_run_step==9'hef) || (r_sys_run_step==9'h105) || (r_sys_run_step==9'h115)) begin
										r_sys_tmp85_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h84) || (r_sys_run_step==9'h8b) || (r_sys_run_step==9'h92) || (r_sys_run_step==9'h98) || (r_sys_run_step==9'ha2) || (r_sys_run_step==9'had) || (r_sys_run_step==9'hb9) || (r_sys_run_step==9'hbf)) begin
										r_sys_tmp86_float <= w_fld_u_0_dataout_1;

									end
									else
									if((r_sys_run_step==9'ha1)) begin
										r_sys_tmp86_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==9'h7) || (r_sys_run_step==9'h17)) begin
										r_sys_tmp86_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'hd) || (r_sys_run_step==9'h13) || (r_sys_run_step==9'h21) || (r_sys_run_step==9'h2b) || (r_sys_run_step==9'h34) || (r_sys_run_step==9'h3a) || (r_sys_run_step==9'h59) || (r_sys_run_step==9'h63) || (r_sys_run_step==9'h6c) || (r_sys_run_step==9'h72) || (r_sys_run_step==9'ha4) || (r_sys_run_step==9'haa)) begin
										r_sys_tmp87_float <= w_fld_u_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h13) || (r_sys_run_step==9'h1a) || (r_sys_run_step==9'h21) || (r_sys_run_step==9'h24) || (r_sys_run_step==9'h44) || (r_sys_run_step==9'h4a) || (r_sys_run_step==9'h6d) || (r_sys_run_step==9'h94) || (r_sys_run_step==9'hda) || (r_sys_run_step==9'hf3) || (r_sys_run_step==9'h107) || (r_sys_run_step==9'h119) || (r_sys_run_step==9'h122)) begin
										r_sys_tmp88_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h5) || (r_sys_run_step==9'h8) || (r_sys_run_step==9'h11) || (r_sys_run_step==9'h22) || (r_sys_run_step==9'h3e) || (r_sys_run_step==9'h65) || (r_sys_run_step==9'h93) || (r_sys_run_step==9'hc1) || (r_sys_run_step==9'he8) || (r_sys_run_step==9'h100) || (r_sys_run_step==9'h112) || (r_sys_run_step==9'h11b) || (r_sys_run_step==9'h11e)) begin
										r_sys_tmp89_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h3) || (r_sys_run_step==9'h9) || (r_sys_run_step==9'h24) || (r_sys_run_step==9'h2d) || (r_sys_run_step==9'h33) || (r_sys_run_step==9'h4e) || (r_sys_run_step==9'h57) || (r_sys_run_step==9'h5d) || (r_sys_run_step==9'h86) || (r_sys_run_step==9'h8f) || (r_sys_run_step==9'h95) || (r_sys_run_step==9'hd5) || (r_sys_run_step==9'hdb)) begin
										r_sys_tmp90_float <= w_fld_u_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h8) || (r_sys_run_step==9'h11) || (r_sys_run_step==9'h17) || (r_sys_run_step==9'h2f) || (r_sys_run_step==9'h39) || (r_sys_run_step==9'h42) || (r_sys_run_step==9'h48) || (r_sys_run_step==9'h68) || (r_sys_run_step==9'h6e) || (r_sys_run_step==9'h78) || (r_sys_run_step==9'h81) || (r_sys_run_step==9'h87) || (r_sys_run_step==9'hc0) || (r_sys_run_step==9'hc6)) begin
										r_sys_tmp91_float <= w_fld_u_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h1b) || (r_sys_run_step==9'h22) || (r_sys_run_step==9'h4c) || (r_sys_run_step==9'h53) || (r_sys_run_step==9'h5a) || (r_sys_run_step==9'h61) || (r_sys_run_step==9'h67) || (r_sys_run_step==9'h71) || (r_sys_run_step==9'h7a) || (r_sys_run_step==9'h80) || (r_sys_run_step==9'hb7) || (r_sys_run_step==9'hc2) || (r_sys_run_step==9'hcc) || (r_sys_run_step==9'hd8) || (r_sys_run_step==9'hde)) begin
										r_sys_tmp92_float <= w_fld_u_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h14) || (r_sys_run_step==9'h1a) || (r_sys_run_step==9'h28) || (r_sys_run_step==9'h32) || (r_sys_run_step==9'h3b) || (r_sys_run_step==9'h41) || (r_sys_run_step==9'h60) || (r_sys_run_step==9'h6a) || (r_sys_run_step==9'h73) || (r_sys_run_step==9'h79) || (r_sys_run_step==9'hae) || (r_sys_run_step==9'hb4) || (r_sys_run_step==9'hbe) || (r_sys_run_step==9'hc7) || (r_sys_run_step==9'hcd)) begin
										r_sys_tmp93_float <= w_fld_u_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h6) || (r_sys_run_step==9'hc) || (r_sys_run_step==9'h16) || (r_sys_run_step==9'h1f) || (r_sys_run_step==9'h25) || (r_sys_run_step==9'h3d) || (r_sys_run_step==9'h47) || (r_sys_run_step==9'h50) || (r_sys_run_step==9'h56) || (r_sys_run_step==9'h7d) || (r_sys_run_step==9'h83) || (r_sys_run_step==9'h8d) || (r_sys_run_step==9'h96) || (r_sys_run_step==9'h9c) || (r_sys_run_step==9'hdc)) begin
										r_sys_tmp94_float <= w_fld_u_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h5) || (r_sys_run_step==9'hf) || (r_sys_run_step==9'h18) || (r_sys_run_step==9'h1e) || (r_sys_run_step==9'h36) || (r_sys_run_step==9'h40) || (r_sys_run_step==9'h49) || (r_sys_run_step==9'h4f) || (r_sys_run_step==9'h75) || (r_sys_run_step==9'h7f) || (r_sys_run_step==9'h88) || (r_sys_run_step==9'h8e) || (r_sys_run_step==9'hca) || (r_sys_run_step==9'hd0) || (r_sys_run_step==9'hda)) begin
										r_sys_tmp95_float <= w_fld_u_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'ha) || (r_sys_run_step==9'h10) || (r_sys_run_step==9'h29) || (r_sys_run_step==9'h30) || (r_sys_run_step==9'h37) || (r_sys_run_step==9'h3e) || (r_sys_run_step==9'h44) || (r_sys_run_step==9'h52) || (r_sys_run_step==9'h5c) || (r_sys_run_step==9'h65) || (r_sys_run_step==9'h6b) || (r_sys_run_step==9'h99) || (r_sys_run_step==9'h9f) || (r_sys_run_step==9'ha9) || (r_sys_run_step==9'hb2) || (r_sys_run_step==9'hb8)) begin
										r_sys_tmp96_float <= w_fld_u_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==9'h2) || (r_sys_run_step==9'h1d) || (r_sys_run_step==9'h26) || (r_sys_run_step==9'h2c) || (r_sys_run_step==9'h45) || (r_sys_run_step==9'h4b) || (r_sys_run_step==9'h55) || (r_sys_run_step==9'h5e) || (r_sys_run_step==9'h64) || (r_sys_run_step==9'h91) || (r_sys_run_step==9'h9b) || (r_sys_run_step==9'ha6) || (r_sys_run_step==9'hb0) || (r_sys_run_step==9'hbb) || (r_sys_run_step==9'hc5) || (r_sys_run_step==9'hce) || (r_sys_run_step==9'hd4)) begin
										r_sys_tmp97_float <= w_fld_u_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
