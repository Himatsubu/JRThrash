/*
TimeStamp:	2016/5/26		10:6
*/


module P3_unroll_small(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy	
);

	reg  signed [31:0] r_ip_DivInt_dividend_0;
	reg  signed [31:0] r_ip_DivInt_divisor_0;
	wire signed [31:0] w_ip_DivInt_quotient_0;
	wire signed [31:0] w_ip_DivInt_fractional_0;
	reg  signed [31:0] r_ip_DivInt_dividend_1;
	reg  signed [31:0] r_ip_DivInt_divisor_1;
	wire signed [31:0] w_ip_DivInt_quotient_1;
	wire signed [31:0] w_ip_DivInt_fractional_1;
	reg         [31:0] r_ip_AddFloat_portA_0;
	reg         [31:0] r_ip_AddFloat_portB_0;
	wire        [31:0] w_ip_AddFloat_result_0;
	reg         [31:0] r_ip_MultFloat_multiplicand_0;
	reg         [31:0] r_ip_MultFloat_multiplier_0;
	wire        [31:0] w_ip_MultFloat_product_0;
	reg  signed [31:0] r_ip_FixedToFloat_fixed_0;
	wire        [31:0] w_ip_FixedToFloat_floating_0;
	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 5:0] r_sys_run_phase;
	reg         [ 1:0] r_sys_run_stage;
	reg         [ 7:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 1:0] w_sys_run_stage_p1;
	wire        [ 7:0] w_sys_run_step_p1;
	wire signed [ 9:0] w_fld_T_0_addr_0;
	wire        [31:0] w_fld_T_0_datain_0;
	wire        [31:0] w_fld_T_0_dataout_0;
	wire               w_fld_T_0_r_w_0;
	wire               w_fld_T_0_ce_0;
	reg  signed [ 9:0] r_fld_T_0_addr_1;
	reg         [31:0] r_fld_T_0_datain_1;
	wire        [31:0] w_fld_T_0_dataout_1;
	reg                r_fld_T_0_r_w_1;
	wire               w_fld_T_0_ce_1;
	wire signed [ 9:0] w_fld_TT_1_addr_0;
	wire        [31:0] w_fld_TT_1_datain_0;
	wire        [31:0] w_fld_TT_1_dataout_0;
	wire               w_fld_TT_1_r_w_0;
	wire               w_fld_TT_1_ce_0;
	reg  signed [ 9:0] r_fld_TT_1_addr_1;
	reg         [31:0] r_fld_TT_1_datain_1;
	wire        [31:0] w_fld_TT_1_dataout_1;
	reg                r_fld_TT_1_r_w_1;
	wire               w_fld_TT_1_ce_1;
	wire signed [ 9:0] w_fld_U_2_addr_0;
	wire        [31:0] w_fld_U_2_datain_0;
	wire        [31:0] w_fld_U_2_dataout_0;
	wire               w_fld_U_2_r_w_0;
	wire               w_fld_U_2_ce_0;
	reg  signed [ 9:0] r_fld_U_2_addr_1;
	reg         [31:0] r_fld_U_2_datain_1;
	wire        [31:0] w_fld_U_2_dataout_1;
	reg                r_fld_U_2_r_w_1;
	wire               w_fld_U_2_ce_1;
	wire signed [ 9:0] w_fld_V_3_addr_0;
	wire        [31:0] w_fld_V_3_datain_0;
	wire        [31:0] w_fld_V_3_dataout_0;
	wire               w_fld_V_3_r_w_0;
	wire               w_fld_V_3_ce_0;
	reg  signed [ 9:0] r_fld_V_3_addr_1;
	reg         [31:0] r_fld_V_3_datain_1;
	wire        [31:0] w_fld_V_3_dataout_1;
	reg                r_fld_V_3_r_w_1;
	wire               w_fld_V_3_ce_1;
	reg  signed [31:0] r_run_k_4;
	reg  signed [31:0] r_run_j_5;
	reg  signed [31:0] r_run_n_6;
	reg  signed [31:0] r_run_mx_7;
	reg  signed [31:0] r_run_my_8;
	reg         [31:0] r_run_dt_9;
	reg         [31:0] r_run_dx_10;
	reg         [31:0] r_run_dy_11;
	reg         [31:0] r_run_r1_12;
	reg         [31:0] r_run_r2_13;
	reg         [31:0] r_run_r3_14;
	reg         [31:0] r_run_r4_15;
	reg         [31:0] r_run_YY_16;
	reg  signed [31:0] r_run_kx_17;
	reg  signed [31:0] r_run_ky_18;
	reg  signed [31:0] r_run_nlast_19;
	reg  signed [31:0] r_run_copy0_j_20;
	reg  signed [31:0] r_run_copy1_j_21;
	reg  signed [31:0] r_run_copy2_j_22;
	reg  signed [31:0] r_run_copy0_j_23;
	reg  signed [31:0] r_run_copy0_j_24;
	reg  signed [31:0] r_run_copy1_j_25;
	reg  signed [31:0] r_run_copy2_j_26;
	reg  signed [31:0] r_run_copy3_j_27;
	reg  signed [31:0] r_run_copy4_j_28;
	reg  signed [31:0] r_run_copy5_j_29;
	reg  signed [31:0] r_run_copy6_j_30;
	reg  signed [31:0] r_run_copy7_j_31;
	reg  signed [31:0] r_run_copy8_j_32;
	reg  signed [31:0] r_run_copy9_j_33;
	reg  signed [31:0] r_run_copy10_j_34;
	reg  signed [31:0] r_run_copy11_j_35;
	reg  signed [31:0] r_run_copy12_j_36;
	reg  signed [31:0] r_run_copy0_j_37;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg         [31:0] r_sys_tmp4_float;
	reg         [31:0] r_sys_tmp5_float;
	reg         [31:0] r_sys_tmp6_float;
	reg         [31:0] r_sys_tmp7_float;
	reg         [31:0] r_sys_tmp8_float;
	reg         [31:0] r_sys_tmp9_float;
	reg         [31:0] r_sys_tmp10_float;
	reg         [31:0] r_sys_tmp11_float;
	reg         [31:0] r_sys_tmp12_float;
	reg         [31:0] r_sys_tmp13_float;
	reg         [31:0] r_sys_tmp14_float;
	reg         [31:0] r_sys_tmp15_float;
	reg         [31:0] r_sys_tmp16_float;
	reg         [31:0] r_sys_tmp17_float;
	reg         [31:0] r_sys_tmp18_float;
	reg         [31:0] r_sys_tmp19_float;
	reg         [31:0] r_sys_tmp20_float;
	reg         [31:0] r_sys_tmp21_float;
	reg         [31:0] r_sys_tmp22_float;
	reg         [31:0] r_sys_tmp23_float;
	reg         [31:0] r_sys_tmp24_float;
	reg         [31:0] r_sys_tmp25_float;
	reg         [31:0] r_sys_tmp26_float;
	reg         [31:0] r_sys_tmp27_float;
	reg         [31:0] r_sys_tmp28_float;
	reg         [31:0] r_sys_tmp29_float;
	reg         [31:0] r_sys_tmp30_float;
	reg         [31:0] r_sys_tmp31_float;
	reg         [31:0] r_sys_tmp32_float;
	reg         [31:0] r_sys_tmp33_float;
	reg         [31:0] r_sys_tmp34_float;
	reg         [31:0] r_sys_tmp35_float;
	reg         [31:0] r_sys_tmp36_float;
	reg         [31:0] r_sys_tmp37_float;
	reg         [31:0] r_sys_tmp38_float;
	reg         [31:0] r_sys_tmp39_float;
	reg         [31:0] r_sys_tmp40_float;
	reg         [31:0] r_sys_tmp41_float;
	reg         [31:0] r_sys_tmp42_float;
	reg         [31:0] r_sys_tmp43_float;
	reg         [31:0] r_sys_tmp44_float;
	wire signed [31:0] w_sys_tmp1;
	wire signed [31:0] w_sys_tmp3;
	wire        [31:0] w_sys_tmp5;
	wire        [31:0] w_sys_tmp6;
	wire        [31:0] w_sys_tmp7;
	wire        [31:0] w_sys_tmp8;
	wire        [31:0] w_sys_tmp9;
	wire        [31:0] w_sys_tmp10;
	wire        [31:0] w_sys_tmp11;
	wire               w_sys_tmp12;
	wire               w_sys_tmp13;
	wire signed [31:0] w_sys_tmp14;
	wire               w_sys_tmp15;
	wire               w_sys_tmp16;
	wire        [31:0] w_sys_tmp18;
	wire        [31:0] w_sys_tmp19;
	wire signed [31:0] w_sys_tmp20;
	wire signed [31:0] w_sys_tmp22;
	wire signed [31:0] w_sys_tmp23;
	wire signed [31:0] w_sys_tmp24;
	wire        [31:0] w_sys_tmp25;
	wire signed [31:0] w_sys_tmp27;
	wire signed [31:0] w_sys_tmp28;
	wire signed [31:0] w_sys_tmp32;
	wire signed [31:0] w_sys_tmp33;
	wire        [31:0] w_sys_tmp36;
	wire        [31:0] w_sys_tmp37;
	wire        [31:0] w_sys_tmp38;
	wire signed [31:0] w_sys_tmp41;
	wire signed [31:0] w_sys_tmp42;
	wire signed [31:0] w_sys_tmp45;
	wire signed [31:0] w_sys_tmp46;
	wire signed [31:0] w_sys_tmp47;
	wire signed [31:0] w_sys_tmp48;
	wire        [31:0] w_sys_tmp128;
	wire        [31:0] w_sys_tmp157;
	wire        [31:0] w_sys_tmp185;
	wire        [31:0] w_sys_tmp213;
	wire        [31:0] w_sys_tmp269;
	wire        [31:0] w_sys_tmp297;
	wire               w_sys_tmp560;
	wire               w_sys_tmp561;
	wire signed [31:0] w_sys_tmp562;
	wire               w_sys_tmp563;
	wire               w_sys_tmp564;
	wire signed [31:0] w_sys_tmp567;
	wire signed [31:0] w_sys_tmp568;
	wire        [31:0] w_sys_tmp569;
	wire signed [31:0] w_sys_tmp571;
	wire signed [31:0] w_sys_tmp572;
	wire        [31:0] w_sys_tmp574;
	wire signed [31:0] w_sys_tmp575;
	wire signed [31:0] w_sys_tmp576;
	wire signed [31:0] w_sys_tmp577;
	wire signed [31:0] w_sys_tmp579;
	wire               w_sys_tmp580;
	wire               w_sys_tmp581;
	wire signed [31:0] w_sys_tmp584;
	wire signed [31:0] w_sys_tmp585;
	wire signed [31:0] w_sys_tmp586;
	wire        [31:0] w_sys_tmp587;
	wire signed [31:0] w_sys_tmp589;
	wire signed [31:0] w_sys_tmp590;
	wire signed [31:0] w_sys_tmp593;
	wire signed [31:0] w_sys_tmp594;
	wire signed [31:0] w_sys_tmp811;
	wire signed [31:0] w_sys_tmp812;
	wire               w_sys_tmp813;
	wire               w_sys_tmp814;
	wire signed [31:0] w_sys_tmp815;
	wire signed [31:0] w_sys_tmp816;
	wire signed [31:0] w_sys_tmp819;
	wire signed [31:0] w_sys_tmp820;
	wire signed [31:0] w_sys_tmp821;
	wire        [31:0] w_sys_tmp822;
	wire signed [31:0] w_sys_tmp823;
	wire signed [31:0] w_sys_tmp932;
	wire               w_sys_tmp933;
	wire               w_sys_tmp934;
	wire signed [31:0] w_sys_tmp935;
	wire signed [31:0] w_sys_tmp936;
	wire signed [31:0] w_sys_tmp937;
	wire               w_sys_tmp938;
	wire               w_sys_tmp939;
	wire signed [31:0] w_sys_tmp940;
	wire signed [31:0] w_sys_tmp943;
	wire signed [31:0] w_sys_tmp944;
	wire signed [31:0] w_sys_tmp945;
	wire        [31:0] w_sys_tmp946;
	wire signed [31:0] w_sys_tmp947;
	wire signed [31:0] w_sys_tmp948;
	wire        [31:0] w_sys_tmp950;
	wire signed [31:0] w_sys_tmp951;
	wire signed [31:0] w_sys_tmp952;
	wire signed [31:0] w_sys_tmp954;
	wire signed [31:0] w_sys_tmp955;
	wire signed [31:0] w_sys_tmp956;
	wire        [31:0] w_sys_tmp958;
	wire signed [31:0] w_sys_tmp959;
	wire signed [31:0] w_sys_tmp960;
	wire signed [31:0] w_sys_tmp961;
	wire signed [31:0] w_sys_tmp963;
	wire signed [31:0] w_sys_tmp964;
	wire signed [31:0] w_sys_tmp966;
	wire signed [31:0] w_sys_tmp967;
	wire signed [31:0] w_sys_tmp968;
	wire signed [31:0] w_sys_tmp971;
	wire signed [31:0] w_sys_tmp972;
	wire signed [31:0] w_sys_tmp973;
	wire signed [31:0] w_sys_tmp975;
	wire signed [31:0] w_sys_tmp976;
	wire signed [31:0] w_sys_tmp977;
	wire        [31:0] w_sys_tmp979;
	wire        [31:0] w_sys_tmp980;
	wire signed [31:0] w_sys_tmp982;
	wire signed [31:0] w_sys_tmp983;
	wire signed [31:0] w_sys_tmp985;
	wire signed [31:0] w_sys_tmp986;
	wire signed [31:0] w_sys_tmp987;
	wire signed [31:0] w_sys_tmp991;
	wire signed [31:0] w_sys_tmp992;
	wire signed [31:0] w_sys_tmp993;
	wire signed [31:0] w_sys_tmp997;
	wire signed [31:0] w_sys_tmp998;
	wire signed [31:0] w_sys_tmp1000;
	wire signed [31:0] w_sys_tmp1001;
	wire signed [31:0] w_sys_tmp1002;
	wire signed [31:0] w_sys_tmp1004;
	wire signed [31:0] w_sys_tmp1005;
	wire signed [31:0] w_sys_tmp1006;
	wire signed [31:0] w_sys_tmp1007;
	wire signed [31:0] w_sys_tmp1008;
	wire signed [31:0] w_sys_tmp1010;
	wire signed [31:0] w_sys_tmp1011;
	wire signed [31:0] w_sys_tmp1012;
	wire signed [31:0] w_sys_tmp1013;
	wire signed [31:0] w_sys_tmp1015;
	wire signed [31:0] w_sys_tmp1016;
	wire signed [31:0] w_sys_tmp1017;
	wire signed [31:0] w_sys_tmp2463;
	wire               w_sys_tmp2464;
	wire               w_sys_tmp2465;
	wire signed [31:0] w_sys_tmp2466;
	wire signed [31:0] w_sys_tmp2467;
	wire signed [31:0] w_sys_tmp2468;
	wire               w_sys_tmp2469;
	wire               w_sys_tmp2470;
	wire signed [31:0] w_sys_tmp2471;
	wire signed [31:0] w_sys_tmp2474;
	wire signed [31:0] w_sys_tmp2475;
	wire signed [31:0] w_sys_tmp2476;
	wire        [31:0] w_sys_tmp2477;
	wire signed [31:0] w_sys_tmp2478;
	wire signed [31:0] w_sys_tmp2479;
	wire signed [31:0] w_sys_tmp2481;
	wire signed [31:0] w_sys_tmp2482;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 2'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 8'h1);
	assign w_fld_T_0_addr_0 = 10'sh0;
	assign w_fld_T_0_datain_0 = 32'h0;
	assign w_fld_T_0_r_w_0 = 1'h0;
	assign w_fld_T_0_ce_0 = w_sys_ce;
	assign w_fld_T_0_ce_1 = w_sys_ce;
	assign w_fld_TT_1_addr_0 = 10'sh0;
	assign w_fld_TT_1_datain_0 = 32'h0;
	assign w_fld_TT_1_r_w_0 = 1'h0;
	assign w_fld_TT_1_ce_0 = w_sys_ce;
	assign w_fld_TT_1_ce_1 = w_sys_ce;
	assign w_fld_U_2_addr_0 = 10'sh0;
	assign w_fld_U_2_datain_0 = 32'h0;
	assign w_fld_U_2_r_w_0 = 1'h0;
	assign w_fld_U_2_ce_0 = w_sys_ce;
	assign w_fld_U_2_ce_1 = w_sys_ce;
	assign w_fld_V_3_addr_0 = 10'sh0;
	assign w_fld_V_3_datain_0 = 32'h0;
	assign w_fld_V_3_r_w_0 = 1'h0;
	assign w_fld_V_3_ce_0 = w_sys_ce;
	assign w_fld_V_3_ce_1 = w_sys_ce;
	assign w_sys_tmp1 = 32'sh0000000a;
	assign w_sys_tmp3 = 32'sh0000000b;
	assign w_sys_tmp5 = 32'h3a03126f;
	assign w_sys_tmp6 = 32'h3ecccccd;
	assign w_sys_tmp7 = 32'h3dcccccd;
	assign w_sys_tmp8 = 32'h3a23d70b;
	assign w_sys_tmp9 = 32'h3b23d70b;
	assign w_sys_tmp10 = 32'h3b4ccccc;
	assign w_sys_tmp11 = 32'h3d4ccccc;
	assign w_sys_tmp12 = ( !w_sys_tmp13 );
	assign w_sys_tmp13 = (r_run_my_8 < r_run_k_4);
	assign w_sys_tmp14 = (r_run_k_4 + w_sys_intOne);
	assign w_sys_tmp15 = ( !w_sys_tmp16 );
	assign w_sys_tmp16 = (r_run_mx_7 < r_run_j_5);
	assign w_sys_tmp18 = w_ip_MultFloat_product_0;
	assign w_sys_tmp19 = w_ip_FixedToFloat_floating_0;
	assign w_sys_tmp20 = (r_run_k_4 - w_sys_intOne);
	assign w_sys_tmp22 = (w_sys_tmp23 + r_run_k_4);
	assign w_sys_tmp23 = (r_run_j_5 * w_sys_tmp24);
	assign w_sys_tmp24 = 32'sh0000000b;
	assign w_sys_tmp25 = 32'h0;
	assign w_sys_tmp27 = (w_sys_tmp28 + r_run_k_4);
	assign w_sys_tmp28 = (r_run_copy2_j_22 * w_sys_tmp24);
	assign w_sys_tmp32 = (w_sys_tmp33 + r_run_k_4);
	assign w_sys_tmp33 = (r_run_copy1_j_21 * w_sys_tmp24);
	assign w_sys_tmp36 = 32'h42200000;
	assign w_sys_tmp37 = w_sys_tmp18;
	assign w_sys_tmp38 = 32'h3f800000;
	assign w_sys_tmp41 = (w_sys_tmp42 + r_run_k_4);
	assign w_sys_tmp42 = (r_run_copy0_j_20 * w_sys_tmp24);
	assign w_sys_tmp45 = (r_run_copy0_j_20 + w_sys_intOne);
	assign w_sys_tmp46 = (r_run_copy1_j_21 + w_sys_intOne);
	assign w_sys_tmp47 = (r_run_copy2_j_22 + w_sys_intOne);
	assign w_sys_tmp48 = (r_run_j_5 + w_sys_intOne);
	assign w_sys_tmp128 = r_sys_tmp16_float;
	assign w_sys_tmp157 = r_sys_tmp15_float;
	assign w_sys_tmp185 = r_sys_tmp13_float;
	assign w_sys_tmp213 = r_sys_tmp10_float;
	assign w_sys_tmp269 = r_sys_tmp8_float;
	assign w_sys_tmp297 = r_sys_tmp5_float;
	assign w_sys_tmp560 = ( !w_sys_tmp561 );
	assign w_sys_tmp561 = (r_run_nlast_19 < r_run_n_6);
	assign w_sys_tmp562 = (r_run_n_6 + w_sys_intOne);
	assign w_sys_tmp563 = ( !w_sys_tmp564 );
	assign w_sys_tmp564 = (r_run_my_8 < r_run_k_4);
	assign w_sys_tmp567 = (w_sys_tmp568 + r_run_k_4);
	assign w_sys_tmp568 = 32'sh0000000b;
	assign w_sys_tmp569 = 32'h0;
	assign w_sys_tmp571 = (w_sys_tmp572 + r_run_k_4);
	assign w_sys_tmp572 = (r_run_mx_7 * w_sys_tmp568);
	assign w_sys_tmp574 = w_fld_T_0_dataout_1;
	assign w_sys_tmp575 = (w_sys_tmp576 + r_run_k_4);
	assign w_sys_tmp576 = (w_sys_tmp577 * w_sys_tmp568);
	assign w_sys_tmp577 = (r_run_mx_7 - w_sys_intOne);
	assign w_sys_tmp579 = (r_run_k_4 + w_sys_intOne);
	assign w_sys_tmp580 = ( !w_sys_tmp581 );
	assign w_sys_tmp581 = (r_run_mx_7 < r_run_j_5);
	assign w_sys_tmp584 = (w_sys_tmp585 + w_sys_intOne);
	assign w_sys_tmp585 = (r_run_j_5 * w_sys_tmp586);
	assign w_sys_tmp586 = 32'sh0000000b;
	assign w_sys_tmp587 = 32'h0;
	assign w_sys_tmp589 = (w_sys_tmp590 + r_run_my_8);
	assign w_sys_tmp590 = (r_run_copy0_j_23 * w_sys_tmp586);
	assign w_sys_tmp593 = (r_run_copy0_j_23 + w_sys_intOne);
	assign w_sys_tmp594 = (r_run_j_5 + w_sys_intOne);
	assign w_sys_tmp811 = w_ip_DivInt_quotient_0;
	assign w_sys_tmp812 = 32'sh00000004;
	assign w_sys_tmp813 = ( !w_sys_tmp814 );
	assign w_sys_tmp814 = (w_sys_tmp815 < r_run_j_5);
	assign w_sys_tmp815 = w_ip_DivInt_quotient_1;
	assign w_sys_tmp816 = 32'sh00000002;
	assign w_sys_tmp819 = (w_sys_tmp820 + w_sys_intOne);
	assign w_sys_tmp820 = (r_run_j_5 * w_sys_tmp821);
	assign w_sys_tmp821 = 32'sh0000000b;
	assign w_sys_tmp822 = 32'h3f800000;
	assign w_sys_tmp823 = (r_run_j_5 + w_sys_intOne);
	assign w_sys_tmp932 = 32'sh00000002;
	assign w_sys_tmp933 = ( !w_sys_tmp934 );
	assign w_sys_tmp934 = (w_sys_tmp935 < r_run_k_4);
	assign w_sys_tmp935 = (r_run_my_8 - w_sys_intOne);
	assign w_sys_tmp936 = (r_run_k_4 + w_sys_intOne);
	assign w_sys_tmp937 = 32'sh00000002;
	assign w_sys_tmp938 = ( !w_sys_tmp939 );
	assign w_sys_tmp939 = (w_sys_tmp940 < r_run_j_5);
	assign w_sys_tmp940 = (r_run_mx_7 - w_sys_intOne);
	assign w_sys_tmp943 = (w_sys_tmp944 + r_run_k_4);
	assign w_sys_tmp944 = (r_run_j_5 * w_sys_tmp945);
	assign w_sys_tmp945 = 32'sh0000000b;
	assign w_sys_tmp946 = w_ip_AddFloat_result_0;
	assign w_sys_tmp947 = (w_sys_tmp948 + r_run_k_4);
	assign w_sys_tmp948 = (r_run_copy12_j_36 * w_sys_tmp945);
	assign w_sys_tmp950 = w_fld_U_2_dataout_1;
	assign w_sys_tmp951 = (w_sys_tmp952 + r_run_k_4);
	assign w_sys_tmp952 = (r_run_copy11_j_35 * w_sys_tmp945);
	assign w_sys_tmp954 = (w_sys_tmp955 + r_run_k_4);
	assign w_sys_tmp955 = (w_sys_tmp956 * w_sys_tmp945);
	assign w_sys_tmp956 = (r_run_copy10_j_34 + w_sys_intOne);
	assign w_sys_tmp958 = w_fld_T_0_dataout_1;
	assign w_sys_tmp959 = (w_sys_tmp960 + r_run_k_4);
	assign w_sys_tmp960 = (w_sys_tmp961 * w_sys_tmp945);
	assign w_sys_tmp961 = (r_run_copy9_j_33 - w_sys_intOne);
	assign w_sys_tmp963 = (w_sys_tmp964 + r_run_k_4);
	assign w_sys_tmp964 = (r_run_copy8_j_32 * w_sys_tmp945);
	assign w_sys_tmp966 = (w_sys_tmp967 + w_sys_intOne);
	assign w_sys_tmp967 = (w_sys_tmp968 + r_run_k_4);
	assign w_sys_tmp968 = (r_run_copy7_j_31 * w_sys_tmp945);
	assign w_sys_tmp971 = (w_sys_tmp972 - w_sys_intOne);
	assign w_sys_tmp972 = (w_sys_tmp973 + r_run_k_4);
	assign w_sys_tmp973 = (r_run_copy6_j_30 * w_sys_tmp945);
	assign w_sys_tmp975 = (w_sys_tmp976 + r_run_k_4);
	assign w_sys_tmp976 = (w_sys_tmp977 * w_sys_tmp945);
	assign w_sys_tmp977 = (r_run_copy5_j_29 + w_sys_intOne);
	assign w_sys_tmp979 = w_ip_MultFloat_product_0;
	assign w_sys_tmp980 = 32'h40000000;
	assign w_sys_tmp982 = (w_sys_tmp983 + r_run_k_4);
	assign w_sys_tmp983 = (r_run_copy4_j_28 * w_sys_tmp945);
	assign w_sys_tmp985 = (w_sys_tmp986 + r_run_k_4);
	assign w_sys_tmp986 = (w_sys_tmp987 * w_sys_tmp945);
	assign w_sys_tmp987 = (r_run_copy3_j_27 - w_sys_intOne);
	assign w_sys_tmp991 = (w_sys_tmp992 + w_sys_intOne);
	assign w_sys_tmp992 = (w_sys_tmp993 + r_run_k_4);
	assign w_sys_tmp993 = (r_run_copy2_j_26 * w_sys_tmp945);
	assign w_sys_tmp997 = (w_sys_tmp998 + r_run_k_4);
	assign w_sys_tmp998 = (r_run_copy1_j_25 * w_sys_tmp945);
	assign w_sys_tmp1000 = (w_sys_tmp1001 - w_sys_intOne);
	assign w_sys_tmp1001 = (w_sys_tmp1002 + r_run_k_4);
	assign w_sys_tmp1002 = (r_run_copy0_j_24 * w_sys_tmp945);
	assign w_sys_tmp1004 = (r_run_copy0_j_24 + w_sys_intOne);
	assign w_sys_tmp1005 = (r_run_copy1_j_25 + w_sys_intOne);
	assign w_sys_tmp1006 = (r_run_copy2_j_26 + w_sys_intOne);
	assign w_sys_tmp1007 = (r_run_copy3_j_27 + w_sys_intOne);
	assign w_sys_tmp1008 = (r_run_copy4_j_28 + w_sys_intOne);
	assign w_sys_tmp1010 = (r_run_copy6_j_30 + w_sys_intOne);
	assign w_sys_tmp1011 = (r_run_copy7_j_31 + w_sys_intOne);
	assign w_sys_tmp1012 = (r_run_copy8_j_32 + w_sys_intOne);
	assign w_sys_tmp1013 = (r_run_copy9_j_33 + w_sys_intOne);
	assign w_sys_tmp1015 = (r_run_copy11_j_35 + w_sys_intOne);
	assign w_sys_tmp1016 = (r_run_copy12_j_36 + w_sys_intOne);
	assign w_sys_tmp1017 = (r_run_j_5 + w_sys_intOne);
	assign w_sys_tmp2463 = 32'sh00000002;
	assign w_sys_tmp2464 = ( !w_sys_tmp2465 );
	assign w_sys_tmp2465 = (w_sys_tmp2466 < r_run_k_4);
	assign w_sys_tmp2466 = (r_run_my_8 - w_sys_intOne);
	assign w_sys_tmp2467 = (r_run_k_4 + w_sys_intOne);
	assign w_sys_tmp2468 = 32'sh00000002;
	assign w_sys_tmp2469 = ( !w_sys_tmp2470 );
	assign w_sys_tmp2470 = (w_sys_tmp2471 < r_run_j_5);
	assign w_sys_tmp2471 = (r_run_mx_7 - w_sys_intOne);
	assign w_sys_tmp2474 = (w_sys_tmp2475 + r_run_k_4);
	assign w_sys_tmp2475 = (r_run_j_5 * w_sys_tmp2476);
	assign w_sys_tmp2476 = 32'sh0000000b;
	assign w_sys_tmp2477 = w_fld_TT_1_dataout_1;
	assign w_sys_tmp2478 = (w_sys_tmp2479 + r_run_k_4);
	assign w_sys_tmp2479 = (r_run_copy0_j_37 * w_sys_tmp2476);
	assign w_sys_tmp2481 = (r_run_copy0_j_37 + w_sys_intOne);
	assign w_sys_tmp2482 = (r_run_j_5 + w_sys_intOne);


	DualPortRAM #(.DWIDTH(32), .AWIDTH(10), .WORDS(1024) )
		dpram_T_0(
			.clk (clock),
			.ce_0 (w_fld_T_0_ce_0),
			.addr_0 (w_fld_T_0_addr_0),
			.datain_0 (w_fld_T_0_datain_0),
			.dataout_0 (w_fld_T_0_dataout_0),
			.r_w_0 (w_fld_T_0_r_w_0),
			.ce_1 (w_fld_T_0_ce_1),
			.addr_1 (r_fld_T_0_addr_1),
			.datain_1 (r_fld_T_0_datain_1),
			.dataout_1 (w_fld_T_0_dataout_1),
			.r_w_1 (r_fld_T_0_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(10), .WORDS(1024) )
		dpram_TT_1(
			.clk (clock),
			.ce_0 (w_fld_TT_1_ce_0),
			.addr_0 (w_fld_TT_1_addr_0),
			.datain_0 (w_fld_TT_1_datain_0),
			.dataout_0 (w_fld_TT_1_dataout_0),
			.r_w_0 (w_fld_TT_1_r_w_0),
			.ce_1 (w_fld_TT_1_ce_1),
			.addr_1 (r_fld_TT_1_addr_1),
			.datain_1 (r_fld_TT_1_datain_1),
			.dataout_1 (w_fld_TT_1_dataout_1),
			.r_w_1 (r_fld_TT_1_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(10), .WORDS(1024) )
		dpram_U_2(
			.clk (clock),
			.ce_0 (w_fld_U_2_ce_0),
			.addr_0 (w_fld_U_2_addr_0),
			.datain_0 (w_fld_U_2_datain_0),
			.dataout_0 (w_fld_U_2_dataout_0),
			.r_w_0 (w_fld_U_2_r_w_0),
			.ce_1 (w_fld_U_2_ce_1),
			.addr_1 (r_fld_U_2_addr_1),
			.datain_1 (r_fld_U_2_datain_1),
			.dataout_1 (w_fld_U_2_dataout_1),
			.r_w_1 (r_fld_U_2_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(10), .WORDS(1024) )
		dpram_V_3(
			.clk (clock),
			.ce_0 (w_fld_V_3_ce_0),
			.addr_0 (w_fld_V_3_addr_0),
			.datain_0 (w_fld_V_3_datain_0),
			.dataout_0 (w_fld_V_3_dataout_0),
			.r_w_0 (w_fld_V_3_r_w_0),
			.ce_1 (w_fld_V_3_ce_1),
			.addr_1 (r_fld_V_3_addr_1),
			.datain_1 (r_fld_V_3_datain_1),
			.dataout_1 (w_fld_V_3_dataout_1),
			.r_w_1 (r_fld_V_3_r_w_1)
		);

	DivInt
		DivInt_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.dividend (r_ip_DivInt_dividend_0),
			.divisor (r_ip_DivInt_divisor_0),
			.fractional (w_ip_DivInt_fractional_0),
			.quotient (w_ip_DivInt_quotient_0)
		);

	DivInt
		DivInt_inst_1(
			.clk (clock),
			.ce (w_sys_ce),
			.dividend (r_ip_DivInt_dividend_1),
			.divisor (r_ip_DivInt_divisor_1),
			.fractional (w_ip_DivInt_fractional_1),
			.quotient (w_ip_DivInt_quotient_1)
		);

	AddFloat
		AddFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_AddFloat_portA_0),
			.b (r_ip_AddFloat_portB_0),
			.result (w_ip_AddFloat_result_0)
		);

	MultFloat
		MultFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_MultFloat_multiplicand_0),
			.b (r_ip_MultFloat_multiplier_0),
			.result (w_ip_MultFloat_product_0)
		);

	FixedToFloat
		FixedToFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_FixedToFloat_fixed_0),
			.result (w_ip_FixedToFloat_floating_0)
		);

	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h20: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_ip_DivInt_dividend_0 <= r_run_mx_7;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h20: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_ip_DivInt_divisor_0 <= w_sys_tmp812;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h21: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_ip_DivInt_dividend_1 <= r_run_mx_7;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h21: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_ip_DivInt_divisor_1 <= w_sys_tmp816;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hc) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h32) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h38)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp38;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h17) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h3e) || (r_sys_run_step==8'h3f) || (r_sys_run_step==8'h41) || (r_sys_run_step==8'h49) || (r_sys_run_step==8'h4a) || (r_sys_run_step==8'h4c) || (r_sys_run_step==8'h54) || (r_sys_run_step==8'h55) || (r_sys_run_step==8'h57) || (r_sys_run_step==8'h5f) || (r_sys_run_step==8'h60) || (r_sys_run_step==8'h62) || (r_sys_run_step==8'h6a) || (r_sys_run_step==8'h6b) || (r_sys_run_step==8'h6d) || (r_sys_run_step==8'h75) || (r_sys_run_step==8'h76) || (r_sys_run_step==8'h78) || (r_sys_run_step==8'h80) || (r_sys_run_step==8'h81) || (r_sys_run_step==8'h83) || (r_sys_run_step==8'h8b) || (r_sys_run_step==8'h8c) || (r_sys_run_step==8'h8e) || (r_sys_run_step==8'h96) || (r_sys_run_step==8'h97) || (r_sys_run_step==8'h99) || (r_sys_run_step==8'ha1) || (r_sys_run_step==8'ha2) || (r_sys_run_step==8'ha4) || (r_sys_run_step==8'hac) || (r_sys_run_step==8'had) || (r_sys_run_step==8'haf) || (r_sys_run_step==8'hb7) || (r_sys_run_step==8'hb8) || (r_sys_run_step==8'hba) || (r_sys_run_step==8'hc2) || (r_sys_run_step==8'hc3) || (r_sys_run_step==8'hc5) || (r_sys_run_step==8'hcd) || (r_sys_run_step==8'hce) || (r_sys_run_step==8'hd0) || (r_sys_run_step==8'hd8) || (r_sys_run_step==8'hd9) || (r_sys_run_step==8'hdb) || (r_sys_run_step==8'hdf) || (r_sys_run_step==8'he7)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp946;

									end
									else
									if((r_sys_run_step==8'h4e)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp26_float;

									end
									else
									if((r_sys_run_step==8'h37)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp33_float;

									end
									else
									if((r_sys_run_step==8'h35) || (r_sys_run_step==8'h40) || (r_sys_run_step==8'h58)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp31_float;

									end
									else
									if((r_sys_run_step==8'h42) || (r_sys_run_step==8'h4b) || (r_sys_run_step==8'h56) || (r_sys_run_step==8'h61) || (r_sys_run_step==8'h6c) || (r_sys_run_step==8'h77) || (r_sys_run_step==8'h82) || (r_sys_run_step==8'h8d) || (r_sys_run_step==8'h98) || (r_sys_run_step==8'ha3) || (r_sys_run_step==8'hae) || (r_sys_run_step==8'hb9) || (r_sys_run_step==8'hc4) || (r_sys_run_step==8'hcf) || (r_sys_run_step==8'hda) || (r_sys_run_step==8'he2)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp44_float;

									end
									else
									if((r_sys_run_step==8'h10) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h3b) || (r_sys_run_step==8'h3d) || (r_sys_run_step==8'h44) || (r_sys_run_step==8'h50) || (r_sys_run_step==8'h51) || (r_sys_run_step==8'h53) || (r_sys_run_step==8'h5a) || (r_sys_run_step==8'h66) || (r_sys_run_step==8'h67) || (r_sys_run_step==8'h69) || (r_sys_run_step==8'h70) || (r_sys_run_step==8'h7c) || (r_sys_run_step==8'h7d) || (r_sys_run_step==8'h7f) || (r_sys_run_step==8'h86) || (r_sys_run_step==8'h92) || (r_sys_run_step==8'h93) || (r_sys_run_step==8'h95) || (r_sys_run_step==8'h9c) || (r_sys_run_step==8'ha8) || (r_sys_run_step==8'ha9) || (r_sys_run_step==8'hab) || (r_sys_run_step==8'hb2) || (r_sys_run_step==8'hbe) || (r_sys_run_step==8'hbf) || (r_sys_run_step==8'hc1) || (r_sys_run_step==8'hc8) || (r_sys_run_step==8'hd4)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp42_float;

									end
									else
									if((r_sys_run_step==8'h38) || (r_sys_run_step==8'h4d)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp22_float;

									end
									else
									if((r_sys_run_step==8'hf) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h59) || (r_sys_run_step==8'h63) || (r_sys_run_step==8'h6e) || (r_sys_run_step==8'h79) || (r_sys_run_step==8'h84) || (r_sys_run_step==8'h8f) || (r_sys_run_step==8'h9a) || (r_sys_run_step==8'ha5) || (r_sys_run_step==8'hb0) || (r_sys_run_step==8'hbb) || (r_sys_run_step==8'hc6) || (r_sys_run_step==8'hd1) || (r_sys_run_step==8'hd5)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp41_float;

									end
									else
									if((r_sys_run_step==8'h12) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h3c) || (r_sys_run_step==8'h47) || (r_sys_run_step==8'h52) || (r_sys_run_step==8'h5d) || (r_sys_run_step==8'h68) || (r_sys_run_step==8'h73) || (r_sys_run_step==8'h7e) || (r_sys_run_step==8'h89) || (r_sys_run_step==8'h94) || (r_sys_run_step==8'h9f) || (r_sys_run_step==8'haa) || (r_sys_run_step==8'hb5) || (r_sys_run_step==8'hc0) || (r_sys_run_step==8'hcb) || (r_sys_run_step==8'hd6)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp40_float;

									end
									else
									if((r_sys_run_step==8'h4) || (r_sys_run_step==8'h6) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h2f) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h32) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h45) || (r_sys_run_step==8'h46) || (r_sys_run_step==8'h48) || (r_sys_run_step==8'h4f) || (r_sys_run_step==8'h5b) || (r_sys_run_step==8'h5c) || (r_sys_run_step==8'h5e) || (r_sys_run_step==8'h65) || (r_sys_run_step==8'h71) || (r_sys_run_step==8'h72) || (r_sys_run_step==8'h74) || (r_sys_run_step==8'h7b) || (r_sys_run_step==8'h87) || (r_sys_run_step==8'h88) || (r_sys_run_step==8'h8a) || (r_sys_run_step==8'h91) || (r_sys_run_step==8'h9d) || (r_sys_run_step==8'h9e) || (r_sys_run_step==8'ha0) || (r_sys_run_step==8'ha7) || (r_sys_run_step==8'hb3) || (r_sys_run_step==8'hb4) || (r_sys_run_step==8'hb6) || (r_sys_run_step==8'hbd) || (r_sys_run_step==8'hc9) || (r_sys_run_step==8'hca) || (r_sys_run_step==8'hcc) || (r_sys_run_step==8'hd3)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp43_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hc)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp269[31], w_sys_tmp269[30:0] };

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
									else
									if((r_sys_run_step==8'h32)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp297[31], w_sys_tmp297[30:0] };

									end
									else
									if((r_sys_run_step==8'h36)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp269[31], w_sys_tmp269[30:0] };

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp185[31], w_sys_tmp185[30:0] };

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp269[31], w_sys_tmp269[30:0] };

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp128[31], w_sys_tmp128[30:0] };

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp185[31], w_sys_tmp185[30:0] };

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp213[31], w_sys_tmp213[30:0] };

									end
									else
									if((r_sys_run_step==8'h34)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp185[31], w_sys_tmp185[30:0] };

									end
									else
									if((r_sys_run_step==8'h30)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp269[31], w_sys_tmp269[30:0] };

									end
									else
									if((r_sys_run_step==8'h21)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp297[31], w_sys_tmp297[30:0] };

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp185[31], w_sys_tmp185[30:0] };

									end
									else
									if((r_sys_run_step==8'h38)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp157[31], w_sys_tmp157[30:0] };

									end
									else
									if((r_sys_run_step==8'h2d)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp185[31], w_sys_tmp185[30:0] };

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp157[31], w_sys_tmp157[30:0] };

									end
									else
									if((r_sys_run_step==8'h2a)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp297[31], w_sys_tmp297[30:0] };

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h18)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'hd3)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'h76)) begin
										r_ip_AddFloat_portB_0 <= { ~r_sys_tmp37_float[31], r_sys_tmp37_float[30:0] };

									end
									else
									if((r_sys_run_step==8'hca)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'h4a)) begin
										r_ip_AddFloat_portB_0 <= { ~r_sys_tmp27_float[31], r_sys_tmp27_float[30:0] };

									end
									else
									if((r_sys_run_step==8'h2f)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'haa)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h39)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h31)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h86)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'hd6)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'h7e)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h30)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'ha8)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h5e)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_ip_AddFloat_portB_0 <= { ~r_sys_tmp34_float[31], r_sys_tmp34_float[30:0] };

									end
									else
									if((r_sys_run_step==8'h52)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h56)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp40_float;

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h89)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'hc9)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'hb6)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'h95)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'h9e)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'h84) || (r_sys_run_step==8'h9a) || (r_sys_run_step==8'hb0) || (r_sys_run_step==8'hc6) || (r_sys_run_step==8'hd5) || (r_sys_run_step==8'hdf) || (r_sys_run_step==8'he7)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp37_float;

									end
									else
									if((r_sys_run_step==8'h91)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h63) || (r_sys_run_step==8'h79) || (r_sys_run_step==8'h8f) || (r_sys_run_step==8'ha5) || (r_sys_run_step==8'hbb) || (r_sys_run_step==8'hd1) || (r_sys_run_step==8'hda)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp36_float;

									end
									else
									if((r_sys_run_step==8'hb3)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h93)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'hb4)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'h53)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'h7f)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'hc8)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'had)) begin
										r_ip_AddFloat_portB_0 <= { ~r_sys_tmp36_float[31], r_sys_tmp36_float[30:0] };

									end
									else
									if((r_sys_run_step==8'h40)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp32_float;

									end
									else
									if((r_sys_run_step==8'hbf)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'hd4)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h38) || (r_sys_run_step==8'h42) || (r_sys_run_step==8'he2)) begin
										r_ip_AddFloat_portB_0 <= w_sys_tmp979;

									end
									else
									if((r_sys_run_step==8'h13) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h3e) || (r_sys_run_step==8'h49) || (r_sys_run_step==8'h54) || (r_sys_run_step==8'h5f) || (r_sys_run_step==8'h6a) || (r_sys_run_step==8'h75) || (r_sys_run_step==8'h80) || (r_sys_run_step==8'h8b) || (r_sys_run_step==8'h96) || (r_sys_run_step==8'ha1) || (r_sys_run_step==8'hac) || (r_sys_run_step==8'hb7) || (r_sys_run_step==8'hc2) || (r_sys_run_step==8'hcd) || (r_sys_run_step==8'hd8)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp39_float;

									end
									else
									if((r_sys_run_step==8'h51)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'h87)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_ip_AddFloat_portB_0 <= { ~r_sys_tmp24_float[31], r_sys_tmp24_float[30:0] };

									end
									else
									if((r_sys_run_step==8'hb8)) begin
										r_ip_AddFloat_portB_0 <= { ~r_sys_tmp37_float[31], r_sys_tmp37_float[30:0] };

									end
									else
									if((r_sys_run_step==8'h2e)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h66)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h37)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp21_float;

									end
									else
									if((r_sys_run_step==8'h7c)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h6b)) begin
										r_ip_AddFloat_portB_0 <= { ~r_sys_tmp36_float[31], r_sys_tmp36_float[30:0] };

									end
									else
									if((r_sys_run_step==8'h3d)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'h55)) begin
										r_ip_AddFloat_portB_0 <= { ~r_sys_tmp34_float[31], r_sys_tmp34_float[30:0] };

									end
									else
									if((r_sys_run_step==8'h17) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h41) || (r_sys_run_step==8'h4c) || (r_sys_run_step==8'h57) || (r_sys_run_step==8'h62) || (r_sys_run_step==8'h6d) || (r_sys_run_step==8'h78) || (r_sys_run_step==8'h83) || (r_sys_run_step==8'h8e) || (r_sys_run_step==8'h99) || (r_sys_run_step==8'ha4) || (r_sys_run_step==8'haf) || (r_sys_run_step==8'hba) || (r_sys_run_step==8'hc5) || (r_sys_run_step==8'hd0) || (r_sys_run_step==8'hdb)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp38_float;

									end
									else
									if((r_sys_run_step==8'ha0)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'h74)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'hbd)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h9c)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'h72)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'h65)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h34)) begin
										r_ip_AddFloat_portB_0 <= { ~r_sys_tmp29_float[31], r_sys_tmp29_float[30:0] };

									end
									else
									if((r_sys_run_step==8'h50)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'hab)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'ha9)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'hcb)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'hcc)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'h70)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'hc0)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h47)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'hce)) begin
										r_ip_AddFloat_portB_0 <= { ~r_sys_tmp37_float[31], r_sys_tmp37_float[30:0] };

									end
									else
									if((r_sys_run_step==8'h5d)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h5c)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'h88)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'h3a)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h3b)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h8a)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'h4f)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h3f)) begin
										r_ip_AddFloat_portB_0 <= { ~r_sys_tmp32_float[31], r_sys_tmp32_float[30:0] };

									end
									else
									if((r_sys_run_step==8'hb5)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h29)) begin
										r_ip_AddFloat_portB_0 <= { ~r_sys_tmp23_float[31], r_sys_tmp23_float[30:0] };

									end
									else
									if((r_sys_run_step==8'h5b)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h94)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h4d) || (r_sys_run_step==8'h58)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp28_float;

									end
									else
									if((r_sys_run_step==8'h46)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'h92)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'hb2)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h21)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_ip_AddFloat_portB_0 <= { ~r_sys_tmp34_float[31], r_sys_tmp34_float[30:0] };

									end
									else
									if((r_sys_run_step==8'h73)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h71)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h59) || (r_sys_run_step==8'h6e) || (r_sys_run_step==8'h77) || (r_sys_run_step==8'h82) || (r_sys_run_step==8'h8d) || (r_sys_run_step==8'h98) || (r_sys_run_step==8'ha3) || (r_sys_run_step==8'hae) || (r_sys_run_step==8'hb9) || (r_sys_run_step==8'hc4) || (r_sys_run_step==8'hcf)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp35_float;

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h7d)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'h67)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'h4b)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp33_float;

									end
									else
									if((r_sys_run_step==8'h48)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'hc3)) begin
										r_ip_AddFloat_portB_0 <= { ~r_sys_tmp36_float[31], r_sys_tmp36_float[30:0] };

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h5a)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'ha2)) begin
										r_ip_AddFloat_portB_0 <= { ~r_sys_tmp37_float[31], r_sys_tmp37_float[30:0] };

									end
									else
									if((r_sys_run_step==8'h81)) begin
										r_ip_AddFloat_portB_0 <= { ~r_sys_tmp36_float[31], r_sys_tmp36_float[30:0] };

									end
									else
									if((r_sys_run_step==8'ha7)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h7b)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h44)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'hbe)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h9f)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'hc1)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'h35)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp30_float;

									end
									else
									if((r_sys_run_step==8'h9d)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'h3c)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h60)) begin
										r_ip_AddFloat_portB_0 <= { ~r_sys_tmp35_float[31], r_sys_tmp35_float[30:0] };

									end
									else
									if((r_sys_run_step==8'h69)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'h97)) begin
										r_ip_AddFloat_portB_0 <= { ~r_sys_tmp36_float[31], r_sys_tmp36_float[30:0] };

									end
									else
									if((r_sys_run_step==8'h8c)) begin
										r_ip_AddFloat_portB_0 <= { ~r_sys_tmp37_float[31], r_sys_tmp37_float[30:0] };

									end
									else
									if((r_sys_run_step==8'h32)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp958[31], w_sys_tmp958[30:0] };

									end
									else
									if((r_sys_run_step==8'hd9)) begin
										r_ip_AddFloat_portB_0 <= { ~r_sys_tmp37_float[31], r_sys_tmp37_float[30:0] };

									end
									else
									if((r_sys_run_step==8'h45)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp979[31], w_sys_tmp979[30:0] };

									end
									else
									if((r_sys_run_step==8'h4e) || (r_sys_run_step==8'h61) || (r_sys_run_step==8'h6c)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp34_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hc) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h32) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h3a)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp36;

									end
									else
									if((r_sys_run_step==8'h16) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h2f) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h3c) || (r_sys_run_step==8'h3e)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp16_float;

									end
									else
									if((8'h7<=r_sys_run_step && r_sys_run_step<=8'hb) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h2e)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_dy_11;

									end
									else
									if((r_sys_run_step==8'h20) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h37)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==8'h3f)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp18;

									end
									else
									if((r_sys_run_step==8'h3b)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==8'h1a) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h2c) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h3d)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp15_float;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h3d) || (r_sys_run_step==8'h41) || (r_sys_run_step==8'h46) || (r_sys_run_step==8'h48) || (r_sys_run_step==8'h49) || (r_sys_run_step==8'h51) || (r_sys_run_step==8'h5c) || (r_sys_run_step==8'h67) || (r_sys_run_step==8'h72) || (r_sys_run_step==8'h7d) || (r_sys_run_step==8'h88) || (r_sys_run_step==8'h93) || (r_sys_run_step==8'h9e) || (r_sys_run_step==8'ha9) || (r_sys_run_step==8'hb4) || (r_sys_run_step==8'hbf) || (r_sys_run_step==8'hca) || (r_sys_run_step==8'hd5) || (r_sys_run_step==8'he0)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_r4_15;

									end
									else
									if((r_sys_run_step==8'h8) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h2c) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h37) || (r_sys_run_step==8'h3f) || (r_sys_run_step==8'h42) || (r_sys_run_step==8'h4a) || (r_sys_run_step==8'h4d) || (r_sys_run_step==8'h55) || (r_sys_run_step==8'h58) || (r_sys_run_step==8'h60) || (r_sys_run_step==8'h63) || (r_sys_run_step==8'h6b) || (r_sys_run_step==8'h6e) || (r_sys_run_step==8'h76) || (r_sys_run_step==8'h79) || (r_sys_run_step==8'h81) || (r_sys_run_step==8'h84) || (r_sys_run_step==8'h8c) || (r_sys_run_step==8'h8f) || (r_sys_run_step==8'h97) || (r_sys_run_step==8'h9a) || (r_sys_run_step==8'ha2) || (r_sys_run_step==8'ha5) || (r_sys_run_step==8'had) || (r_sys_run_step==8'hb0) || (r_sys_run_step==8'hb8) || (r_sys_run_step==8'hbb) || (r_sys_run_step==8'hc3) || (r_sys_run_step==8'hc6) || (r_sys_run_step==8'hce) || (r_sys_run_step==8'hd1)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp980;

									end
									else
									if((r_sys_run_step==8'hb1)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp32_float;

									end
									else
									if((r_sys_run_step==8'h85)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==8'hcf)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp25_float;

									end
									else
									if((r_sys_run_step==8'h1f) || (r_sys_run_step==8'h4e)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp35_float;

									end
									else
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h6) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h2f) || (r_sys_run_step==8'h32) || (r_sys_run_step==8'h39)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_r1_12;

									end
									else
									if((r_sys_run_step==8'h61)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==8'h77)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp24_float;

									end
									else
									if((r_sys_run_step==8'hd2)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp33_float;

									end
									else
									if((r_sys_run_step==8'h22) || (r_sys_run_step==8'h59)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h3b) || (r_sys_run_step==8'h3c) || (r_sys_run_step==8'h3e) || (r_sys_run_step==8'h45) || (r_sys_run_step==8'h47)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_r2_13;

									end
									else
									if((r_sys_run_step==8'h64)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp18_float;

									end
									else
									if((r_sys_run_step==8'h38) || (r_sys_run_step==8'h9b)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==8'h40) || (r_sys_run_step==8'ha6)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==8'ha3)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==8'hc7)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp27_float;

									end
									else
									if((r_sys_run_step==8'h8d)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==8'h35) || (r_sys_run_step==8'hc4)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp21_float;

									end
									else
									if((r_sys_run_step==8'h90)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp30_float;

									end
									else
									if((r_sys_run_step==8'ha) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h6f)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp37_float;

									end
									else
									if((r_sys_run_step==8'h2d) || (r_sys_run_step==8'hae)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==8'h82)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==8'h14) || (r_sys_run_step==8'h56)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp36_float;

									end
									else
									if((r_sys_run_step==8'h1c) || (r_sys_run_step==8'h43) || (r_sys_run_step==8'hbc)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp20_float;

									end
									else
									if((r_sys_run_step==8'hb9)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp29_float;

									end
									else
									if((r_sys_run_step==8'h2b) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h44) || (r_sys_run_step==8'h4f) || (r_sys_run_step==8'h5a) || (r_sys_run_step==8'h65) || (r_sys_run_step==8'h70) || (r_sys_run_step==8'h7b) || (r_sys_run_step==8'h86) || (r_sys_run_step==8'h91) || (r_sys_run_step==8'h9c) || (r_sys_run_step==8'ha7) || (r_sys_run_step==8'hb2) || (r_sys_run_step==8'hbd) || (r_sys_run_step==8'hc8) || (r_sys_run_step==8'hd3) || (r_sys_run_step==8'hdd)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_r3_14;

									end
									else
									if((r_sys_run_step==8'h18) || (r_sys_run_step==8'h6c)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp14_float;

									end
									else
									if((r_sys_run_step==8'h98)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp23_float;

									end
									else
									if((r_sys_run_step==8'h7a)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==8'h4b)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp34_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h2b)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==8'h23) || (r_sys_run_step==8'h2f) || (r_sys_run_step==8'h37)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==8'h17) || (r_sys_run_step==8'h28)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==8'h10) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h1f)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==8'hd) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h2e)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp1_float;

									end
									else
									if((8'h7<=r_sys_run_step && r_sys_run_step<=8'hb)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp19;

									end
									else
									if((r_sys_run_step==8'h1d) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h3c)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==8'he) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h32) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h3a)) begin
										r_ip_MultFloat_multiplier_0 <= r_run_YY_16;

									end
									else
									if((r_sys_run_step==8'h16) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h2c) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h3b) || (r_sys_run_step==8'h3e)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp14_float;

									end
									else
									if((r_sys_run_step==8'h1a) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h3d) || (r_sys_run_step==8'h3f)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp37;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h14) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h40) || (r_sys_run_step==8'h4b) || (r_sys_run_step==8'h51) || (r_sys_run_step==8'h56) || (r_sys_run_step==8'h5c) || (r_sys_run_step==8'h61) || (r_sys_run_step==8'h67) || (r_sys_run_step==8'h6c) || (r_sys_run_step==8'h72) || (r_sys_run_step==8'h77) || (r_sys_run_step==8'h7d) || (r_sys_run_step==8'h82) || (r_sys_run_step==8'h88) || (r_sys_run_step==8'h8d) || (r_sys_run_step==8'h93) || (r_sys_run_step==8'h98) || (r_sys_run_step==8'h9e) || (r_sys_run_step==8'ha3) || (r_sys_run_step==8'ha9) || (r_sys_run_step==8'hae) || (r_sys_run_step==8'hb4) || (r_sys_run_step==8'hb9) || (r_sys_run_step==8'hbf) || (r_sys_run_step==8'hc4) || (r_sys_run_step==8'hca) || (r_sys_run_step==8'hcf) || (r_sys_run_step==8'hd5) || (r_sys_run_step==8'hdd) || (r_sys_run_step==8'he0)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp946;

									end
									else
									if((r_sys_run_step==8'h2f)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==8'h15) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h3d)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp26_float;

									end
									else
									if((r_sys_run_step==8'h36)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==8'h47)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==8'hd) || (r_sys_run_step==8'h1b)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp31_float;

									end
									else
									if((r_sys_run_step==8'h45)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp22_float;

									end
									else
									if((r_sys_run_step==8'h3c)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==8'h9) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h24)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp32_float;

									end
									else
									if((r_sys_run_step==8'h32)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==8'h10) || (r_sys_run_step==8'h3b)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp25_float;

									end
									else
									if((r_sys_run_step==8'h2e)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp24_float;

									end
									else
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h48)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp33_float;

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp18_float;

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==8'h11) || (r_sys_run_step==8'h28)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp27_float;

									end
									else
									if((r_sys_run_step==8'h1a) || (r_sys_run_step==8'h41)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp19_float;

									end
									else
									if((r_sys_run_step==8'h39)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==8'ha) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h43) || (r_sys_run_step==8'h44) || (r_sys_run_step==8'h4e) || (r_sys_run_step==8'h4f) || (r_sys_run_step==8'h59) || (r_sys_run_step==8'h5a) || (r_sys_run_step==8'h64) || (r_sys_run_step==8'h65) || (r_sys_run_step==8'h6f) || (r_sys_run_step==8'h70) || (r_sys_run_step==8'h7a) || (r_sys_run_step==8'h7b) || (r_sys_run_step==8'h85) || (r_sys_run_step==8'h86) || (r_sys_run_step==8'h90) || (r_sys_run_step==8'h91) || (r_sys_run_step==8'h9b) || (r_sys_run_step==8'h9c) || (r_sys_run_step==8'ha6) || (r_sys_run_step==8'ha7) || (r_sys_run_step==8'hb1) || (r_sys_run_step==8'hb2) || (r_sys_run_step==8'hbc) || (r_sys_run_step==8'hbd) || (r_sys_run_step==8'hc7) || (r_sys_run_step==8'hc8) || (r_sys_run_step==8'hd2) || (r_sys_run_step==8'hd3)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp44_float;

									end
									else
									if((r_sys_run_step==8'hc) || (r_sys_run_step==8'h27)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp30_float;

									end
									else
									if((r_sys_run_step==8'h22) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h46) || (r_sys_run_step==8'h49)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp41_float;

									end
									else
									if((r_sys_run_step==8'he) || (r_sys_run_step==8'h31)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp29_float;

									end
									else
									if((r_sys_run_step==8'h8) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h2c) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h37) || (r_sys_run_step==8'h3f) || (r_sys_run_step==8'h42) || (r_sys_run_step==8'h4a) || (r_sys_run_step==8'h4d) || (r_sys_run_step==8'h55) || (r_sys_run_step==8'h58) || (r_sys_run_step==8'h60) || (r_sys_run_step==8'h63) || (r_sys_run_step==8'h6b) || (r_sys_run_step==8'h6e) || (r_sys_run_step==8'h76) || (r_sys_run_step==8'h79) || (r_sys_run_step==8'h81) || (r_sys_run_step==8'h84) || (r_sys_run_step==8'h8c) || (r_sys_run_step==8'h8f) || (r_sys_run_step==8'h97) || (r_sys_run_step==8'h9a) || (r_sys_run_step==8'ha2) || (r_sys_run_step==8'ha5) || (r_sys_run_step==8'had) || (r_sys_run_step==8'hb0) || (r_sys_run_step==8'hb8) || (r_sys_run_step==8'hbb) || (r_sys_run_step==8'hc3) || (r_sys_run_step==8'hc6) || (r_sys_run_step==8'hce) || (r_sys_run_step==8'hd1)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp958;

									end
									else
									if((r_sys_run_step==8'h12) || (r_sys_run_step==8'h3e)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp28_float;

									end
									else
									if((r_sys_run_step==8'h20)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp23_float;

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp16_float;

									end
									else
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp950;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h12)) begin
										r_ip_FixedToFloat_fixed_0 <= w_sys_tmp20;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h3c: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 6'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_phase <= 6'h2;
						end

						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h4;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp12) ? 6'h9 : 6'hf);

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'ha;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp15) ? 6'hd : 6'h6);

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h44)) begin
										r_sys_run_phase <= 6'ha;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h10;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp560) ? 6'h14 : 6'h3c);

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h10;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h15;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp563) ? 6'h18 : 6'h1a);

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_run_phase <= 6'h15;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h1b;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp580) ? 6'h1e : 6'h20);

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h25)) begin
										r_sys_run_phase <= 6'h1b;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h21;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h25)) begin
										r_sys_run_phase <= ((w_sys_tmp813) ? 6'h24 : 6'h26);

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h12)) begin
										r_sys_run_phase <= 6'h21;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h27;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp933) ? 6'h2b : 6'h31);

									end
								end

							endcase
						end

						6'h28: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h27;

									end
								end

							endcase
						end

						6'h2b: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h2c;

									end
								end

							endcase
						end

						6'h2c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp938) ? 6'h2f : 6'h28);

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hec)) begin
										r_sys_run_phase <= 6'h2c;

									end
								end

							endcase
						end

						6'h31: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h32;

									end
								end

							endcase
						end

						6'h32: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2464) ? 6'h36 : 6'h11);

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h32;

									end
								end

							endcase
						end

						6'h36: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h37;

									end
								end

							endcase
						end

						6'h37: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2469) ? 6'h3a : 6'h33);

									end
								end

							endcase
						end

						6'h3a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h14)) begin
										r_sys_run_phase <= 6'h37;

									end
								end

							endcase
						end

						6'h3c: begin
							r_sys_run_phase <= 6'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h44)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h25)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h25)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h25)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h12)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h28: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h2b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h2c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hec)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h31: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h32: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h36: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h37: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h3a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h14)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 8'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h43)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==8'h44)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h1) || (r_sys_run_step==8'h2)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h25)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h24)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h25)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h24)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h24)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h12)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h11)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h28: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h2b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h2c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hec)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'heb)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h31: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h32: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h36: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h37: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h3a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h13)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						6'h3c: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_T_0_addr_1 <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h12)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp22[9:0] );

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp571[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp575[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp567[9:0] );

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h1) || (r_sys_run_step==8'h3) || (r_sys_run_step==8'h5) || (r_sys_run_step==8'h7) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h25)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp589[9:0] );

									end
									else
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h2) || (r_sys_run_step==8'h4) || (r_sys_run_step==8'h6) || (r_sys_run_step==8'h8) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h24)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp584[9:0] );

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h12)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp819[9:0] );

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h1) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h43) || (r_sys_run_step==8'h4e) || (r_sys_run_step==8'h59) || (r_sys_run_step==8'h64) || (r_sys_run_step==8'h6f) || (r_sys_run_step==8'h7a) || (r_sys_run_step==8'h85) || (r_sys_run_step==8'h90) || (r_sys_run_step==8'h9b) || (r_sys_run_step==8'ha6) || (r_sys_run_step==8'hb1) || (r_sys_run_step==8'hbc) || (r_sys_run_step==8'hc7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp954[9:0] );

									end
									else
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h3e) || (r_sys_run_step==8'h49) || (r_sys_run_step==8'h54) || (r_sys_run_step==8'h5f) || (r_sys_run_step==8'h6a) || (r_sys_run_step==8'h75) || (r_sys_run_step==8'h80) || (r_sys_run_step==8'h8b) || (r_sys_run_step==8'h96) || (r_sys_run_step==8'ha1) || (r_sys_run_step==8'hac) || (r_sys_run_step==8'hb7) || (r_sys_run_step==8'hc2) || (r_sys_run_step==8'hcd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp985[9:0] );

									end
									else
									if((r_sys_run_step==8'h6) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h32) || (r_sys_run_step==8'h3d) || (r_sys_run_step==8'h48) || (r_sys_run_step==8'h53) || (r_sys_run_step==8'h5e) || (r_sys_run_step==8'h69) || (r_sys_run_step==8'h74) || (r_sys_run_step==8'h7f) || (r_sys_run_step==8'h8a) || (r_sys_run_step==8'h95) || (r_sys_run_step==8'ha0) || (r_sys_run_step==8'hab) || (r_sys_run_step==8'hb6) || (r_sys_run_step==8'hc1) || (r_sys_run_step==8'hcc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp982[9:0] );

									end
									else
									if((r_sys_run_step==8'h4) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h3b) || (r_sys_run_step==8'h46) || (r_sys_run_step==8'h51) || (r_sys_run_step==8'h5c) || (r_sys_run_step==8'h67) || (r_sys_run_step==8'h72) || (r_sys_run_step==8'h7d) || (r_sys_run_step==8'h88) || (r_sys_run_step==8'h93) || (r_sys_run_step==8'h9e) || (r_sys_run_step==8'ha9) || (r_sys_run_step==8'hb4) || (r_sys_run_step==8'hbf) || (r_sys_run_step==8'hca)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp971[9:0] );

									end
									else
									if((r_sys_run_step==8'h5) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h3c) || (r_sys_run_step==8'h47) || (r_sys_run_step==8'h52) || (r_sys_run_step==8'h5d) || (r_sys_run_step==8'h68) || (r_sys_run_step==8'h73) || (r_sys_run_step==8'h7e) || (r_sys_run_step==8'h89) || (r_sys_run_step==8'h94) || (r_sys_run_step==8'h9f) || (r_sys_run_step==8'haa) || (r_sys_run_step==8'hb5) || (r_sys_run_step==8'hc0) || (r_sys_run_step==8'hcb)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp975[9:0] );

									end
									else
									if((r_sys_run_step==8'h3) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h2f) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h45) || (r_sys_run_step==8'h50) || (r_sys_run_step==8'h5b) || (r_sys_run_step==8'h66) || (r_sys_run_step==8'h71) || (r_sys_run_step==8'h7c) || (r_sys_run_step==8'h87) || (r_sys_run_step==8'h92) || (r_sys_run_step==8'h9d) || (r_sys_run_step==8'ha8) || (r_sys_run_step==8'hb3) || (r_sys_run_step==8'hbe) || (r_sys_run_step==8'hc9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp966[9:0] );

									end
									else
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h2c) || (r_sys_run_step==8'h37) || (r_sys_run_step==8'h42) || (r_sys_run_step==8'h4d) || (r_sys_run_step==8'h58) || (r_sys_run_step==8'h63) || (r_sys_run_step==8'h6e) || (r_sys_run_step==8'h79) || (r_sys_run_step==8'h84) || (r_sys_run_step==8'h8f) || (r_sys_run_step==8'h9a) || (r_sys_run_step==8'ha5) || (r_sys_run_step==8'hb0) || (r_sys_run_step==8'hbb) || (r_sys_run_step==8'hc6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp947[9:0] );

									end
									else
									if((r_sys_run_step==8'h9) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h40) || (r_sys_run_step==8'h4b) || (r_sys_run_step==8'h56) || (r_sys_run_step==8'h61) || (r_sys_run_step==8'h6c) || (r_sys_run_step==8'h77) || (r_sys_run_step==8'h82) || (r_sys_run_step==8'h8d) || (r_sys_run_step==8'h98) || (r_sys_run_step==8'ha3) || (r_sys_run_step==8'hae) || (r_sys_run_step==8'hb9) || (r_sys_run_step==8'hc4) || (r_sys_run_step==8'hcf)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp997[9:0] );

									end
									else
									if((r_sys_run_step==8'ha) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h41) || (r_sys_run_step==8'h4c) || (r_sys_run_step==8'h57) || (r_sys_run_step==8'h62) || (r_sys_run_step==8'h6d) || (r_sys_run_step==8'h78) || (r_sys_run_step==8'h83) || (r_sys_run_step==8'h8e) || (r_sys_run_step==8'h99) || (r_sys_run_step==8'ha4) || (r_sys_run_step==8'haf) || (r_sys_run_step==8'hba) || (r_sys_run_step==8'hc5) || (r_sys_run_step==8'hd0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1000[9:0] );

									end
									else
									if((r_sys_run_step==8'h2) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h44) || (r_sys_run_step==8'h4f) || (r_sys_run_step==8'h5a) || (r_sys_run_step==8'h65) || (r_sys_run_step==8'h70) || (r_sys_run_step==8'h7b) || (r_sys_run_step==8'h86) || (r_sys_run_step==8'h91) || (r_sys_run_step==8'h9c) || (r_sys_run_step==8'ha7) || (r_sys_run_step==8'hb2) || (r_sys_run_step==8'hbd) || (r_sys_run_step==8'hc8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp959[9:0] );

									end
									else
									if((r_sys_run_step==8'h8) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h3f) || (r_sys_run_step==8'h4a) || (r_sys_run_step==8'h55) || (r_sys_run_step==8'h60) || (r_sys_run_step==8'h6b) || (r_sys_run_step==8'h76) || (r_sys_run_step==8'h81) || (r_sys_run_step==8'h8c) || (r_sys_run_step==8'h97) || (r_sys_run_step==8'ha2) || (r_sys_run_step==8'had) || (r_sys_run_step==8'hb8) || (r_sys_run_step==8'hc3) || (r_sys_run_step==8'hce)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp991[9:0] );

									end
								end

							endcase
						end

						6'h3a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h14)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2474[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h12)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp25;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp574;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp569;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h25)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp587;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h12)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp822;

									end
								end

							endcase
						end

						6'h3a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h14)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp2477;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_T_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h12)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h3)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h25)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h12)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'hd0)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h14)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h3c: begin
							r_fld_T_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_TT_1_addr_1 <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h12)) begin
										r_fld_TT_1_addr_1 <= $signed( w_sys_tmp27[9:0] );

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h47) || (r_sys_run_step==8'h52) || (r_sys_run_step==8'h53) || (r_sys_run_step==8'h5d) || (r_sys_run_step==8'h5e) || (r_sys_run_step==8'h68) || (r_sys_run_step==8'h73) || (r_sys_run_step==8'h7e) || (r_sys_run_step==8'h89) || (r_sys_run_step==8'h94) || (r_sys_run_step==8'h9f) || (r_sys_run_step==8'haa) || (r_sys_run_step==8'hb5) || (r_sys_run_step==8'hc0) || (r_sys_run_step==8'hcb) || (r_sys_run_step==8'hd6) || (r_sys_run_step==8'hda) || (r_sys_run_step==8'he4) || (r_sys_run_step==8'hec)) begin
										r_fld_TT_1_addr_1 <= $signed( w_sys_tmp943[9:0] );

									end
								end

							endcase
						end

						6'h3a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h12)) begin
										r_fld_TT_1_addr_1 <= $signed( w_sys_tmp2478[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h12)) begin
										r_fld_TT_1_datain_1 <= w_sys_tmp25;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h47) || (r_sys_run_step==8'h52) || (r_sys_run_step==8'h53) || (r_sys_run_step==8'h5d) || (r_sys_run_step==8'h5e) || (r_sys_run_step==8'h68) || (r_sys_run_step==8'h73) || (r_sys_run_step==8'h7e) || (r_sys_run_step==8'h89) || (r_sys_run_step==8'h94) || (r_sys_run_step==8'h9f) || (r_sys_run_step==8'haa) || (r_sys_run_step==8'hb5) || (r_sys_run_step==8'hc0) || (r_sys_run_step==8'hcb) || (r_sys_run_step==8'hd6) || (r_sys_run_step==8'hda) || (r_sys_run_step==8'he4) || (r_sys_run_step==8'hec)) begin
										r_fld_TT_1_datain_1 <= w_sys_tmp946;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_TT_1_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h12)) begin
										r_fld_TT_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h47) || (r_sys_run_step==8'h52) || (r_sys_run_step==8'h53) || (r_sys_run_step==8'h5d) || (r_sys_run_step==8'h5e) || (r_sys_run_step==8'h68) || (r_sys_run_step==8'h73) || (r_sys_run_step==8'h7e) || (r_sys_run_step==8'h89) || (r_sys_run_step==8'h94) || (r_sys_run_step==8'h9f) || (r_sys_run_step==8'haa) || (r_sys_run_step==8'hb5) || (r_sys_run_step==8'hc0) || (r_sys_run_step==8'hcb) || (r_sys_run_step==8'hd6) || (r_sys_run_step==8'hda) || (r_sys_run_step==8'he4) || (r_sys_run_step==8'hec)) begin
										r_fld_TT_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h3a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h12)) begin
										r_fld_TT_1_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3c: begin
							r_fld_TT_1_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_U_2_addr_1 <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h1b) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h3c) || (r_sys_run_step==8'h3e) || (8'h40<=r_sys_run_step && r_sys_run_step<=8'h44)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp32[9:0] );

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h12)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp951[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h1b) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h3c) || (r_sys_run_step==8'h3e) || (8'h40<=r_sys_run_step && r_sys_run_step<=8'h44)) begin
										r_fld_U_2_datain_1 <= w_sys_tmp18;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_U_2_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h1b) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h3c) || (r_sys_run_step==8'h3e) || (8'h40<=r_sys_run_step && r_sys_run_step<=8'h44)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h12)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3c: begin
							r_fld_U_2_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_V_3_addr_1 <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h12)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp41[9:0] );

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h12)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp963[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h12)) begin
										r_fld_V_3_datain_1 <= w_sys_tmp25;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_V_3_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h12)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h12)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3c: begin
							r_fld_V_3_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_4 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_4 <= w_sys_tmp14;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_4 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_run_k_4 <= w_sys_tmp579;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_4 <= w_sys_tmp932;

									end
								end

							endcase
						end

						6'h28: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_4 <= w_sys_tmp936;

									end
								end

							endcase
						end

						6'h31: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_4 <= w_sys_tmp2463;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_4 <= w_sys_tmp2467;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_j_5 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h12)) begin
										r_run_j_5 <= w_sys_tmp48;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_j_5 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h2) || (r_sys_run_step==8'h4) || (r_sys_run_step==8'h6) || (r_sys_run_step==8'h8) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h24)) begin
										r_run_j_5 <= w_sys_tmp594;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h25)) begin
										r_run_j_5 <= w_sys_tmp811;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h12)) begin
										r_run_j_5 <= w_sys_tmp823;

									end
								end

							endcase
						end

						6'h2b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_j_5 <= w_sys_tmp937;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h47) || (r_sys_run_step==8'h52) || (r_sys_run_step==8'h53) || (r_sys_run_step==8'h5d) || (r_sys_run_step==8'h5e) || (r_sys_run_step==8'h68) || (r_sys_run_step==8'h73) || (r_sys_run_step==8'h7e) || (r_sys_run_step==8'h89) || (r_sys_run_step==8'h94) || (r_sys_run_step==8'h9f) || (r_sys_run_step==8'haa) || (r_sys_run_step==8'hb5) || (r_sys_run_step==8'hc0) || (r_sys_run_step==8'hcb) || (r_sys_run_step==8'hd6) || (r_sys_run_step==8'hda) || (r_sys_run_step==8'he4) || (r_sys_run_step==8'hec)) begin
										r_run_j_5 <= w_sys_tmp1017;

									end
								end

							endcase
						end

						6'h36: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_j_5 <= w_sys_tmp2468;

									end
								end

							endcase
						end

						6'h3a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h14)) begin
										r_run_j_5 <= w_sys_tmp2482;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_n_6 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_n_6 <= w_sys_tmp562;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_mx_7 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_my_8 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_dt_9 <= w_sys_tmp5;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_dx_10 <= w_sys_tmp6;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_dy_11 <= w_sys_tmp7;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_r1_12 <= w_sys_tmp8;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_r2_13 <= w_sys_tmp9;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_r3_14 <= w_sys_tmp10;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_r4_15 <= w_sys_tmp11;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h1e) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h36)) begin
										r_run_YY_16 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_run_YY_16 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==8'h21) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h32)) begin
										r_run_YY_16 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_run_YY_16 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==8'h15) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h34)) begin
										r_run_YY_16 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==8'hc) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'he)) begin
										r_run_YY_16 <= w_sys_tmp18;

									end
									else
									if((r_sys_run_step==8'h13) || (r_sys_run_step==8'h38)) begin
										r_run_YY_16 <= r_sys_tmp15_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_kx_17 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_ky_18 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_nlast_19 <= w_sys_intOne;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy0_j_20 <= r_run_j_5;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h12)) begin
										r_run_copy0_j_20 <= w_sys_tmp45;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy1_j_21 <= r_run_j_5;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h1b) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h3c) || (r_sys_run_step==8'h3e) || (8'h40<=r_sys_run_step && r_sys_run_step<=8'h44)) begin
										r_run_copy1_j_21 <= w_sys_tmp46;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy2_j_22 <= r_run_j_5;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h12)) begin
										r_run_copy2_j_22 <= w_sys_tmp47;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1a: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy0_j_23 <= r_run_j_5;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h1) || (r_sys_run_step==8'h3) || (r_sys_run_step==8'h5) || (r_sys_run_step==8'h7) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h25)) begin
										r_run_copy0_j_23 <= w_sys_tmp593;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2b: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy0_j_24 <= r_run_j_5;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'ha) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h41) || (r_sys_run_step==8'h4c) || (r_sys_run_step==8'h57) || (r_sys_run_step==8'h62) || (r_sys_run_step==8'h6d) || (r_sys_run_step==8'h78) || (r_sys_run_step==8'h83) || (r_sys_run_step==8'h8e) || (r_sys_run_step==8'h99) || (r_sys_run_step==8'ha4) || (r_sys_run_step==8'haf) || (r_sys_run_step==8'hba) || (r_sys_run_step==8'hc5) || (r_sys_run_step==8'hd0)) begin
										r_run_copy0_j_24 <= w_sys_tmp1004;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2b: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy1_j_25 <= r_run_j_5;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h9) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h40) || (r_sys_run_step==8'h4b) || (r_sys_run_step==8'h56) || (r_sys_run_step==8'h61) || (r_sys_run_step==8'h6c) || (r_sys_run_step==8'h77) || (r_sys_run_step==8'h82) || (r_sys_run_step==8'h8d) || (r_sys_run_step==8'h98) || (r_sys_run_step==8'ha3) || (r_sys_run_step==8'hae) || (r_sys_run_step==8'hb9) || (r_sys_run_step==8'hc4) || (r_sys_run_step==8'hcf)) begin
										r_run_copy1_j_25 <= w_sys_tmp1005;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2b: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy2_j_26 <= r_run_j_5;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h8) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h3f) || (r_sys_run_step==8'h4a) || (r_sys_run_step==8'h55) || (r_sys_run_step==8'h60) || (r_sys_run_step==8'h6b) || (r_sys_run_step==8'h76) || (r_sys_run_step==8'h81) || (r_sys_run_step==8'h8c) || (r_sys_run_step==8'h97) || (r_sys_run_step==8'ha2) || (r_sys_run_step==8'had) || (r_sys_run_step==8'hb8) || (r_sys_run_step==8'hc3) || (r_sys_run_step==8'hce)) begin
										r_run_copy2_j_26 <= w_sys_tmp1006;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2b: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy3_j_27 <= r_run_j_5;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h3e) || (r_sys_run_step==8'h49) || (r_sys_run_step==8'h54) || (r_sys_run_step==8'h5f) || (r_sys_run_step==8'h6a) || (r_sys_run_step==8'h75) || (r_sys_run_step==8'h80) || (r_sys_run_step==8'h8b) || (r_sys_run_step==8'h96) || (r_sys_run_step==8'ha1) || (r_sys_run_step==8'hac) || (r_sys_run_step==8'hb7) || (r_sys_run_step==8'hc2) || (r_sys_run_step==8'hcd)) begin
										r_run_copy3_j_27 <= w_sys_tmp1007;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2b: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy4_j_28 <= r_run_j_5;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h6) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h32) || (r_sys_run_step==8'h3d) || (r_sys_run_step==8'h48) || (r_sys_run_step==8'h53) || (r_sys_run_step==8'h5e) || (r_sys_run_step==8'h69) || (r_sys_run_step==8'h74) || (r_sys_run_step==8'h7f) || (r_sys_run_step==8'h8a) || (r_sys_run_step==8'h95) || (r_sys_run_step==8'ha0) || (r_sys_run_step==8'hab) || (r_sys_run_step==8'hb6) || (r_sys_run_step==8'hc1) || (r_sys_run_step==8'hcc)) begin
										r_run_copy4_j_28 <= w_sys_tmp1008;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2b: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy5_j_29 <= r_run_j_5;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h5) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h3c) || (r_sys_run_step==8'h47) || (r_sys_run_step==8'h52) || (r_sys_run_step==8'h5d) || (r_sys_run_step==8'h68) || (r_sys_run_step==8'h73) || (r_sys_run_step==8'h7e) || (r_sys_run_step==8'h89) || (r_sys_run_step==8'h94) || (r_sys_run_step==8'h9f) || (r_sys_run_step==8'haa) || (r_sys_run_step==8'hb5) || (r_sys_run_step==8'hc0) || (r_sys_run_step==8'hcb)) begin
										r_run_copy5_j_29 <= w_sys_tmp977;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2b: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy6_j_30 <= r_run_j_5;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h4) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h3b) || (r_sys_run_step==8'h46) || (r_sys_run_step==8'h51) || (r_sys_run_step==8'h5c) || (r_sys_run_step==8'h67) || (r_sys_run_step==8'h72) || (r_sys_run_step==8'h7d) || (r_sys_run_step==8'h88) || (r_sys_run_step==8'h93) || (r_sys_run_step==8'h9e) || (r_sys_run_step==8'ha9) || (r_sys_run_step==8'hb4) || (r_sys_run_step==8'hbf) || (r_sys_run_step==8'hca)) begin
										r_run_copy6_j_30 <= w_sys_tmp1010;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2b: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy7_j_31 <= r_run_j_5;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h3) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h2f) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h45) || (r_sys_run_step==8'h50) || (r_sys_run_step==8'h5b) || (r_sys_run_step==8'h66) || (r_sys_run_step==8'h71) || (r_sys_run_step==8'h7c) || (r_sys_run_step==8'h87) || (r_sys_run_step==8'h92) || (r_sys_run_step==8'h9d) || (r_sys_run_step==8'ha8) || (r_sys_run_step==8'hb3) || (r_sys_run_step==8'hbe) || (r_sys_run_step==8'hc9)) begin
										r_run_copy7_j_31 <= w_sys_tmp1011;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2b: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy8_j_32 <= r_run_j_5;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h12)) begin
										r_run_copy8_j_32 <= w_sys_tmp1012;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2b: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy9_j_33 <= r_run_j_5;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h2) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h44) || (r_sys_run_step==8'h4f) || (r_sys_run_step==8'h5a) || (r_sys_run_step==8'h65) || (r_sys_run_step==8'h70) || (r_sys_run_step==8'h7b) || (r_sys_run_step==8'h86) || (r_sys_run_step==8'h91) || (r_sys_run_step==8'h9c) || (r_sys_run_step==8'ha7) || (r_sys_run_step==8'hb2) || (r_sys_run_step==8'hbd) || (r_sys_run_step==8'hc8)) begin
										r_run_copy9_j_33 <= w_sys_tmp1013;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2b: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy10_j_34 <= r_run_j_5;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h1) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h43) || (r_sys_run_step==8'h4e) || (r_sys_run_step==8'h59) || (r_sys_run_step==8'h64) || (r_sys_run_step==8'h6f) || (r_sys_run_step==8'h7a) || (r_sys_run_step==8'h85) || (r_sys_run_step==8'h90) || (r_sys_run_step==8'h9b) || (r_sys_run_step==8'ha6) || (r_sys_run_step==8'hb1) || (r_sys_run_step==8'hbc) || (r_sys_run_step==8'hc7)) begin
										r_run_copy10_j_34 <= w_sys_tmp956;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2b: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy11_j_35 <= r_run_j_5;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h12)) begin
										r_run_copy11_j_35 <= w_sys_tmp1015;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2b: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy12_j_36 <= r_run_j_5;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h2c) || (r_sys_run_step==8'h37) || (r_sys_run_step==8'h42) || (r_sys_run_step==8'h4d) || (r_sys_run_step==8'h58) || (r_sys_run_step==8'h63) || (r_sys_run_step==8'h6e) || (r_sys_run_step==8'h79) || (r_sys_run_step==8'h84) || (r_sys_run_step==8'h8f) || (r_sys_run_step==8'h9a) || (r_sys_run_step==8'ha5) || (r_sys_run_step==8'hb0) || (r_sys_run_step==8'hbb) || (r_sys_run_step==8'hc6)) begin
										r_run_copy12_j_36 <= w_sys_tmp1016;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h36: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy0_j_37 <= r_run_j_5;

									end
								end

							endcase
						end

						6'h3a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h12)) begin
										r_run_copy0_j_37 <= w_sys_tmp2481;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h18)) begin
										r_sys_tmp0_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h25)) begin
										r_sys_tmp0_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h16)) begin
										r_sys_tmp1_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h20)) begin
										r_sys_tmp1_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h15)) begin
										r_sys_tmp2_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h16)) begin
										r_sys_tmp2_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h13)) begin
										r_sys_tmp3_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h14)) begin
										r_sys_tmp3_float <= w_fld_U_2_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h11) || (r_sys_run_step==8'h17)) begin
										r_sys_tmp4_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h14)) begin
										r_sys_tmp4_float <= w_fld_V_3_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h19) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h2a)) begin
										r_sys_tmp5_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h13)) begin
										r_sys_tmp5_float <= w_fld_V_3_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h18) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h2f)) begin
										r_sys_tmp6_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h12)) begin
										r_sys_tmp6_float <= w_fld_U_2_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'he) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h14)) begin
										r_sys_tmp7_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h11)) begin
										r_sys_tmp7_float <= w_fld_V_3_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h17) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h30)) begin
										r_sys_tmp8_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hf)) begin
										r_sys_tmp8_float <= w_fld_V_3_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h13) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h37)) begin
										r_sys_tmp9_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hd)) begin
										r_sys_tmp9_float <= w_fld_V_3_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h14) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h32)) begin
										r_sys_tmp10_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h17) || (r_sys_run_step==8'h3b)) begin
										r_sys_tmp10_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hc) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h19)) begin
										r_sys_tmp11_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h15) || (r_sys_run_step==8'h2d)) begin
										r_sys_tmp11_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h12) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h32) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h3d)) begin
										r_sys_tmp12_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h13) || (r_sys_run_step==8'h22)) begin
										r_sys_tmp12_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h12) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h37)) begin
										r_sys_tmp13_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'he) || (r_sys_run_step==8'h40)) begin
										r_sys_tmp13_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h11) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h2c) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h3b)) begin
										r_sys_tmp14_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hc) || (r_sys_run_step==8'h1a)) begin
										r_sys_tmp14_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h10) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h2c) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h3b)) begin
										r_sys_tmp15_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h33)) begin
										r_sys_tmp15_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_sys_tmp15_float <= w_fld_U_2_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hf) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h2f) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h3d)) begin
										r_sys_tmp16_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h2c)) begin
										r_sys_tmp16_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_sys_tmp16_float <= w_fld_V_3_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h2b)) begin
										r_sys_tmp17_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_sys_tmp17_float <= w_fld_V_3_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h28)) begin
										r_sys_tmp18_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_sys_tmp18_float <= w_fld_V_3_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h25)) begin
										r_sys_tmp19_float <= w_ip_AddFloat_result_0;

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_sys_tmp19_float <= w_fld_V_3_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h11) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h43)) begin
										r_sys_tmp20_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hb) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h37)) begin
										r_sys_tmp21_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h2e) || (r_sys_run_step==8'h3c)) begin
										r_sys_tmp22_float <= w_ip_AddFloat_result_0;

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_sys_tmp22_float <= w_fld_U_2_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h27) || (r_sys_run_step==8'h29)) begin
										r_sys_tmp23_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_sys_tmp23_float <= w_fld_U_2_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h1d) || (r_sys_run_step==8'h1e)) begin
										r_sys_tmp24_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_sys_tmp24_float <= w_fld_U_2_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h3e)) begin
										r_sys_tmp25_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==8'h5) || (r_sys_run_step==8'h10)) begin
										r_sys_tmp25_float <= w_fld_V_3_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h16) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h3d)) begin
										r_sys_tmp26_float <= w_ip_AddFloat_result_0;

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_sys_tmp26_float <= w_fld_U_2_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h48) || (r_sys_run_step==8'h4a)) begin
										r_sys_tmp27_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==8'ha) || (r_sys_run_step==8'h11)) begin
										r_sys_tmp27_float <= w_fld_U_2_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h46) || (r_sys_run_step==8'h4d)) begin
										r_sys_tmp28_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==8'h6) || (r_sys_run_step==8'h12)) begin
										r_sys_tmp28_float <= w_fld_V_3_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h32) || (r_sys_run_step==8'h34)) begin
										r_sys_tmp29_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==8'h4) || (r_sys_run_step==8'he)) begin
										r_sys_tmp29_float <= w_fld_V_3_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h30) || (r_sys_run_step==8'h36)) begin
										r_sys_tmp30_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==8'h3) || (r_sys_run_step==8'hc)) begin
										r_sys_tmp30_float <= w_fld_V_3_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h23) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h45)) begin
										r_sys_tmp31_float <= w_ip_AddFloat_result_0;

									end
									else
									if((r_sys_run_step==8'h8) || (r_sys_run_step==8'hd)) begin
										r_sys_tmp31_float <= w_fld_U_2_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h3d) || (r_sys_run_step==8'h3f) || (r_sys_run_step==8'h41)) begin
										r_sys_tmp32_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'hf)) begin
										r_sys_tmp32_float <= w_fld_U_2_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h49) || (r_sys_run_step==8'h4c)) begin
										r_sys_tmp33_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==8'h26) || (r_sys_run_step==8'h3b)) begin
										r_sys_tmp33_float <= w_ip_AddFloat_result_0;

									end
									else
									if((r_sys_run_step==8'h2) || (r_sys_run_step==8'h7)) begin
										r_sys_tmp33_float <= w_fld_V_3_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hf) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h4b) || (r_sys_run_step==8'h53) || (r_sys_run_step==8'h5f) || (r_sys_run_step==8'h6a)) begin
										r_sys_tmp34_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h9) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h4e) || (r_sys_run_step==8'h5e) || (r_sys_run_step==8'h61) || (r_sys_run_step==8'h75) || (r_sys_run_step==8'h80) || (r_sys_run_step==8'h8b) || (r_sys_run_step==8'h96) || (r_sys_run_step==8'ha1) || (r_sys_run_step==8'hac) || (r_sys_run_step==8'hb7) || (r_sys_run_step==8'hc2) || (r_sys_run_step==8'hcd)) begin
										r_sys_tmp35_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h8) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h56) || (r_sys_run_step==8'h69) || (r_sys_run_step==8'h6c) || (r_sys_run_step==8'h7f) || (r_sys_run_step==8'h82) || (r_sys_run_step==8'h95) || (r_sys_run_step==8'h98) || (r_sys_run_step==8'hab) || (r_sys_run_step==8'hae) || (r_sys_run_step==8'hc1) || (r_sys_run_step==8'hc4) || (r_sys_run_step==8'hd8)) begin
										r_sys_tmp36_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h74) || (r_sys_run_step==8'h77) || (r_sys_run_step==8'h8a) || (r_sys_run_step==8'h8d) || (r_sys_run_step==8'ha0) || (r_sys_run_step==8'ha3) || (r_sys_run_step==8'hb6) || (r_sys_run_step==8'hb9) || (r_sys_run_step==8'hcc) || (r_sys_run_step==8'hcf) || (r_sys_run_step==8'hd7) || (r_sys_run_step==8'hda) || (r_sys_run_step==8'he5)) begin
										r_sys_tmp37_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hc) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h43) || (r_sys_run_step==8'h4e) || (r_sys_run_step==8'h59) || (r_sys_run_step==8'h64) || (r_sys_run_step==8'h6f) || (r_sys_run_step==8'h7a) || (r_sys_run_step==8'h85) || (r_sys_run_step==8'h90) || (r_sys_run_step==8'h9b) || (r_sys_run_step==8'ha6) || (r_sys_run_step==8'hb1) || (r_sys_run_step==8'hbc) || (r_sys_run_step==8'hc7) || (r_sys_run_step==8'hd2)) begin
										r_sys_tmp38_float <= w_fld_T_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h9) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h40) || (r_sys_run_step==8'h4b) || (r_sys_run_step==8'h56) || (r_sys_run_step==8'h61) || (r_sys_run_step==8'h6c) || (r_sys_run_step==8'h77) || (r_sys_run_step==8'h82) || (r_sys_run_step==8'h8d) || (r_sys_run_step==8'h98) || (r_sys_run_step==8'ha3) || (r_sys_run_step==8'hae) || (r_sys_run_step==8'hb9) || (r_sys_run_step==8'hc4) || (r_sys_run_step==8'hcf)) begin
										r_sys_tmp39_float <= w_fld_T_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h54)) begin
										r_sys_tmp40_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==8'ha) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h41) || (r_sys_run_step==8'h4c) || (r_sys_run_step==8'h57) || (r_sys_run_step==8'h62) || (r_sys_run_step==8'h6d) || (r_sys_run_step==8'h78) || (r_sys_run_step==8'h83) || (r_sys_run_step==8'h8e) || (r_sys_run_step==8'h99) || (r_sys_run_step==8'ha4) || (r_sys_run_step==8'haf) || (r_sys_run_step==8'hba) || (r_sys_run_step==8'hc5) || (r_sys_run_step==8'hd0)) begin
										r_sys_tmp40_float <= w_fld_T_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h12) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h46) || (r_sys_run_step==8'h50) || (r_sys_run_step==8'h5b) || (r_sys_run_step==8'h66) || (r_sys_run_step==8'h71) || (r_sys_run_step==8'h7c) || (r_sys_run_step==8'h87) || (r_sys_run_step==8'h92) || (r_sys_run_step==8'h9d) || (r_sys_run_step==8'ha8) || (r_sys_run_step==8'hb3) || (r_sys_run_step==8'hbe) || (r_sys_run_step==8'hc9) || (r_sys_run_step==8'hd4)) begin
										r_sys_tmp41_float <= w_ip_AddFloat_result_0;

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_sys_tmp41_float <= w_fld_T_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h2) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h3c) || (r_sys_run_step==8'h3e) || (r_sys_run_step==8'h44) || (r_sys_run_step==8'h50) || (r_sys_run_step==8'h52) || (r_sys_run_step==8'h54) || (r_sys_run_step==8'h5a) || (r_sys_run_step==8'h66) || (r_sys_run_step==8'h68) || (r_sys_run_step==8'h6a) || (r_sys_run_step==8'h70) || (r_sys_run_step==8'h7c) || (r_sys_run_step==8'h7e) || (r_sys_run_step==8'h80) || (r_sys_run_step==8'h86) || (r_sys_run_step==8'h92) || (r_sys_run_step==8'h94) || (r_sys_run_step==8'h96) || (r_sys_run_step==8'h9c) || (r_sys_run_step==8'ha8) || (r_sys_run_step==8'haa) || (r_sys_run_step==8'hac) || (r_sys_run_step==8'hb2) || (r_sys_run_step==8'hbe) || (r_sys_run_step==8'hc0) || (r_sys_run_step==8'hc2) || (r_sys_run_step==8'hc8)) begin
										r_sys_tmp42_float <= w_fld_T_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h3) || (r_sys_run_step==8'h5) || (r_sys_run_step==8'h7) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h2f) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h45) || (r_sys_run_step==8'h47) || (r_sys_run_step==8'h49) || (r_sys_run_step==8'h4f) || (r_sys_run_step==8'h5b) || (r_sys_run_step==8'h5d) || (r_sys_run_step==8'h5f) || (r_sys_run_step==8'h65) || (r_sys_run_step==8'h71) || (r_sys_run_step==8'h73) || (r_sys_run_step==8'h75) || (r_sys_run_step==8'h7b) || (r_sys_run_step==8'h87) || (r_sys_run_step==8'h89) || (r_sys_run_step==8'h8b) || (r_sys_run_step==8'h91) || (r_sys_run_step==8'h9d) || (r_sys_run_step==8'h9f) || (r_sys_run_step==8'ha1) || (r_sys_run_step==8'ha7) || (r_sys_run_step==8'hb3) || (r_sys_run_step==8'hb5) || (r_sys_run_step==8'hb7) || (r_sys_run_step==8'hbd) || (r_sys_run_step==8'hc9) || (r_sys_run_step==8'hcb) || (r_sys_run_step==8'hcd)) begin
										r_sys_tmp43_float <= w_fld_T_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h9) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h2c) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h37) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h42) || (r_sys_run_step==8'h43) || (r_sys_run_step==8'h44) || (r_sys_run_step==8'h4d) || (r_sys_run_step==8'h4e) || (r_sys_run_step==8'h4f) || (r_sys_run_step==8'h58) || (r_sys_run_step==8'h59) || (r_sys_run_step==8'h5a) || (r_sys_run_step==8'h63) || (r_sys_run_step==8'h64) || (r_sys_run_step==8'h65) || (r_sys_run_step==8'h6e) || (r_sys_run_step==8'h6f) || (r_sys_run_step==8'h70) || (r_sys_run_step==8'h79) || (r_sys_run_step==8'h7a) || (r_sys_run_step==8'h7b) || (r_sys_run_step==8'h84) || (r_sys_run_step==8'h85) || (r_sys_run_step==8'h86) || (r_sys_run_step==8'h8f) || (r_sys_run_step==8'h90) || (r_sys_run_step==8'h91) || (r_sys_run_step==8'h9a) || (r_sys_run_step==8'h9b) || (r_sys_run_step==8'h9c) || (r_sys_run_step==8'ha5) || (r_sys_run_step==8'ha6) || (r_sys_run_step==8'ha7) || (r_sys_run_step==8'hb0) || (r_sys_run_step==8'hb1) || (r_sys_run_step==8'hb2) || (r_sys_run_step==8'hbb) || (r_sys_run_step==8'hbc) || (r_sys_run_step==8'hbd) || (r_sys_run_step==8'hc6) || (r_sys_run_step==8'hc7) || (r_sys_run_step==8'hc8) || (r_sys_run_step==8'hd1) || (r_sys_run_step==8'hd2) || (r_sys_run_step==8'hd3) || (r_sys_run_step==8'hde)) begin
										r_sys_tmp44_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
