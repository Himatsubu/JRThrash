/*
TimeStamp:	2016/5/10		14:30
*/


module c1_test02(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy	
);

	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 5:0] r_sys_run_phase;
	reg         [ 2:0] r_sys_run_stage;
	reg         [ 4:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 2:0] w_sys_run_stage_p1;
	wire        [ 4:0] w_sys_run_step_p1;
	wire signed [ 8:0] w_fld_u_0_addr_0;
	wire        [31:0] w_fld_u_0_datain_0;
	wire        [31:0] w_fld_u_0_dataout_0;
	wire               w_fld_u_0_r_w_0;
	wire               w_fld_u_0_ce_0;
	reg  signed [ 8:0] r_fld_u_0_addr_1;
	reg         [31:0] r_fld_u_0_datain_1;
	wire        [31:0] w_fld_u_0_dataout_1;
	reg                r_fld_u_0_r_w_1;
	wire               w_fld_u_0_ce_1;
	reg  signed [31:0] r_run_k_5;
	reg  signed [31:0] r_run_j_6;
	reg  signed [31:0] r_run_n_7;
	reg  signed [31:0] r_run_mx_8;
	reg  signed [31:0] r_run_my_9;
	reg  signed [31:0] r_run_nlast_10;
	reg         [31:0] r_run_dx_11;
	reg         [31:0] r_run_dy_12;
	reg  signed [31:0] r_run_copy0_j_13;
	reg  signed [31:0] r_run_copy1_j_14;
	reg  signed [31:0] r_run_copy2_j_15;
	reg                r_sub03_run_req;
	wire               w_sub03_run_busy;
	wire signed [ 8:0] w_sub03_u_addr;
	reg  signed [ 8:0] r_sub03_u_addr;
	wire        [31:0] w_sub03_u_datain;
	reg         [31:0] r_sub03_u_datain;
	wire        [31:0] w_sub03_u_dataout;
	wire               w_sub03_u_r_w;
	reg                r_sub03_u_r_w;
	wire signed [ 8:0] w_sub03_result_addr;
	reg  signed [ 8:0] r_sub03_result_addr;
	wire        [31:0] w_sub03_result_datain;
	reg         [31:0] r_sub03_result_datain;
	wire        [31:0] w_sub03_result_dataout;
	wire               w_sub03_result_r_w;
	reg                r_sub03_result_r_w;
	reg                r_sub02_run_req;
	wire               w_sub02_run_busy;
	wire signed [ 8:0] w_sub02_u_addr;
	reg  signed [ 8:0] r_sub02_u_addr;
	wire        [31:0] w_sub02_u_datain;
	reg         [31:0] r_sub02_u_datain;
	wire        [31:0] w_sub02_u_dataout;
	wire               w_sub02_u_r_w;
	reg                r_sub02_u_r_w;
	wire signed [ 8:0] w_sub02_result_addr;
	reg  signed [ 8:0] r_sub02_result_addr;
	wire        [31:0] w_sub02_result_datain;
	reg         [31:0] r_sub02_result_datain;
	wire        [31:0] w_sub02_result_dataout;
	wire               w_sub02_result_r_w;
	reg                r_sub02_result_r_w;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [ 9:0] w_sub01_u_addr;
	reg  signed [ 9:0] r_sub01_u_addr;
	wire        [31:0] w_sub01_u_datain;
	reg         [31:0] r_sub01_u_datain;
	wire        [31:0] w_sub01_u_dataout;
	wire               w_sub01_u_r_w;
	reg                r_sub01_u_r_w;
	wire signed [ 9:0] w_sub01_result_addr;
	reg  signed [ 9:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [ 8:0] w_sub00_u_addr;
	reg  signed [ 8:0] r_sub00_u_addr;
	wire        [31:0] w_sub00_u_datain;
	reg         [31:0] r_sub00_u_datain;
	wire        [31:0] w_sub00_u_dataout;
	wire               w_sub00_u_r_w;
	reg                r_sub00_u_r_w;
	wire signed [ 8:0] w_sub00_result_addr;
	reg  signed [ 8:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	wire signed [31:0] w_sys_tmp1;
	wire        [31:0] w_sys_tmp3;
	wire signed [31:0] w_sys_tmp5;
	wire               w_sys_tmp6;
	wire               w_sys_tmp7;
	wire signed [31:0] w_sys_tmp8;
	wire               w_sys_tmp9;
	wire               w_sys_tmp10;
	wire signed [31:0] w_sys_tmp13;
	wire signed [31:0] w_sys_tmp14;
	wire signed [31:0] w_sys_tmp15;
	wire        [31:0] w_sys_tmp16;
	wire signed [31:0] w_sys_tmp17;
	wire               w_sys_tmp54;
	wire               w_sys_tmp55;
	wire signed [31:0] w_sys_tmp56;
	wire               w_sys_tmp57;
	wire               w_sys_tmp58;
	wire signed [31:0] w_sys_tmp61;
	wire signed [31:0] w_sys_tmp62;
	wire        [31:0] w_sys_tmp63;
	wire signed [31:0] w_sys_tmp65;
	wire signed [31:0] w_sys_tmp66;
	wire        [31:0] w_sys_tmp68;
	wire signed [31:0] w_sys_tmp70;
	wire signed [31:0] w_sys_tmp71;
	wire        [31:0] w_sys_tmp73;
	wire signed [31:0] w_sys_tmp75;
	wire signed [31:0] w_sys_tmp76;
	wire signed [31:0] w_sys_tmp79;
	wire signed [31:0] w_sys_tmp80;
	wire signed [31:0] w_sys_tmp81;
	wire signed [31:0] w_sys_tmp82;
	wire signed [31:0] w_sys_tmp221;
	wire               w_sys_tmp222;
	wire               w_sys_tmp223;
	wire signed [31:0] w_sys_tmp226;
	wire signed [31:0] w_sys_tmp227;
	wire        [31:0] w_sys_tmp228;
	wire signed [31:0] w_sys_tmp232;
	wire signed [31:0] w_sys_tmp233;
	wire signed [31:0] w_sys_tmp238;
	wire signed [31:0] w_sys_tmp239;
	wire signed [31:0] w_sys_tmp244;
	wire signed [31:0] w_sys_tmp245;
	wire signed [31:0] w_sys_tmp250;
	wire signed [31:0] w_sys_tmp251;
	wire signed [31:0] w_sys_tmp256;
	wire signed [31:0] w_sys_tmp257;
	wire signed [31:0] w_sys_tmp274;
	wire signed [31:0] w_sys_tmp275;
	wire signed [31:0] w_sys_tmp280;
	wire signed [31:0] w_sys_tmp281;
	wire signed [31:0] w_sys_tmp286;
	wire signed [31:0] w_sys_tmp287;
	wire signed [31:0] w_sys_tmp292;
	wire signed [31:0] w_sys_tmp293;
	wire signed [31:0] w_sys_tmp298;
	wire signed [31:0] w_sys_tmp299;
	wire signed [31:0] w_sys_tmp303;
	wire               w_sys_tmp304;
	wire               w_sys_tmp305;
	wire signed [31:0] w_sys_tmp306;
	wire signed [31:0] w_sys_tmp309;
	wire signed [31:0] w_sys_tmp310;
	wire        [31:0] w_sys_tmp311;
	wire signed [31:0] w_sys_tmp315;
	wire signed [31:0] w_sys_tmp316;
	wire signed [31:0] w_sys_tmp321;
	wire signed [31:0] w_sys_tmp322;
	wire signed [31:0] w_sys_tmp327;
	wire signed [31:0] w_sys_tmp328;
	wire signed [31:0] w_sys_tmp333;
	wire signed [31:0] w_sys_tmp334;
	wire signed [31:0] w_sys_tmp339;
	wire signed [31:0] w_sys_tmp340;
	wire signed [31:0] w_sys_tmp357;
	wire signed [31:0] w_sys_tmp358;
	wire signed [31:0] w_sys_tmp363;
	wire signed [31:0] w_sys_tmp364;
	wire signed [31:0] w_sys_tmp369;
	wire signed [31:0] w_sys_tmp370;
	wire signed [31:0] w_sys_tmp375;
	wire signed [31:0] w_sys_tmp376;
	wire signed [31:0] w_sys_tmp381;
	wire signed [31:0] w_sys_tmp382;
	wire signed [31:0] w_sys_tmp386;
	wire signed [31:0] w_sys_tmp387;
	wire               w_sys_tmp388;
	wire               w_sys_tmp389;
	wire signed [31:0] w_sys_tmp390;
	wire signed [31:0] w_sys_tmp393;
	wire signed [31:0] w_sys_tmp394;
	wire        [31:0] w_sys_tmp395;
	wire signed [31:0] w_sys_tmp399;
	wire signed [31:0] w_sys_tmp400;
	wire signed [31:0] w_sys_tmp405;
	wire signed [31:0] w_sys_tmp406;
	wire signed [31:0] w_sys_tmp411;
	wire signed [31:0] w_sys_tmp412;
	wire signed [31:0] w_sys_tmp422;
	wire signed [31:0] w_sys_tmp423;
	wire signed [31:0] w_sys_tmp427;
	wire signed [31:0] w_sys_tmp428;
	wire signed [31:0] w_sys_tmp432;
	wire signed [31:0] w_sys_tmp433;
	wire signed [31:0] w_sys_tmp437;
	wire signed [31:0] w_sys_tmp438;
	wire signed [31:0] w_sys_tmp442;
	wire signed [31:0] w_sys_tmp443;
	wire signed [31:0] w_sys_tmp446;
	wire signed [31:0] w_sys_tmp447;
	wire               w_sys_tmp448;
	wire               w_sys_tmp449;
	wire signed [31:0] w_sys_tmp450;
	wire signed [31:0] w_sys_tmp453;
	wire signed [31:0] w_sys_tmp454;
	wire        [31:0] w_sys_tmp455;
	wire signed [31:0] w_sys_tmp459;
	wire signed [31:0] w_sys_tmp460;
	wire signed [31:0] w_sys_tmp465;
	wire signed [31:0] w_sys_tmp466;
	wire signed [31:0] w_sys_tmp471;
	wire signed [31:0] w_sys_tmp472;
	wire signed [31:0] w_sys_tmp482;
	wire signed [31:0] w_sys_tmp483;
	wire signed [31:0] w_sys_tmp487;
	wire signed [31:0] w_sys_tmp488;
	wire signed [31:0] w_sys_tmp492;
	wire signed [31:0] w_sys_tmp493;
	wire signed [31:0] w_sys_tmp497;
	wire signed [31:0] w_sys_tmp498;
	wire signed [31:0] w_sys_tmp502;
	wire signed [31:0] w_sys_tmp503;
	wire signed [31:0] w_sys_tmp506;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 3'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 5'h1);
	assign w_fld_u_0_addr_0 = 9'sh0;
	assign w_fld_u_0_datain_0 = 32'h0;
	assign w_fld_u_0_r_w_0 = 1'h0;
	assign w_fld_u_0_ce_0 = w_sys_ce;
	assign w_fld_u_0_ce_1 = w_sys_ce;
	assign w_sub03_u_addr = ( (|r_sys_processing_methodID) ? r_sub03_u_addr : 9'sh0 ) ;
	assign w_sub03_u_datain = ( (|r_sys_processing_methodID) ? r_sub03_u_datain : 32'h0 ) ;
	assign w_sub03_u_r_w = ( (|r_sys_processing_methodID) ? r_sub03_u_r_w : 1'h0 ) ;
	assign w_sub03_result_addr = ( (|r_sys_processing_methodID) ? r_sub03_result_addr : 9'sh0 ) ;
	assign w_sub03_result_datain = ( (|r_sys_processing_methodID) ? r_sub03_result_datain : 32'h0 ) ;
	assign w_sub03_result_r_w = ( (|r_sys_processing_methodID) ? r_sub03_result_r_w : 1'h0 ) ;
	assign w_sub02_u_addr = ( (|r_sys_processing_methodID) ? r_sub02_u_addr : 9'sh0 ) ;
	assign w_sub02_u_datain = ( (|r_sys_processing_methodID) ? r_sub02_u_datain : 32'h0 ) ;
	assign w_sub02_u_r_w = ( (|r_sys_processing_methodID) ? r_sub02_u_r_w : 1'h0 ) ;
	assign w_sub02_result_addr = ( (|r_sys_processing_methodID) ? r_sub02_result_addr : 9'sh0 ) ;
	assign w_sub02_result_datain = ( (|r_sys_processing_methodID) ? r_sub02_result_datain : 32'h0 ) ;
	assign w_sub02_result_r_w = ( (|r_sys_processing_methodID) ? r_sub02_result_r_w : 1'h0 ) ;
	assign w_sub01_u_addr = ( (|r_sys_processing_methodID) ? r_sub01_u_addr : 10'sh0 ) ;
	assign w_sub01_u_datain = ( (|r_sys_processing_methodID) ? r_sub01_u_datain : 32'h0 ) ;
	assign w_sub01_u_r_w = ( (|r_sys_processing_methodID) ? r_sub01_u_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 10'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub00_u_addr = ( (|r_sys_processing_methodID) ? r_sub00_u_addr : 9'sh0 ) ;
	assign w_sub00_u_datain = ( (|r_sys_processing_methodID) ? r_sub00_u_datain : 32'h0 ) ;
	assign w_sub00_u_r_w = ( (|r_sys_processing_methodID) ? r_sub00_u_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 9'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh0000000b;
	assign w_sys_tmp3 = 32'h3d4ccccd;
	assign w_sys_tmp5 = 32'sh00000190;
	assign w_sys_tmp6 = ( !w_sys_tmp7 );
	assign w_sys_tmp7 = (r_run_my_9 < r_run_k_5);
	assign w_sys_tmp8 = (r_run_k_5 + w_sys_intOne);
	assign w_sys_tmp9 = ( !w_sys_tmp10 );
	assign w_sys_tmp10 = (r_run_mx_8 < r_run_j_6);
	assign w_sys_tmp13 = (w_sys_tmp14 + r_run_k_5);
	assign w_sys_tmp14 = (r_run_j_6 * w_sys_tmp15);
	assign w_sys_tmp15 = 32'sh0000000b;
	assign w_sys_tmp16 = 32'h0;
	assign w_sys_tmp17 = (r_run_j_6 + w_sys_intOne);
	assign w_sys_tmp54 = ( !w_sys_tmp55 );
	assign w_sys_tmp55 = (r_run_nlast_10 < r_run_n_7);
	assign w_sys_tmp56 = (r_run_n_7 + w_sys_intOne);
	assign w_sys_tmp57 = ( !w_sys_tmp58 );
	assign w_sys_tmp58 = (r_run_my_9 < r_run_j_6);
	assign w_sys_tmp61 = (w_sys_tmp62 + r_run_j_6);
	assign w_sys_tmp62 = 32'sh0000000b;
	assign w_sys_tmp63 = 32'h3f000000;
	assign w_sys_tmp65 = (w_sys_tmp66 + r_run_copy2_j_15);
	assign w_sys_tmp66 = (r_run_mx_8 * w_sys_tmp62);
	assign w_sys_tmp68 = 32'h0;
	assign w_sys_tmp70 = (w_sys_tmp71 + w_sys_intOne);
	assign w_sys_tmp71 = (r_run_copy1_j_14 * w_sys_tmp62);
	assign w_sys_tmp73 = 32'h3f800000;
	assign w_sys_tmp75 = (w_sys_tmp76 + r_run_my_9);
	assign w_sys_tmp76 = (r_run_copy0_j_13 * w_sys_tmp62);
	assign w_sys_tmp79 = (r_run_copy0_j_13 + w_sys_intOne);
	assign w_sys_tmp80 = (r_run_copy1_j_14 + w_sys_intOne);
	assign w_sys_tmp81 = (r_run_copy2_j_15 + w_sys_intOne);
	assign w_sys_tmp82 = (r_run_j_6 + w_sys_intOne);
	assign w_sys_tmp221 = 32'sh00000005;
	assign w_sys_tmp222 = ( !w_sys_tmp223 );
	assign w_sys_tmp223 = (r_run_my_9 < r_run_k_5);
	assign w_sys_tmp226 = (w_sys_tmp227 + r_run_k_5);
	assign w_sys_tmp227 = 32'sh0000000b;
	assign w_sys_tmp228 = w_fld_u_0_dataout_1;
	assign w_sys_tmp232 = (w_sys_tmp233 + r_run_k_5);
	assign w_sys_tmp233 = 32'sh00000016;
	assign w_sys_tmp238 = (w_sys_tmp239 + r_run_k_5);
	assign w_sys_tmp239 = 32'sh00000021;
	assign w_sys_tmp244 = (w_sys_tmp245 + r_run_k_5);
	assign w_sys_tmp245 = 32'sh0000002c;
	assign w_sys_tmp250 = (w_sys_tmp251 + r_run_k_5);
	assign w_sys_tmp251 = 32'sh00000037;
	assign w_sys_tmp256 = (w_sys_tmp257 + r_run_k_5);
	assign w_sys_tmp257 = 32'sh00000042;
	assign w_sys_tmp274 = (w_sys_tmp275 + r_run_k_5);
	assign w_sys_tmp275 = 32'sh0000004d;
	assign w_sys_tmp280 = (w_sys_tmp281 + r_run_k_5);
	assign w_sys_tmp281 = 32'sh00000058;
	assign w_sys_tmp286 = (w_sys_tmp287 + r_run_k_5);
	assign w_sys_tmp287 = 32'sh00000063;
	assign w_sys_tmp292 = (w_sys_tmp293 + r_run_k_5);
	assign w_sys_tmp293 = 32'sh0000006e;
	assign w_sys_tmp298 = (w_sys_tmp299 + r_run_k_5);
	assign w_sys_tmp299 = 32'sh00000079;
	assign w_sys_tmp303 = (r_run_k_5 + w_sys_intOne);
	assign w_sys_tmp304 = ( !w_sys_tmp305 );
	assign w_sys_tmp305 = (w_sys_tmp306 < r_run_k_5);
	assign w_sys_tmp306 = 32'sh00000006;
	assign w_sys_tmp309 = (w_sys_tmp310 + r_run_k_5);
	assign w_sys_tmp310 = 32'sh0000000b;
	assign w_sys_tmp311 = w_fld_u_0_dataout_1;
	assign w_sys_tmp315 = (w_sys_tmp316 + r_run_k_5);
	assign w_sys_tmp316 = 32'sh00000016;
	assign w_sys_tmp321 = (w_sys_tmp322 + r_run_k_5);
	assign w_sys_tmp322 = 32'sh00000021;
	assign w_sys_tmp327 = (w_sys_tmp328 + r_run_k_5);
	assign w_sys_tmp328 = 32'sh0000002c;
	assign w_sys_tmp333 = (w_sys_tmp334 + r_run_k_5);
	assign w_sys_tmp334 = 32'sh00000037;
	assign w_sys_tmp339 = (w_sys_tmp340 + r_run_k_5);
	assign w_sys_tmp340 = 32'sh00000042;
	assign w_sys_tmp357 = (w_sys_tmp358 + r_run_k_5);
	assign w_sys_tmp358 = 32'sh0000004d;
	assign w_sys_tmp363 = (w_sys_tmp364 + r_run_k_5);
	assign w_sys_tmp364 = 32'sh00000058;
	assign w_sys_tmp369 = (w_sys_tmp370 + r_run_k_5);
	assign w_sys_tmp370 = 32'sh00000063;
	assign w_sys_tmp375 = (w_sys_tmp376 + r_run_k_5);
	assign w_sys_tmp376 = 32'sh0000006e;
	assign w_sys_tmp381 = (w_sys_tmp382 + r_run_k_5);
	assign w_sys_tmp382 = 32'sh00000079;
	assign w_sys_tmp386 = (r_run_k_5 + w_sys_intOne);
	assign w_sys_tmp387 = 32'sh00000002;
	assign w_sys_tmp388 = ( !w_sys_tmp389 );
	assign w_sys_tmp389 = (w_sys_tmp390 < r_run_k_5);
	assign w_sys_tmp390 = 32'sh00000005;
	assign w_sys_tmp393 = (w_sys_tmp394 + r_run_k_5);
	assign w_sys_tmp394 = 32'sh00000016;
	assign w_sys_tmp395 = w_sub00_result_dataout;
	assign w_sys_tmp399 = (w_sys_tmp400 + r_run_k_5);
	assign w_sys_tmp400 = 32'sh00000021;
	assign w_sys_tmp405 = (w_sys_tmp406 + r_run_k_5);
	assign w_sys_tmp406 = 32'sh0000002c;
	assign w_sys_tmp411 = (w_sys_tmp412 + r_run_k_5);
	assign w_sys_tmp412 = 32'sh00000037;
	assign w_sys_tmp422 = (w_sys_tmp423 + r_run_k_5);
	assign w_sys_tmp423 = 32'sh00000042;
	assign w_sys_tmp427 = (w_sys_tmp428 + r_run_k_5);
	assign w_sys_tmp428 = 32'sh0000004d;
	assign w_sys_tmp432 = (w_sys_tmp433 + r_run_k_5);
	assign w_sys_tmp433 = 32'sh00000058;
	assign w_sys_tmp437 = (w_sys_tmp438 + r_run_k_5);
	assign w_sys_tmp438 = 32'sh00000063;
	assign w_sys_tmp442 = (w_sys_tmp443 + r_run_k_5);
	assign w_sys_tmp443 = 32'sh0000006e;
	assign w_sys_tmp446 = (r_run_k_5 + w_sys_intOne);
	assign w_sys_tmp447 = 32'sh00000006;
	assign w_sys_tmp448 = ( !w_sys_tmp449 );
	assign w_sys_tmp449 = (w_sys_tmp450 < r_run_k_5);
	assign w_sys_tmp450 = 32'sh0000000a;
	assign w_sys_tmp453 = (w_sys_tmp454 + r_run_k_5);
	assign w_sys_tmp454 = 32'sh00000016;
	assign w_sys_tmp455 = w_sub02_result_dataout;
	assign w_sys_tmp459 = (w_sys_tmp460 + r_run_k_5);
	assign w_sys_tmp460 = 32'sh00000021;
	assign w_sys_tmp465 = (w_sys_tmp466 + r_run_k_5);
	assign w_sys_tmp466 = 32'sh0000002c;
	assign w_sys_tmp471 = (w_sys_tmp472 + r_run_k_5);
	assign w_sys_tmp472 = 32'sh00000037;
	assign w_sys_tmp482 = (w_sys_tmp483 + r_run_k_5);
	assign w_sys_tmp483 = 32'sh00000042;
	assign w_sys_tmp487 = (w_sys_tmp488 + r_run_k_5);
	assign w_sys_tmp488 = 32'sh0000004d;
	assign w_sys_tmp492 = (w_sys_tmp493 + r_run_k_5);
	assign w_sys_tmp493 = 32'sh00000058;
	assign w_sys_tmp497 = (w_sys_tmp498 + r_run_k_5);
	assign w_sys_tmp498 = 32'sh00000063;
	assign w_sys_tmp502 = (w_sys_tmp503 + r_run_k_5);
	assign w_sys_tmp503 = 32'sh0000006e;
	assign w_sys_tmp506 = (r_run_k_5 + w_sys_intOne);


	sub03
		sub03_inst(
			.i_fld_result_1_addr_0 (w_sub03_result_addr),
			.i_fld_result_1_datain_0 (w_sub03_result_datain),
			.o_fld_result_1_dataout_0 (w_sub03_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub03_result_r_w),
			.i_fld_u_0_addr_0 (w_sub03_u_addr),
			.i_fld_u_0_datain_0 (w_sub03_u_datain),
			.o_fld_u_0_dataout_0 (w_sub03_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub03_u_r_w),
			.o_run_busy (w_sub03_run_busy),
			.i_run_req (r_sub03_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub02
		sub02_inst(
			.i_fld_result_1_addr_0 (w_sub02_result_addr),
			.i_fld_result_1_datain_0 (w_sub02_result_datain),
			.o_fld_result_1_dataout_0 (w_sub02_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub02_result_r_w),
			.i_fld_u_0_addr_0 (w_sub02_u_addr),
			.i_fld_u_0_datain_0 (w_sub02_u_datain),
			.o_fld_u_0_dataout_0 (w_sub02_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub02_u_r_w),
			.o_run_busy (w_sub02_run_busy),
			.i_run_req (r_sub02_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub01
		sub01_inst(
			.i_fld_result_1_addr_0 (w_sub01_result_addr),
			.i_fld_result_1_datain_0 (w_sub01_result_datain),
			.o_fld_result_1_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub01_result_r_w),
			.i_fld_u_0_addr_0 (w_sub01_u_addr),
			.i_fld_u_0_datain_0 (w_sub01_u_datain),
			.o_fld_u_0_dataout_0 (w_sub01_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub01_u_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub00
		sub00_inst(
			.i_fld_result_1_addr_0 (w_sub00_result_addr),
			.i_fld_result_1_datain_0 (w_sub00_result_datain),
			.o_fld_result_1_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub00_result_r_w),
			.i_fld_u_0_addr_0 (w_sub00_u_addr),
			.i_fld_u_0_datain_0 (w_sub00_u_datain),
			.o_fld_u_0_dataout_0 (w_sub00_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub00_u_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(9), .WORDS(484) )
		dpram_u_0(
			.clk (clock),
			.ce_0 (w_fld_u_0_ce_0),
			.addr_0 (w_fld_u_0_addr_0),
			.datain_0 (w_fld_u_0_datain_0),
			.dataout_0 (w_fld_u_0_dataout_0),
			.r_w_0 (w_fld_u_0_r_w_0),
			.ce_1 (w_fld_u_0_ce_1),
			.addr_1 (r_fld_u_0_addr_1),
			.datain_1 (r_fld_u_0_datain_1),
			.dataout_1 (w_fld_u_0_dataout_1),
			.r_w_1 (r_fld_u_0_r_w_1)
		);

	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h36: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 6'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_phase <= 6'h2;
						end

						6'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 6'h4;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6) ? 6'h9 : 6'hf);

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 6'ha;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp9) ? 6'hd : 6'h6);

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h6)) begin
										r_sys_run_phase <= 6'ha;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 6'h10;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp54) ? 6'h14 : 6'h36);

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 6'h10;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 6'h15;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp57) ? 6'h18 : 6'h1a);

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1b)) begin
										r_sys_run_phase <= 6'h15;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 6'h1b;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp222) ? 6'h1e : 6'h1f);

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'he)) begin
										r_sys_run_phase <= 6'h1b;

									end
								end

							endcase
						end

						6'h1f: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_phase <= 6'h21;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 6'h22;

									end
								end

							endcase
						end

						6'h22: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp304) ? 6'h25 : 6'h26);

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'he)) begin
										r_sys_run_phase <= 6'h22;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_phase <= 6'h28;

									end
								end

							endcase
						end

						6'h28: begin

							case(r_sys_run_stage) 
								3'h3: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_phase <= 6'h2a;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 6'h2b;

									end
								end

							endcase
						end

						6'h2b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp388) ? 6'h2e : 6'h30);

									end
								end

							endcase
						end

						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'hb)) begin
										r_sys_run_phase <= 6'h2b;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 6'h31;

									end
								end

							endcase
						end

						6'h31: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp448) ? 6'h34 : 6'h11);

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'hb)) begin
										r_sys_run_phase <= 6'h31;

									end
								end

							endcase
						end

						6'h36: begin
							r_sys_run_phase <= 6'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 3'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h6)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1b)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'he)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h22: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'he)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h28: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h2b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'hb)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h31: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'hb)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 5'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h6)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h5)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1b)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h1a)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'he)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'hd)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h22: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'he)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'hd)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h28: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub00_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub01_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub02_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub03_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h2b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'ha)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'hb)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h31: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'hb)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'ha)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						6'h36: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_addr_1 <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp13[8:0] );

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h3) || (r_sys_run_step==5'h7) || (r_sys_run_step==5'hb) || (r_sys_run_step==5'hf) || (r_sys_run_step==5'h13) || (r_sys_run_step==5'h17) || (r_sys_run_step==5'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp75[8:0] );

									end
									else
									if((r_sys_run_step==5'h1) || (r_sys_run_step==5'h5) || (r_sys_run_step==5'h9) || (r_sys_run_step==5'hd) || (r_sys_run_step==5'h11) || (r_sys_run_step==5'h15) || (r_sys_run_step==5'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp65[8:0] );

									end
									else
									if((r_sys_run_step==5'h0) || (r_sys_run_step==5'h4) || (r_sys_run_step==5'h8) || (r_sys_run_step==5'hc) || (r_sys_run_step==5'h10) || (r_sys_run_step==5'h14) || (r_sys_run_step==5'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp61[8:0] );

									end
									else
									if((r_sys_run_step==5'h2) || (r_sys_run_step==5'h6) || (r_sys_run_step==5'ha) || (r_sys_run_step==5'he) || (r_sys_run_step==5'h12) || (r_sys_run_step==5'h16) || (r_sys_run_step==5'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp70[8:0] );

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp274[8:0] );

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp226[8:0] );

									end
									else
									if((r_sys_run_step==5'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp298[8:0] );

									end
									else
									if((r_sys_run_step==5'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp244[8:0] );

									end
									else
									if((r_sys_run_step==5'h5) || (r_sys_run_step==5'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp256[8:0] );

									end
									else
									if((r_sys_run_step==5'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp286[8:0] );

									end
									else
									if((r_sys_run_step==5'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp292[8:0] );

									end
									else
									if((r_sys_run_step==5'h4) || (r_sys_run_step==5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp250[8:0] );

									end
									else
									if((r_sys_run_step==5'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp280[8:0] );

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp232[8:0] );

									end
									else
									if((r_sys_run_step==5'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp238[8:0] );

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp369[8:0] );

									end
									else
									if((r_sys_run_step==5'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp363[8:0] );

									end
									else
									if((r_sys_run_step==5'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp381[8:0] );

									end
									else
									if((r_sys_run_step==5'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp375[8:0] );

									end
									else
									if((r_sys_run_step==5'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp327[8:0] );

									end
									else
									if((r_sys_run_step==5'h4) || (r_sys_run_step==5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp333[8:0] );

									end
									else
									if((r_sys_run_step==5'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp321[8:0] );

									end
									else
									if((r_sys_run_step==5'h5) || (r_sys_run_step==5'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp339[8:0] );

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp309[8:0] );

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp357[8:0] );

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp315[8:0] );

									end
								end

							endcase
						end

						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp437[8:0] );

									end
									else
									if((r_sys_run_step==5'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp405[8:0] );

									end
									else
									if((r_sys_run_step==5'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp399[8:0] );

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp427[8:0] );

									end
									else
									if((r_sys_run_step==5'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp422[8:0] );

									end
									else
									if((r_sys_run_step==5'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp442[8:0] );

									end
									else
									if((r_sys_run_step==5'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp432[8:0] );

									end
									else
									if((r_sys_run_step==5'h5) || (r_sys_run_step==5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp411[8:0] );

									end
									else
									if((r_sys_run_step==5'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp393[8:0] );

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp492[8:0] );

									end
									else
									if((r_sys_run_step==5'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp465[8:0] );

									end
									else
									if((r_sys_run_step==5'h5) || (r_sys_run_step==5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp471[8:0] );

									end
									else
									if((r_sys_run_step==5'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp482[8:0] );

									end
									else
									if((r_sys_run_step==5'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp502[8:0] );

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp487[8:0] );

									end
									else
									if((r_sys_run_step==5'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp459[8:0] );

									end
									else
									if((r_sys_run_step==5'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp453[8:0] );

									end
									else
									if((r_sys_run_step==5'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp497[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp16;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h2) || (r_sys_run_step==5'h6) || (r_sys_run_step==5'ha) || (r_sys_run_step==5'he) || (r_sys_run_step==5'h12) || (r_sys_run_step==5'h16) || (r_sys_run_step==5'h1a)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp73;

									end
									else
									if((r_sys_run_step==5'h0) || (r_sys_run_step==5'h4) || (r_sys_run_step==5'h8) || (r_sys_run_step==5'hc) || (r_sys_run_step==5'h10) || (r_sys_run_step==5'h14) || (r_sys_run_step==5'h18)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp63;

									end
									else
									if((r_sys_run_step==5'h1) || (r_sys_run_step==5'h3) || (r_sys_run_step==5'h5) || (r_sys_run_step==5'h7) || (r_sys_run_step==5'h9) || (r_sys_run_step==5'hb) || (r_sys_run_step==5'hd) || (r_sys_run_step==5'hf) || (r_sys_run_step==5'h11) || (r_sys_run_step==5'h13) || (r_sys_run_step==5'h15) || (r_sys_run_step==5'h17) || (r_sys_run_step==5'h19) || (r_sys_run_step==5'h1b)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp68;

									end
								end

							endcase
						end

						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h9)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==5'h6) || (r_sys_run_step==5'ha)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp3_float;

									end
									else
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h5)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp395;

									end
									else
									if((r_sys_run_step==5'h7) || (r_sys_run_step==5'hb)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp1_float;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h9)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==5'h6) || (r_sys_run_step==5'ha)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp3_float;

									end
									else
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h5)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp455;

									end
									else
									if((r_sys_run_step==5'h7) || (r_sys_run_step==5'hb)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp1_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h1b)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'hc)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'hc)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'hb)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'hb)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h36: begin
							r_fld_u_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h4: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_5 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_5 <= w_sys_tmp8;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_5 <= w_sys_tmp221;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'he)) begin
										r_run_k_5 <= w_sys_tmp303;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_5 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'he)) begin
										r_run_k_5 <= w_sys_tmp386;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_5 <= w_sys_tmp387;

									end
								end

							endcase
						end

						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'hb)) begin
										r_run_k_5 <= w_sys_tmp446;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_5 <= w_sys_tmp447;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'hb)) begin
										r_run_k_5 <= w_sys_tmp506;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_6 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_j_6 <= w_sys_tmp17;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_6 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0) || (r_sys_run_step==5'h4) || (r_sys_run_step==5'h8) || (r_sys_run_step==5'hc) || (r_sys_run_step==5'h10) || (r_sys_run_step==5'h14) || (r_sys_run_step==5'h18)) begin
										r_run_j_6 <= w_sys_tmp82;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_n_7 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_n_7 <= w_sys_tmp56;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_mx_8 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_my_9 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_nlast_10 <= w_sys_tmp5;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_dx_11 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_dy_12 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_13 <= r_run_j_6;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h3) || (r_sys_run_step==5'h7) || (r_sys_run_step==5'hb) || (r_sys_run_step==5'hf) || (r_sys_run_step==5'h13) || (r_sys_run_step==5'h17) || (r_sys_run_step==5'h1b)) begin
										r_run_copy0_j_13 <= w_sys_tmp79;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy1_j_14 <= r_run_j_6;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h2) || (r_sys_run_step==5'h6) || (r_sys_run_step==5'ha) || (r_sys_run_step==5'he) || (r_sys_run_step==5'h12) || (r_sys_run_step==5'h16) || (r_sys_run_step==5'h1a)) begin
										r_run_copy1_j_14 <= w_sys_tmp80;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy2_j_15 <= r_run_j_6;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1) || (r_sys_run_step==5'h5) || (r_sys_run_step==5'h9) || (r_sys_run_step==5'hd) || (r_sys_run_step==5'h11) || (r_sys_run_step==5'h15) || (r_sys_run_step==5'h19)) begin
										r_run_copy2_j_15 <= w_sys_tmp81;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1f: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'ha)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp274[8:0] );

									end
									else
									if((r_sys_run_step==5'he)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp298[8:0] );

									end
									else
									if((r_sys_run_step==5'h9)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp256[8:0] );

									end
									else
									if((r_sys_run_step==5'hc)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp286[8:0] );

									end
									else
									if((r_sys_run_step==5'hd)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp292[8:0] );

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp250[8:0] );

									end
									else
									if((r_sys_run_step==5'hb)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp280[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h8<=r_sys_run_step && r_sys_run_step<=5'he)) begin
										r_sub03_u_datain <= w_sys_tmp228;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h8<=r_sys_run_step && r_sys_run_step<=5'he)) begin
										r_sub03_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h36: begin
							r_sub03_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h3)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp492[8:0] );

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp471[8:0] );

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp482[8:0] );

									end
									else
									if((r_sys_run_step==5'h5)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp502[8:0] );

									end
									else
									if((r_sys_run_step==5'h2)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp487[8:0] );

									end
									else
									if((r_sys_run_step==5'h4)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp497[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h5)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h36: begin
							r_sub03_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h2)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp226[8:0] );

									end
									else
									if((r_sys_run_step==5'h5)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp244[8:0] );

									end
									else
									if((r_sys_run_step==5'h7)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp256[8:0] );

									end
									else
									if((r_sys_run_step==5'h6)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp250[8:0] );

									end
									else
									if((r_sys_run_step==5'h3)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp232[8:0] );

									end
									else
									if((r_sys_run_step==5'h4)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp238[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sub02_u_datain <= w_sys_tmp228;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sub02_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h36: begin
							r_sub02_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h2)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp465[8:0] );

									end
									else
									if((r_sys_run_step==5'h3)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp471[8:0] );

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp459[8:0] );

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp453[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h3)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h36: begin
							r_sub02_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h26: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'hc)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp369[9:0] );

									end
									else
									if((r_sys_run_step==5'hb)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp363[9:0] );

									end
									else
									if((r_sys_run_step==5'he)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp381[9:0] );

									end
									else
									if((r_sys_run_step==5'hd)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp375[9:0] );

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp333[9:0] );

									end
									else
									if((r_sys_run_step==5'h9)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp339[9:0] );

									end
									else
									if((r_sys_run_step==5'ha)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp357[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h8<=r_sys_run_step && r_sys_run_step<=5'he)) begin
										r_sub01_u_datain <= w_sys_tmp311;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h8<=r_sys_run_step && r_sys_run_step<=5'he)) begin
										r_sub01_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h36: begin
							r_sub01_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h4)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp437[9:0] );

									end
									else
									if((r_sys_run_step==5'h2)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp427[9:0] );

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp422[9:0] );

									end
									else
									if((r_sys_run_step==5'h5)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp442[9:0] );

									end
									else
									if((r_sys_run_step==5'h3)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp432[9:0] );

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp411[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h5)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h36: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h26: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h5)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp327[8:0] );

									end
									else
									if((r_sys_run_step==5'h6)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp333[8:0] );

									end
									else
									if((r_sys_run_step==5'h4)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp321[8:0] );

									end
									else
									if((r_sys_run_step==5'h7)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp339[8:0] );

									end
									else
									if((r_sys_run_step==5'h2)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp309[8:0] );

									end
									else
									if((r_sys_run_step==5'h3)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp315[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sub00_u_datain <= w_sys_tmp311;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sub00_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h36: begin
							r_sub00_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h2)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp405[8:0] );

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp399[8:0] );

									end
									else
									if((r_sys_run_step==5'h3)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp411[8:0] );

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp393[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h3)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h36: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h5)) begin
										r_sys_tmp0_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h5)) begin
										r_sys_tmp0_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h4)) begin
										r_sys_tmp1_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h4)) begin
										r_sys_tmp1_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h3) || (r_sys_run_step==5'h7)) begin
										r_sys_tmp2_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h3) || (r_sys_run_step==5'h7)) begin
										r_sys_tmp2_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h2) || (r_sys_run_step==5'h6)) begin
										r_sys_tmp3_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h2) || (r_sys_run_step==5'h6)) begin
										r_sys_tmp3_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
