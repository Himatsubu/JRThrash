/*
TimeStamp:	2016/10/5		20:33
*/


module c1(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy	
);

	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 8:0] r_sys_run_phase;
	reg         [ 4:0] r_sys_run_stage;
	reg         [ 5:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 4:0] w_sys_run_stage_p1;
	wire        [ 5:0] w_sys_run_step_p1;
	wire signed [14:0] w_fld_u_0_addr_0;
	wire        [31:0] w_fld_u_0_datain_0;
	wire        [31:0] w_fld_u_0_dataout_0;
	wire               w_fld_u_0_r_w_0;
	wire               w_fld_u_0_ce_0;
	reg  signed [14:0] r_fld_u_0_addr_1;
	reg         [31:0] r_fld_u_0_datain_1;
	wire        [31:0] w_fld_u_0_dataout_1;
	reg                r_fld_u_0_r_w_1;
	wire               w_fld_u_0_ce_1;
	reg  signed [31:0] r_run_k_17;
	reg  signed [31:0] r_run_j_18;
	reg  signed [31:0] r_run_n_19;
	reg  signed [31:0] r_run_mx_20;
	reg  signed [31:0] r_run_my_21;
	reg  signed [31:0] r_run_nlast_22;
	reg  signed [31:0] r_run_copy0_j_23;
	reg  signed [31:0] r_run_copy0_j_24;
	reg  signed [31:0] r_run_copy0_j_25;
	reg  signed [31:0] r_run_copy0_j_26;
	reg  signed [31:0] r_run_copy0_j_27;
	reg  signed [31:0] r_run_copy0_j_28;
	reg  signed [31:0] r_run_copy0_j_29;
	reg  signed [31:0] r_run_copy0_j_30;
	reg  signed [31:0] r_run_copy0_j_31;
	reg  signed [31:0] r_run_copy0_j_32;
	reg  signed [31:0] r_run_copy0_j_33;
	reg  signed [31:0] r_run_copy0_j_34;
	reg  signed [31:0] r_run_copy0_j_35;
	reg  signed [31:0] r_run_copy0_j_36;
	reg  signed [31:0] r_run_copy0_j_37;
	reg  signed [31:0] r_run_copy0_j_38;
	reg  signed [31:0] r_run_copy0_j_39;
	reg  signed [31:0] r_run_copy1_j_40;
	reg  signed [31:0] r_run_copy2_j_41;
	reg  signed [31:0] r_run_copy3_j_42;
	reg  signed [31:0] r_run_copy4_j_43;
	reg  signed [31:0] r_run_copy5_j_44;
	reg  signed [31:0] r_run_copy6_j_45;
	reg  signed [31:0] r_run_copy7_j_46;
	reg  signed [31:0] r_run_copy8_j_47;
	reg  signed [31:0] r_run_copy9_j_48;
	reg  signed [31:0] r_run_copy10_j_49;
	reg  signed [31:0] r_run_copy0_j_50;
	reg  signed [31:0] r_run_copy1_j_51;
	reg  signed [31:0] r_run_copy2_j_52;
	reg  signed [31:0] r_run_copy3_j_53;
	reg  signed [31:0] r_run_copy4_j_54;
	reg  signed [31:0] r_run_copy5_j_55;
	reg  signed [31:0] r_run_copy6_j_56;
	reg  signed [31:0] r_run_copy7_j_57;
	reg  signed [31:0] r_run_copy8_j_58;
	reg  signed [31:0] r_run_copy9_j_59;
	reg  signed [31:0] r_run_copy10_j_60;
	reg  signed [31:0] r_run_copy0_j_61;
	reg  signed [31:0] r_run_copy1_j_62;
	reg  signed [31:0] r_run_copy2_j_63;
	reg  signed [31:0] r_run_copy3_j_64;
	reg  signed [31:0] r_run_copy4_j_65;
	reg  signed [31:0] r_run_copy5_j_66;
	reg  signed [31:0] r_run_copy6_j_67;
	reg  signed [31:0] r_run_copy7_j_68;
	reg  signed [31:0] r_run_copy8_j_69;
	reg  signed [31:0] r_run_copy9_j_70;
	reg  signed [31:0] r_run_copy10_j_71;
	reg  signed [31:0] r_run_copy0_j_72;
	reg  signed [31:0] r_run_copy1_j_73;
	reg  signed [31:0] r_run_copy2_j_74;
	reg  signed [31:0] r_run_copy3_j_75;
	reg  signed [31:0] r_run_copy4_j_76;
	reg  signed [31:0] r_run_copy5_j_77;
	reg  signed [31:0] r_run_copy6_j_78;
	reg  signed [31:0] r_run_copy7_j_79;
	reg  signed [31:0] r_run_copy8_j_80;
	reg  signed [31:0] r_run_copy9_j_81;
	reg  signed [31:0] r_run_copy10_j_82;
	reg  signed [31:0] r_run_copy0_j_83;
	reg  signed [31:0] r_run_copy0_j_84;
	reg  signed [31:0] r_run_copy0_j_85;
	reg  signed [31:0] r_run_copy0_j_86;
	reg  signed [31:0] r_run_copy0_j_87;
	reg  signed [31:0] r_run_copy0_j_88;
	reg  signed [31:0] r_run_copy0_j_89;
	reg  signed [31:0] r_run_copy0_j_90;
	reg  signed [31:0] r_run_copy0_j_91;
	reg  signed [31:0] r_run_copy0_j_92;
	reg  signed [31:0] r_run_copy0_j_93;
	reg  signed [31:0] r_run_copy0_j_94;
	reg  signed [31:0] r_run_copy0_j_95;
	reg  signed [31:0] r_run_copy0_j_96;
	reg  signed [31:0] r_run_copy0_j_97;
	reg  signed [31:0] r_run_copy0_j_98;
	reg                r_sub09_run_req;
	wire               w_sub09_run_busy;
	wire signed [12:0] w_sub09_u_addr;
	reg  signed [12:0] r_sub09_u_addr;
	wire        [31:0] w_sub09_u_datain;
	reg         [31:0] r_sub09_u_datain;
	wire        [31:0] w_sub09_u_dataout;
	wire               w_sub09_u_r_w;
	reg                r_sub09_u_r_w;
	wire signed [12:0] w_sub09_result_addr;
	reg  signed [12:0] r_sub09_result_addr;
	wire        [31:0] w_sub09_result_datain;
	reg         [31:0] r_sub09_result_datain;
	wire        [31:0] w_sub09_result_dataout;
	wire               w_sub09_result_r_w;
	reg                r_sub09_result_r_w;
	reg                r_sub08_run_req;
	wire               w_sub08_run_busy;
	wire signed [12:0] w_sub08_u_addr;
	reg  signed [12:0] r_sub08_u_addr;
	wire        [31:0] w_sub08_u_datain;
	reg         [31:0] r_sub08_u_datain;
	wire        [31:0] w_sub08_u_dataout;
	wire               w_sub08_u_r_w;
	reg                r_sub08_u_r_w;
	wire signed [12:0] w_sub08_result_addr;
	reg  signed [12:0] r_sub08_result_addr;
	wire        [31:0] w_sub08_result_datain;
	reg         [31:0] r_sub08_result_datain;
	wire        [31:0] w_sub08_result_dataout;
	wire               w_sub08_result_r_w;
	reg                r_sub08_result_r_w;
	reg                r_sub12_run_req;
	wire               w_sub12_run_busy;
	wire signed [12:0] w_sub12_u_addr;
	reg  signed [12:0] r_sub12_u_addr;
	wire        [31:0] w_sub12_u_datain;
	reg         [31:0] r_sub12_u_datain;
	wire        [31:0] w_sub12_u_dataout;
	wire               w_sub12_u_r_w;
	reg                r_sub12_u_r_w;
	wire signed [12:0] w_sub12_result_addr;
	reg  signed [12:0] r_sub12_result_addr;
	wire        [31:0] w_sub12_result_datain;
	reg         [31:0] r_sub12_result_datain;
	wire        [31:0] w_sub12_result_dataout;
	wire               w_sub12_result_r_w;
	reg                r_sub12_result_r_w;
	reg                r_sub03_run_req;
	wire               w_sub03_run_busy;
	wire signed [12:0] w_sub03_u_addr;
	reg  signed [12:0] r_sub03_u_addr;
	wire        [31:0] w_sub03_u_datain;
	reg         [31:0] r_sub03_u_datain;
	wire        [31:0] w_sub03_u_dataout;
	wire               w_sub03_u_r_w;
	reg                r_sub03_u_r_w;
	wire signed [12:0] w_sub03_result_addr;
	reg  signed [12:0] r_sub03_result_addr;
	wire        [31:0] w_sub03_result_datain;
	reg         [31:0] r_sub03_result_datain;
	wire        [31:0] w_sub03_result_dataout;
	wire               w_sub03_result_r_w;
	reg                r_sub03_result_r_w;
	reg                r_sub02_run_req;
	wire               w_sub02_run_busy;
	wire signed [12:0] w_sub02_u_addr;
	reg  signed [12:0] r_sub02_u_addr;
	wire        [31:0] w_sub02_u_datain;
	reg         [31:0] r_sub02_u_datain;
	wire        [31:0] w_sub02_u_dataout;
	wire               w_sub02_u_r_w;
	reg                r_sub02_u_r_w;
	wire signed [12:0] w_sub02_result_addr;
	reg  signed [12:0] r_sub02_result_addr;
	wire        [31:0] w_sub02_result_datain;
	reg         [31:0] r_sub02_result_datain;
	wire        [31:0] w_sub02_result_dataout;
	wire               w_sub02_result_r_w;
	reg                r_sub02_result_r_w;
	reg                r_sub11_run_req;
	wire               w_sub11_run_busy;
	wire signed [12:0] w_sub11_u_addr;
	reg  signed [12:0] r_sub11_u_addr;
	wire        [31:0] w_sub11_u_datain;
	reg         [31:0] r_sub11_u_datain;
	wire        [31:0] w_sub11_u_dataout;
	wire               w_sub11_u_r_w;
	reg                r_sub11_u_r_w;
	wire signed [12:0] w_sub11_result_addr;
	reg  signed [12:0] r_sub11_result_addr;
	wire        [31:0] w_sub11_result_datain;
	reg         [31:0] r_sub11_result_datain;
	wire        [31:0] w_sub11_result_dataout;
	wire               w_sub11_result_r_w;
	reg                r_sub11_result_r_w;
	reg                r_sub14_run_req;
	wire               w_sub14_run_busy;
	wire signed [12:0] w_sub14_u_addr;
	reg  signed [12:0] r_sub14_u_addr;
	wire        [31:0] w_sub14_u_datain;
	reg         [31:0] r_sub14_u_datain;
	wire        [31:0] w_sub14_u_dataout;
	wire               w_sub14_u_r_w;
	reg                r_sub14_u_r_w;
	wire signed [12:0] w_sub14_result_addr;
	reg  signed [12:0] r_sub14_result_addr;
	wire        [31:0] w_sub14_result_datain;
	reg         [31:0] r_sub14_result_datain;
	wire        [31:0] w_sub14_result_dataout;
	wire               w_sub14_result_r_w;
	reg                r_sub14_result_r_w;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [12:0] w_sub01_u_addr;
	reg  signed [12:0] r_sub01_u_addr;
	wire        [31:0] w_sub01_u_datain;
	reg         [31:0] r_sub01_u_datain;
	wire        [31:0] w_sub01_u_dataout;
	wire               w_sub01_u_r_w;
	reg                r_sub01_u_r_w;
	wire signed [12:0] w_sub01_result_addr;
	reg  signed [12:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub13_run_req;
	wire               w_sub13_run_busy;
	wire signed [12:0] w_sub13_u_addr;
	reg  signed [12:0] r_sub13_u_addr;
	wire        [31:0] w_sub13_u_datain;
	reg         [31:0] r_sub13_u_datain;
	wire        [31:0] w_sub13_u_dataout;
	wire               w_sub13_u_r_w;
	reg                r_sub13_u_r_w;
	wire signed [12:0] w_sub13_result_addr;
	reg  signed [12:0] r_sub13_result_addr;
	wire        [31:0] w_sub13_result_datain;
	reg         [31:0] r_sub13_result_datain;
	wire        [31:0] w_sub13_result_dataout;
	wire               w_sub13_result_r_w;
	reg                r_sub13_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [12:0] w_sub00_u_addr;
	reg  signed [12:0] r_sub00_u_addr;
	wire        [31:0] w_sub00_u_datain;
	reg         [31:0] r_sub00_u_datain;
	wire        [31:0] w_sub00_u_dataout;
	wire               w_sub00_u_r_w;
	reg                r_sub00_u_r_w;
	wire signed [12:0] w_sub00_result_addr;
	reg  signed [12:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	reg                r_sub07_run_req;
	wire               w_sub07_run_busy;
	wire signed [12:0] w_sub07_u_addr;
	reg  signed [12:0] r_sub07_u_addr;
	wire        [31:0] w_sub07_u_datain;
	reg         [31:0] r_sub07_u_datain;
	wire        [31:0] w_sub07_u_dataout;
	wire               w_sub07_u_r_w;
	reg                r_sub07_u_r_w;
	wire signed [12:0] w_sub07_result_addr;
	reg  signed [12:0] r_sub07_result_addr;
	wire        [31:0] w_sub07_result_datain;
	reg         [31:0] r_sub07_result_datain;
	wire        [31:0] w_sub07_result_dataout;
	wire               w_sub07_result_r_w;
	reg                r_sub07_result_r_w;
	reg                r_sub06_run_req;
	wire               w_sub06_run_busy;
	wire signed [12:0] w_sub06_u_addr;
	reg  signed [12:0] r_sub06_u_addr;
	wire        [31:0] w_sub06_u_datain;
	reg         [31:0] r_sub06_u_datain;
	wire        [31:0] w_sub06_u_dataout;
	wire               w_sub06_u_r_w;
	reg                r_sub06_u_r_w;
	wire signed [12:0] w_sub06_result_addr;
	reg  signed [12:0] r_sub06_result_addr;
	wire        [31:0] w_sub06_result_datain;
	reg         [31:0] r_sub06_result_datain;
	wire        [31:0] w_sub06_result_dataout;
	wire               w_sub06_result_r_w;
	reg                r_sub06_result_r_w;
	reg                r_sub15_run_req;
	wire               w_sub15_run_busy;
	wire signed [12:0] w_sub15_u_addr;
	reg  signed [12:0] r_sub15_u_addr;
	wire        [31:0] w_sub15_u_datain;
	reg         [31:0] r_sub15_u_datain;
	wire        [31:0] w_sub15_u_dataout;
	wire               w_sub15_u_r_w;
	reg                r_sub15_u_r_w;
	wire signed [12:0] w_sub15_result_addr;
	reg  signed [12:0] r_sub15_result_addr;
	wire        [31:0] w_sub15_result_datain;
	reg         [31:0] r_sub15_result_datain;
	wire        [31:0] w_sub15_result_dataout;
	wire               w_sub15_result_r_w;
	reg                r_sub15_result_r_w;
	reg                r_sub05_run_req;
	wire               w_sub05_run_busy;
	wire signed [12:0] w_sub05_u_addr;
	reg  signed [12:0] r_sub05_u_addr;
	wire        [31:0] w_sub05_u_datain;
	reg         [31:0] r_sub05_u_datain;
	wire        [31:0] w_sub05_u_dataout;
	wire               w_sub05_u_r_w;
	reg                r_sub05_u_r_w;
	wire signed [12:0] w_sub05_result_addr;
	reg  signed [12:0] r_sub05_result_addr;
	wire        [31:0] w_sub05_result_datain;
	reg         [31:0] r_sub05_result_datain;
	wire        [31:0] w_sub05_result_dataout;
	wire               w_sub05_result_r_w;
	reg                r_sub05_result_r_w;
	reg                r_sub04_run_req;
	wire               w_sub04_run_busy;
	wire signed [12:0] w_sub04_u_addr;
	reg  signed [12:0] r_sub04_u_addr;
	wire        [31:0] w_sub04_u_datain;
	reg         [31:0] r_sub04_u_datain;
	wire        [31:0] w_sub04_u_dataout;
	wire               w_sub04_u_r_w;
	reg                r_sub04_u_r_w;
	wire signed [12:0] w_sub04_result_addr;
	reg  signed [12:0] r_sub04_result_addr;
	wire        [31:0] w_sub04_result_datain;
	reg         [31:0] r_sub04_result_datain;
	wire        [31:0] w_sub04_result_dataout;
	wire               w_sub04_result_r_w;
	reg                r_sub04_result_r_w;
	reg                r_sub10_run_req;
	wire               w_sub10_run_busy;
	wire signed [12:0] w_sub10_u_addr;
	reg  signed [12:0] r_sub10_u_addr;
	wire        [31:0] w_sub10_u_datain;
	reg         [31:0] r_sub10_u_datain;
	wire        [31:0] w_sub10_u_dataout;
	wire               w_sub10_u_r_w;
	reg                r_sub10_u_r_w;
	wire signed [12:0] w_sub10_result_addr;
	reg  signed [12:0] r_sub10_result_addr;
	wire        [31:0] w_sub10_result_datain;
	reg         [31:0] r_sub10_result_datain;
	wire        [31:0] w_sub10_result_dataout;
	wire               w_sub10_result_r_w;
	reg                r_sub10_result_r_w;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	wire signed [31:0] w_sys_tmp1;
	wire signed [31:0] w_sys_tmp3;
	wire               w_sys_tmp4;
	wire               w_sys_tmp5;
	wire signed [31:0] w_sys_tmp6;
	wire               w_sys_tmp7;
	wire               w_sys_tmp8;
	wire signed [31:0] w_sys_tmp11;
	wire signed [31:0] w_sys_tmp12;
	wire signed [31:0] w_sys_tmp13;
	wire        [31:0] w_sys_tmp14;
	wire signed [31:0] w_sys_tmp15;
	wire               w_sys_tmp52;
	wire               w_sys_tmp53;
	wire signed [31:0] w_sys_tmp54;
	wire signed [31:0] w_sys_tmp55;
	wire               w_sys_tmp56;
	wire               w_sys_tmp57;
	wire signed [31:0] w_sys_tmp58;
	wire signed [31:0] w_sys_tmp61;
	wire signed [31:0] w_sys_tmp62;
	wire signed [31:0] w_sys_tmp63;
	wire        [31:0] w_sys_tmp64;
	wire signed [31:0] w_sys_tmp65;
	wire signed [31:0] w_sys_tmp66;
	wire signed [31:0] w_sys_tmp68;
	wire signed [31:0] w_sys_tmp69;
	wire signed [31:0] w_sys_tmp130;
	wire               w_sys_tmp131;
	wire               w_sys_tmp132;
	wire signed [31:0] w_sys_tmp133;
	wire signed [31:0] w_sys_tmp136;
	wire signed [31:0] w_sys_tmp137;
	wire signed [31:0] w_sys_tmp138;
	wire        [31:0] w_sys_tmp139;
	wire signed [31:0] w_sys_tmp140;
	wire signed [31:0] w_sys_tmp141;
	wire signed [31:0] w_sys_tmp142;
	wire signed [31:0] w_sys_tmp143;
	wire signed [31:0] w_sys_tmp144;
	wire signed [31:0] w_sys_tmp205;
	wire               w_sys_tmp206;
	wire               w_sys_tmp207;
	wire signed [31:0] w_sys_tmp208;
	wire signed [31:0] w_sys_tmp211;
	wire signed [31:0] w_sys_tmp212;
	wire signed [31:0] w_sys_tmp213;
	wire        [31:0] w_sys_tmp214;
	wire signed [31:0] w_sys_tmp215;
	wire signed [31:0] w_sys_tmp216;
	wire signed [31:0] w_sys_tmp218;
	wire signed [31:0] w_sys_tmp219;
	wire signed [31:0] w_sys_tmp280;
	wire               w_sys_tmp281;
	wire               w_sys_tmp282;
	wire signed [31:0] w_sys_tmp283;
	wire signed [31:0] w_sys_tmp286;
	wire signed [31:0] w_sys_tmp287;
	wire signed [31:0] w_sys_tmp288;
	wire        [31:0] w_sys_tmp289;
	wire signed [31:0] w_sys_tmp290;
	wire signed [31:0] w_sys_tmp291;
	wire signed [31:0] w_sys_tmp293;
	wire signed [31:0] w_sys_tmp294;
	wire signed [31:0] w_sys_tmp355;
	wire               w_sys_tmp356;
	wire               w_sys_tmp357;
	wire signed [31:0] w_sys_tmp358;
	wire signed [31:0] w_sys_tmp359;
	wire               w_sys_tmp360;
	wire               w_sys_tmp361;
	wire signed [31:0] w_sys_tmp362;
	wire signed [31:0] w_sys_tmp365;
	wire signed [31:0] w_sys_tmp366;
	wire signed [31:0] w_sys_tmp367;
	wire        [31:0] w_sys_tmp368;
	wire signed [31:0] w_sys_tmp369;
	wire signed [31:0] w_sys_tmp370;
	wire signed [31:0] w_sys_tmp372;
	wire signed [31:0] w_sys_tmp373;
	wire signed [31:0] w_sys_tmp434;
	wire               w_sys_tmp435;
	wire               w_sys_tmp436;
	wire signed [31:0] w_sys_tmp437;
	wire signed [31:0] w_sys_tmp440;
	wire signed [31:0] w_sys_tmp441;
	wire signed [31:0] w_sys_tmp442;
	wire        [31:0] w_sys_tmp443;
	wire signed [31:0] w_sys_tmp444;
	wire signed [31:0] w_sys_tmp445;
	wire signed [31:0] w_sys_tmp447;
	wire signed [31:0] w_sys_tmp448;
	wire signed [31:0] w_sys_tmp509;
	wire               w_sys_tmp510;
	wire               w_sys_tmp511;
	wire signed [31:0] w_sys_tmp512;
	wire signed [31:0] w_sys_tmp515;
	wire signed [31:0] w_sys_tmp516;
	wire signed [31:0] w_sys_tmp517;
	wire        [31:0] w_sys_tmp518;
	wire signed [31:0] w_sys_tmp519;
	wire signed [31:0] w_sys_tmp520;
	wire signed [31:0] w_sys_tmp522;
	wire signed [31:0] w_sys_tmp523;
	wire signed [31:0] w_sys_tmp584;
	wire               w_sys_tmp585;
	wire               w_sys_tmp586;
	wire signed [31:0] w_sys_tmp587;
	wire signed [31:0] w_sys_tmp590;
	wire signed [31:0] w_sys_tmp591;
	wire signed [31:0] w_sys_tmp592;
	wire        [31:0] w_sys_tmp593;
	wire signed [31:0] w_sys_tmp594;
	wire signed [31:0] w_sys_tmp595;
	wire signed [31:0] w_sys_tmp597;
	wire signed [31:0] w_sys_tmp598;
	wire signed [31:0] w_sys_tmp659;
	wire               w_sys_tmp660;
	wire               w_sys_tmp661;
	wire signed [31:0] w_sys_tmp662;
	wire signed [31:0] w_sys_tmp663;
	wire               w_sys_tmp664;
	wire               w_sys_tmp665;
	wire signed [31:0] w_sys_tmp666;
	wire signed [31:0] w_sys_tmp669;
	wire signed [31:0] w_sys_tmp670;
	wire signed [31:0] w_sys_tmp671;
	wire        [31:0] w_sys_tmp672;
	wire signed [31:0] w_sys_tmp673;
	wire signed [31:0] w_sys_tmp674;
	wire signed [31:0] w_sys_tmp676;
	wire signed [31:0] w_sys_tmp677;
	wire signed [31:0] w_sys_tmp738;
	wire               w_sys_tmp739;
	wire               w_sys_tmp740;
	wire signed [31:0] w_sys_tmp741;
	wire signed [31:0] w_sys_tmp744;
	wire signed [31:0] w_sys_tmp745;
	wire signed [31:0] w_sys_tmp746;
	wire        [31:0] w_sys_tmp747;
	wire signed [31:0] w_sys_tmp748;
	wire signed [31:0] w_sys_tmp749;
	wire signed [31:0] w_sys_tmp751;
	wire signed [31:0] w_sys_tmp752;
	wire signed [31:0] w_sys_tmp813;
	wire               w_sys_tmp814;
	wire               w_sys_tmp815;
	wire signed [31:0] w_sys_tmp816;
	wire signed [31:0] w_sys_tmp819;
	wire signed [31:0] w_sys_tmp820;
	wire signed [31:0] w_sys_tmp821;
	wire        [31:0] w_sys_tmp822;
	wire signed [31:0] w_sys_tmp823;
	wire signed [31:0] w_sys_tmp824;
	wire signed [31:0] w_sys_tmp826;
	wire signed [31:0] w_sys_tmp827;
	wire signed [31:0] w_sys_tmp888;
	wire               w_sys_tmp889;
	wire               w_sys_tmp890;
	wire signed [31:0] w_sys_tmp891;
	wire signed [31:0] w_sys_tmp894;
	wire signed [31:0] w_sys_tmp895;
	wire signed [31:0] w_sys_tmp896;
	wire        [31:0] w_sys_tmp897;
	wire signed [31:0] w_sys_tmp898;
	wire signed [31:0] w_sys_tmp899;
	wire signed [31:0] w_sys_tmp901;
	wire signed [31:0] w_sys_tmp902;
	wire signed [31:0] w_sys_tmp963;
	wire               w_sys_tmp964;
	wire               w_sys_tmp965;
	wire signed [31:0] w_sys_tmp966;
	wire signed [31:0] w_sys_tmp967;
	wire               w_sys_tmp968;
	wire               w_sys_tmp969;
	wire signed [31:0] w_sys_tmp970;
	wire signed [31:0] w_sys_tmp973;
	wire signed [31:0] w_sys_tmp974;
	wire signed [31:0] w_sys_tmp975;
	wire        [31:0] w_sys_tmp976;
	wire signed [31:0] w_sys_tmp977;
	wire signed [31:0] w_sys_tmp978;
	wire signed [31:0] w_sys_tmp980;
	wire signed [31:0] w_sys_tmp981;
	wire signed [31:0] w_sys_tmp1042;
	wire               w_sys_tmp1043;
	wire               w_sys_tmp1044;
	wire signed [31:0] w_sys_tmp1045;
	wire signed [31:0] w_sys_tmp1048;
	wire signed [31:0] w_sys_tmp1049;
	wire signed [31:0] w_sys_tmp1050;
	wire        [31:0] w_sys_tmp1051;
	wire signed [31:0] w_sys_tmp1052;
	wire signed [31:0] w_sys_tmp1053;
	wire signed [31:0] w_sys_tmp1055;
	wire signed [31:0] w_sys_tmp1056;
	wire signed [31:0] w_sys_tmp1117;
	wire               w_sys_tmp1118;
	wire               w_sys_tmp1119;
	wire signed [31:0] w_sys_tmp1120;
	wire signed [31:0] w_sys_tmp1123;
	wire signed [31:0] w_sys_tmp1124;
	wire signed [31:0] w_sys_tmp1125;
	wire        [31:0] w_sys_tmp1126;
	wire signed [31:0] w_sys_tmp1127;
	wire signed [31:0] w_sys_tmp1128;
	wire signed [31:0] w_sys_tmp1130;
	wire signed [31:0] w_sys_tmp1131;
	wire signed [31:0] w_sys_tmp1192;
	wire               w_sys_tmp1193;
	wire               w_sys_tmp1194;
	wire signed [31:0] w_sys_tmp1195;
	wire signed [31:0] w_sys_tmp1198;
	wire signed [31:0] w_sys_tmp1199;
	wire signed [31:0] w_sys_tmp1200;
	wire        [31:0] w_sys_tmp1201;
	wire signed [31:0] w_sys_tmp1202;
	wire signed [31:0] w_sys_tmp1203;
	wire signed [31:0] w_sys_tmp1205;
	wire signed [31:0] w_sys_tmp1206;
	wire               w_sys_tmp1267;
	wire               w_sys_tmp1268;
	wire signed [31:0] w_sys_tmp1269;
	wire signed [31:0] w_sys_tmp1270;
	wire               w_sys_tmp1271;
	wire               w_sys_tmp1272;
	wire signed [31:0] w_sys_tmp1273;
	wire signed [31:0] w_sys_tmp1276;
	wire signed [31:0] w_sys_tmp1277;
	wire        [31:0] w_sys_tmp1278;
	wire signed [31:0] w_sys_tmp1282;
	wire signed [31:0] w_sys_tmp1283;
	wire        [31:0] w_sys_tmp1284;
	wire signed [31:0] w_sys_tmp1288;
	wire signed [31:0] w_sys_tmp1289;
	wire signed [31:0] w_sys_tmp1293;
	wire signed [31:0] w_sys_tmp1294;
	wire signed [31:0] w_sys_tmp1299;
	wire signed [31:0] w_sys_tmp1300;
	wire signed [31:0] w_sys_tmp1304;
	wire signed [31:0] w_sys_tmp1305;
	wire        [31:0] w_sys_tmp1306;
	wire signed [31:0] w_sys_tmp1309;
	wire signed [31:0] w_sys_tmp1310;
	wire               w_sys_tmp1311;
	wire               w_sys_tmp1312;
	wire signed [31:0] w_sys_tmp1313;
	wire signed [31:0] w_sys_tmp1316;
	wire signed [31:0] w_sys_tmp1317;
	wire        [31:0] w_sys_tmp1318;
	wire signed [31:0] w_sys_tmp1322;
	wire signed [31:0] w_sys_tmp1323;
	wire        [31:0] w_sys_tmp1324;
	wire signed [31:0] w_sys_tmp1328;
	wire signed [31:0] w_sys_tmp1329;
	wire signed [31:0] w_sys_tmp1333;
	wire signed [31:0] w_sys_tmp1334;
	wire signed [31:0] w_sys_tmp1339;
	wire signed [31:0] w_sys_tmp1340;
	wire signed [31:0] w_sys_tmp1344;
	wire signed [31:0] w_sys_tmp1345;
	wire        [31:0] w_sys_tmp1346;
	wire signed [31:0] w_sys_tmp1349;
	wire signed [31:0] w_sys_tmp1350;
	wire               w_sys_tmp1351;
	wire               w_sys_tmp1352;
	wire signed [31:0] w_sys_tmp1353;
	wire signed [31:0] w_sys_tmp1356;
	wire signed [31:0] w_sys_tmp1357;
	wire        [31:0] w_sys_tmp1358;
	wire signed [31:0] w_sys_tmp1362;
	wire signed [31:0] w_sys_tmp1363;
	wire        [31:0] w_sys_tmp1364;
	wire signed [31:0] w_sys_tmp1368;
	wire signed [31:0] w_sys_tmp1369;
	wire signed [31:0] w_sys_tmp1373;
	wire signed [31:0] w_sys_tmp1374;
	wire signed [31:0] w_sys_tmp1379;
	wire signed [31:0] w_sys_tmp1380;
	wire signed [31:0] w_sys_tmp1384;
	wire signed [31:0] w_sys_tmp1385;
	wire        [31:0] w_sys_tmp1386;
	wire signed [31:0] w_sys_tmp1389;
	wire signed [31:0] w_sys_tmp1390;
	wire               w_sys_tmp1391;
	wire               w_sys_tmp1392;
	wire signed [31:0] w_sys_tmp1393;
	wire signed [31:0] w_sys_tmp1396;
	wire signed [31:0] w_sys_tmp1397;
	wire        [31:0] w_sys_tmp1398;
	wire signed [31:0] w_sys_tmp1402;
	wire signed [31:0] w_sys_tmp1403;
	wire        [31:0] w_sys_tmp1404;
	wire signed [31:0] w_sys_tmp1408;
	wire signed [31:0] w_sys_tmp1409;
	wire signed [31:0] w_sys_tmp1413;
	wire signed [31:0] w_sys_tmp1414;
	wire signed [31:0] w_sys_tmp1419;
	wire signed [31:0] w_sys_tmp1420;
	wire signed [31:0] w_sys_tmp1424;
	wire signed [31:0] w_sys_tmp1425;
	wire        [31:0] w_sys_tmp1426;
	wire signed [31:0] w_sys_tmp1429;
	wire signed [31:0] w_sys_tmp1430;
	wire               w_sys_tmp1431;
	wire               w_sys_tmp1432;
	wire signed [31:0] w_sys_tmp1433;
	wire signed [31:0] w_sys_tmp1436;
	wire signed [31:0] w_sys_tmp1437;
	wire signed [31:0] w_sys_tmp1438;
	wire signed [31:0] w_sys_tmp1439;
	wire        [31:0] w_sys_tmp1440;
	wire signed [31:0] w_sys_tmp1441;
	wire signed [31:0] w_sys_tmp1442;
	wire signed [31:0] w_sys_tmp1446;
	wire signed [31:0] w_sys_tmp1447;
	wire signed [31:0] w_sys_tmp1449;
	wire        [31:0] w_sys_tmp1450;
	wire signed [31:0] w_sys_tmp1451;
	wire signed [31:0] w_sys_tmp1452;
	wire signed [31:0] w_sys_tmp1456;
	wire signed [31:0] w_sys_tmp1457;
	wire signed [31:0] w_sys_tmp1459;
	wire signed [31:0] w_sys_tmp1460;
	wire signed [31:0] w_sys_tmp1461;
	wire signed [31:0] w_sys_tmp1465;
	wire signed [31:0] w_sys_tmp1466;
	wire signed [31:0] w_sys_tmp1468;
	wire signed [31:0] w_sys_tmp1470;
	wire signed [31:0] w_sys_tmp1471;
	wire signed [31:0] w_sys_tmp1475;
	wire signed [31:0] w_sys_tmp1476;
	wire signed [31:0] w_sys_tmp1478;
	wire signed [31:0] w_sys_tmp1479;
	wire signed [31:0] w_sys_tmp1480;
	wire signed [31:0] w_sys_tmp1484;
	wire signed [31:0] w_sys_tmp1485;
	wire signed [31:0] w_sys_tmp1487;
	wire        [31:0] w_sys_tmp1488;
	wire signed [31:0] w_sys_tmp1489;
	wire signed [31:0] w_sys_tmp1490;
	wire signed [31:0] w_sys_tmp1493;
	wire signed [31:0] w_sys_tmp1494;
	wire signed [31:0] w_sys_tmp1495;
	wire signed [31:0] w_sys_tmp1496;
	wire signed [31:0] w_sys_tmp1497;
	wire signed [31:0] w_sys_tmp1498;
	wire signed [31:0] w_sys_tmp1499;
	wire signed [31:0] w_sys_tmp1500;
	wire signed [31:0] w_sys_tmp1501;
	wire signed [31:0] w_sys_tmp1502;
	wire signed [31:0] w_sys_tmp1503;
	wire signed [31:0] w_sys_tmp1504;
	wire signed [31:0] w_sys_tmp1931;
	wire               w_sys_tmp1932;
	wire               w_sys_tmp1933;
	wire signed [31:0] w_sys_tmp1934;
	wire signed [31:0] w_sys_tmp1937;
	wire signed [31:0] w_sys_tmp1938;
	wire signed [31:0] w_sys_tmp1939;
	wire signed [31:0] w_sys_tmp1940;
	wire        [31:0] w_sys_tmp1941;
	wire signed [31:0] w_sys_tmp1942;
	wire signed [31:0] w_sys_tmp1943;
	wire signed [31:0] w_sys_tmp1947;
	wire signed [31:0] w_sys_tmp1948;
	wire signed [31:0] w_sys_tmp1950;
	wire        [31:0] w_sys_tmp1951;
	wire signed [31:0] w_sys_tmp1952;
	wire signed [31:0] w_sys_tmp1953;
	wire signed [31:0] w_sys_tmp1957;
	wire signed [31:0] w_sys_tmp1958;
	wire signed [31:0] w_sys_tmp1960;
	wire signed [31:0] w_sys_tmp1961;
	wire signed [31:0] w_sys_tmp1962;
	wire signed [31:0] w_sys_tmp1966;
	wire signed [31:0] w_sys_tmp1967;
	wire signed [31:0] w_sys_tmp1969;
	wire signed [31:0] w_sys_tmp1971;
	wire signed [31:0] w_sys_tmp1972;
	wire signed [31:0] w_sys_tmp1976;
	wire signed [31:0] w_sys_tmp1977;
	wire signed [31:0] w_sys_tmp1979;
	wire signed [31:0] w_sys_tmp1980;
	wire signed [31:0] w_sys_tmp1981;
	wire signed [31:0] w_sys_tmp1985;
	wire signed [31:0] w_sys_tmp1986;
	wire signed [31:0] w_sys_tmp1988;
	wire        [31:0] w_sys_tmp1989;
	wire signed [31:0] w_sys_tmp1990;
	wire signed [31:0] w_sys_tmp1991;
	wire signed [31:0] w_sys_tmp1994;
	wire signed [31:0] w_sys_tmp1995;
	wire signed [31:0] w_sys_tmp1996;
	wire signed [31:0] w_sys_tmp1997;
	wire signed [31:0] w_sys_tmp1998;
	wire signed [31:0] w_sys_tmp1999;
	wire signed [31:0] w_sys_tmp2000;
	wire signed [31:0] w_sys_tmp2001;
	wire signed [31:0] w_sys_tmp2002;
	wire signed [31:0] w_sys_tmp2003;
	wire signed [31:0] w_sys_tmp2004;
	wire signed [31:0] w_sys_tmp2005;
	wire signed [31:0] w_sys_tmp2432;
	wire               w_sys_tmp2433;
	wire               w_sys_tmp2434;
	wire signed [31:0] w_sys_tmp2435;
	wire signed [31:0] w_sys_tmp2438;
	wire signed [31:0] w_sys_tmp2439;
	wire signed [31:0] w_sys_tmp2440;
	wire signed [31:0] w_sys_tmp2441;
	wire        [31:0] w_sys_tmp2442;
	wire signed [31:0] w_sys_tmp2443;
	wire signed [31:0] w_sys_tmp2444;
	wire signed [31:0] w_sys_tmp2448;
	wire signed [31:0] w_sys_tmp2449;
	wire signed [31:0] w_sys_tmp2451;
	wire        [31:0] w_sys_tmp2452;
	wire signed [31:0] w_sys_tmp2453;
	wire signed [31:0] w_sys_tmp2454;
	wire signed [31:0] w_sys_tmp2458;
	wire signed [31:0] w_sys_tmp2459;
	wire signed [31:0] w_sys_tmp2461;
	wire signed [31:0] w_sys_tmp2462;
	wire signed [31:0] w_sys_tmp2463;
	wire signed [31:0] w_sys_tmp2467;
	wire signed [31:0] w_sys_tmp2468;
	wire signed [31:0] w_sys_tmp2470;
	wire signed [31:0] w_sys_tmp2472;
	wire signed [31:0] w_sys_tmp2473;
	wire signed [31:0] w_sys_tmp2477;
	wire signed [31:0] w_sys_tmp2478;
	wire signed [31:0] w_sys_tmp2480;
	wire signed [31:0] w_sys_tmp2481;
	wire signed [31:0] w_sys_tmp2482;
	wire signed [31:0] w_sys_tmp2486;
	wire signed [31:0] w_sys_tmp2487;
	wire signed [31:0] w_sys_tmp2489;
	wire        [31:0] w_sys_tmp2490;
	wire signed [31:0] w_sys_tmp2491;
	wire signed [31:0] w_sys_tmp2492;
	wire signed [31:0] w_sys_tmp2495;
	wire signed [31:0] w_sys_tmp2496;
	wire signed [31:0] w_sys_tmp2497;
	wire signed [31:0] w_sys_tmp2498;
	wire signed [31:0] w_sys_tmp2499;
	wire signed [31:0] w_sys_tmp2500;
	wire signed [31:0] w_sys_tmp2501;
	wire signed [31:0] w_sys_tmp2502;
	wire signed [31:0] w_sys_tmp2503;
	wire signed [31:0] w_sys_tmp2504;
	wire signed [31:0] w_sys_tmp2505;
	wire signed [31:0] w_sys_tmp2506;
	wire signed [31:0] w_sys_tmp2933;
	wire               w_sys_tmp2934;
	wire               w_sys_tmp2935;
	wire signed [31:0] w_sys_tmp2936;
	wire signed [31:0] w_sys_tmp2939;
	wire signed [31:0] w_sys_tmp2940;
	wire signed [31:0] w_sys_tmp2941;
	wire signed [31:0] w_sys_tmp2942;
	wire        [31:0] w_sys_tmp2943;
	wire signed [31:0] w_sys_tmp2944;
	wire signed [31:0] w_sys_tmp2945;
	wire signed [31:0] w_sys_tmp2949;
	wire signed [31:0] w_sys_tmp2950;
	wire signed [31:0] w_sys_tmp2952;
	wire        [31:0] w_sys_tmp2953;
	wire signed [31:0] w_sys_tmp2954;
	wire signed [31:0] w_sys_tmp2955;
	wire signed [31:0] w_sys_tmp2959;
	wire signed [31:0] w_sys_tmp2960;
	wire signed [31:0] w_sys_tmp2962;
	wire signed [31:0] w_sys_tmp2963;
	wire signed [31:0] w_sys_tmp2964;
	wire signed [31:0] w_sys_tmp2968;
	wire signed [31:0] w_sys_tmp2969;
	wire signed [31:0] w_sys_tmp2971;
	wire signed [31:0] w_sys_tmp2973;
	wire signed [31:0] w_sys_tmp2974;
	wire signed [31:0] w_sys_tmp2978;
	wire signed [31:0] w_sys_tmp2979;
	wire signed [31:0] w_sys_tmp2981;
	wire signed [31:0] w_sys_tmp2982;
	wire signed [31:0] w_sys_tmp2983;
	wire signed [31:0] w_sys_tmp2987;
	wire signed [31:0] w_sys_tmp2988;
	wire signed [31:0] w_sys_tmp2990;
	wire        [31:0] w_sys_tmp2991;
	wire signed [31:0] w_sys_tmp2992;
	wire signed [31:0] w_sys_tmp2993;
	wire signed [31:0] w_sys_tmp2996;
	wire signed [31:0] w_sys_tmp2997;
	wire signed [31:0] w_sys_tmp2998;
	wire signed [31:0] w_sys_tmp2999;
	wire signed [31:0] w_sys_tmp3000;
	wire signed [31:0] w_sys_tmp3001;
	wire signed [31:0] w_sys_tmp3002;
	wire signed [31:0] w_sys_tmp3003;
	wire signed [31:0] w_sys_tmp3004;
	wire signed [31:0] w_sys_tmp3005;
	wire signed [31:0] w_sys_tmp3006;
	wire signed [31:0] w_sys_tmp3007;
	wire signed [31:0] w_sys_tmp3434;
	wire               w_sys_tmp3435;
	wire               w_sys_tmp3436;
	wire signed [31:0] w_sys_tmp3437;
	wire signed [31:0] w_sys_tmp3438;
	wire signed [31:0] w_sys_tmp3439;
	wire               w_sys_tmp3440;
	wire               w_sys_tmp3441;
	wire signed [31:0] w_sys_tmp3442;
	wire signed [31:0] w_sys_tmp3445;
	wire signed [31:0] w_sys_tmp3446;
	wire signed [31:0] w_sys_tmp3447;
	wire        [31:0] w_sys_tmp3448;
	wire signed [31:0] w_sys_tmp3449;
	wire signed [31:0] w_sys_tmp3450;
	wire signed [31:0] w_sys_tmp3452;
	wire signed [31:0] w_sys_tmp3453;
	wire signed [31:0] w_sys_tmp3514;
	wire               w_sys_tmp3515;
	wire               w_sys_tmp3516;
	wire signed [31:0] w_sys_tmp3517;
	wire signed [31:0] w_sys_tmp3520;
	wire signed [31:0] w_sys_tmp3521;
	wire signed [31:0] w_sys_tmp3522;
	wire        [31:0] w_sys_tmp3523;
	wire signed [31:0] w_sys_tmp3524;
	wire signed [31:0] w_sys_tmp3525;
	wire signed [31:0] w_sys_tmp3527;
	wire signed [31:0] w_sys_tmp3528;
	wire signed [31:0] w_sys_tmp3589;
	wire               w_sys_tmp3590;
	wire               w_sys_tmp3591;
	wire signed [31:0] w_sys_tmp3592;
	wire signed [31:0] w_sys_tmp3595;
	wire signed [31:0] w_sys_tmp3596;
	wire signed [31:0] w_sys_tmp3597;
	wire        [31:0] w_sys_tmp3598;
	wire signed [31:0] w_sys_tmp3599;
	wire signed [31:0] w_sys_tmp3600;
	wire signed [31:0] w_sys_tmp3602;
	wire signed [31:0] w_sys_tmp3603;
	wire signed [31:0] w_sys_tmp3664;
	wire               w_sys_tmp3665;
	wire               w_sys_tmp3666;
	wire signed [31:0] w_sys_tmp3667;
	wire signed [31:0] w_sys_tmp3670;
	wire signed [31:0] w_sys_tmp3671;
	wire signed [31:0] w_sys_tmp3672;
	wire        [31:0] w_sys_tmp3673;
	wire signed [31:0] w_sys_tmp3674;
	wire signed [31:0] w_sys_tmp3675;
	wire signed [31:0] w_sys_tmp3677;
	wire signed [31:0] w_sys_tmp3678;
	wire signed [31:0] w_sys_tmp3739;
	wire               w_sys_tmp3740;
	wire               w_sys_tmp3741;
	wire signed [31:0] w_sys_tmp3742;
	wire signed [31:0] w_sys_tmp3743;
	wire signed [31:0] w_sys_tmp3744;
	wire               w_sys_tmp3745;
	wire               w_sys_tmp3746;
	wire signed [31:0] w_sys_tmp3747;
	wire signed [31:0] w_sys_tmp3750;
	wire signed [31:0] w_sys_tmp3751;
	wire signed [31:0] w_sys_tmp3752;
	wire        [31:0] w_sys_tmp3753;
	wire signed [31:0] w_sys_tmp3754;
	wire signed [31:0] w_sys_tmp3755;
	wire signed [31:0] w_sys_tmp3757;
	wire signed [31:0] w_sys_tmp3758;
	wire signed [31:0] w_sys_tmp3819;
	wire               w_sys_tmp3820;
	wire               w_sys_tmp3821;
	wire signed [31:0] w_sys_tmp3822;
	wire signed [31:0] w_sys_tmp3825;
	wire signed [31:0] w_sys_tmp3826;
	wire signed [31:0] w_sys_tmp3827;
	wire        [31:0] w_sys_tmp3828;
	wire signed [31:0] w_sys_tmp3829;
	wire signed [31:0] w_sys_tmp3830;
	wire signed [31:0] w_sys_tmp3832;
	wire signed [31:0] w_sys_tmp3833;
	wire signed [31:0] w_sys_tmp3894;
	wire               w_sys_tmp3895;
	wire               w_sys_tmp3896;
	wire signed [31:0] w_sys_tmp3897;
	wire signed [31:0] w_sys_tmp3900;
	wire signed [31:0] w_sys_tmp3901;
	wire signed [31:0] w_sys_tmp3902;
	wire        [31:0] w_sys_tmp3903;
	wire signed [31:0] w_sys_tmp3904;
	wire signed [31:0] w_sys_tmp3905;
	wire signed [31:0] w_sys_tmp3907;
	wire signed [31:0] w_sys_tmp3908;
	wire signed [31:0] w_sys_tmp3969;
	wire               w_sys_tmp3970;
	wire               w_sys_tmp3971;
	wire signed [31:0] w_sys_tmp3972;
	wire signed [31:0] w_sys_tmp3975;
	wire signed [31:0] w_sys_tmp3976;
	wire signed [31:0] w_sys_tmp3977;
	wire        [31:0] w_sys_tmp3978;
	wire signed [31:0] w_sys_tmp3979;
	wire signed [31:0] w_sys_tmp3980;
	wire signed [31:0] w_sys_tmp3982;
	wire signed [31:0] w_sys_tmp3983;
	wire signed [31:0] w_sys_tmp4044;
	wire               w_sys_tmp4045;
	wire               w_sys_tmp4046;
	wire signed [31:0] w_sys_tmp4047;
	wire signed [31:0] w_sys_tmp4048;
	wire signed [31:0] w_sys_tmp4049;
	wire               w_sys_tmp4050;
	wire               w_sys_tmp4051;
	wire signed [31:0] w_sys_tmp4052;
	wire signed [31:0] w_sys_tmp4055;
	wire signed [31:0] w_sys_tmp4056;
	wire signed [31:0] w_sys_tmp4057;
	wire        [31:0] w_sys_tmp4058;
	wire signed [31:0] w_sys_tmp4059;
	wire signed [31:0] w_sys_tmp4060;
	wire signed [31:0] w_sys_tmp4062;
	wire signed [31:0] w_sys_tmp4063;
	wire signed [31:0] w_sys_tmp4124;
	wire               w_sys_tmp4125;
	wire               w_sys_tmp4126;
	wire signed [31:0] w_sys_tmp4127;
	wire signed [31:0] w_sys_tmp4130;
	wire signed [31:0] w_sys_tmp4131;
	wire signed [31:0] w_sys_tmp4132;
	wire        [31:0] w_sys_tmp4133;
	wire signed [31:0] w_sys_tmp4134;
	wire signed [31:0] w_sys_tmp4135;
	wire signed [31:0] w_sys_tmp4137;
	wire signed [31:0] w_sys_tmp4138;
	wire signed [31:0] w_sys_tmp4199;
	wire               w_sys_tmp4200;
	wire               w_sys_tmp4201;
	wire signed [31:0] w_sys_tmp4202;
	wire signed [31:0] w_sys_tmp4205;
	wire signed [31:0] w_sys_tmp4206;
	wire signed [31:0] w_sys_tmp4207;
	wire        [31:0] w_sys_tmp4208;
	wire signed [31:0] w_sys_tmp4209;
	wire signed [31:0] w_sys_tmp4210;
	wire signed [31:0] w_sys_tmp4212;
	wire signed [31:0] w_sys_tmp4213;
	wire signed [31:0] w_sys_tmp4274;
	wire               w_sys_tmp4275;
	wire               w_sys_tmp4276;
	wire signed [31:0] w_sys_tmp4277;
	wire signed [31:0] w_sys_tmp4280;
	wire signed [31:0] w_sys_tmp4281;
	wire signed [31:0] w_sys_tmp4282;
	wire        [31:0] w_sys_tmp4283;
	wire signed [31:0] w_sys_tmp4284;
	wire signed [31:0] w_sys_tmp4285;
	wire signed [31:0] w_sys_tmp4287;
	wire signed [31:0] w_sys_tmp4288;
	wire signed [31:0] w_sys_tmp4349;
	wire               w_sys_tmp4350;
	wire               w_sys_tmp4351;
	wire signed [31:0] w_sys_tmp4352;
	wire signed [31:0] w_sys_tmp4353;
	wire signed [31:0] w_sys_tmp4354;
	wire               w_sys_tmp4355;
	wire               w_sys_tmp4356;
	wire signed [31:0] w_sys_tmp4357;
	wire signed [31:0] w_sys_tmp4360;
	wire signed [31:0] w_sys_tmp4361;
	wire signed [31:0] w_sys_tmp4362;
	wire        [31:0] w_sys_tmp4363;
	wire signed [31:0] w_sys_tmp4364;
	wire signed [31:0] w_sys_tmp4365;
	wire signed [31:0] w_sys_tmp4367;
	wire signed [31:0] w_sys_tmp4368;
	wire signed [31:0] w_sys_tmp4429;
	wire               w_sys_tmp4430;
	wire               w_sys_tmp4431;
	wire signed [31:0] w_sys_tmp4432;
	wire signed [31:0] w_sys_tmp4435;
	wire signed [31:0] w_sys_tmp4436;
	wire signed [31:0] w_sys_tmp4437;
	wire        [31:0] w_sys_tmp4438;
	wire signed [31:0] w_sys_tmp4439;
	wire signed [31:0] w_sys_tmp4440;
	wire signed [31:0] w_sys_tmp4442;
	wire signed [31:0] w_sys_tmp4443;
	wire signed [31:0] w_sys_tmp4504;
	wire               w_sys_tmp4505;
	wire               w_sys_tmp4506;
	wire signed [31:0] w_sys_tmp4507;
	wire signed [31:0] w_sys_tmp4510;
	wire signed [31:0] w_sys_tmp4511;
	wire signed [31:0] w_sys_tmp4512;
	wire        [31:0] w_sys_tmp4513;
	wire signed [31:0] w_sys_tmp4514;
	wire signed [31:0] w_sys_tmp4515;
	wire signed [31:0] w_sys_tmp4517;
	wire signed [31:0] w_sys_tmp4518;
	wire signed [31:0] w_sys_tmp4579;
	wire               w_sys_tmp4580;
	wire               w_sys_tmp4581;
	wire signed [31:0] w_sys_tmp4582;
	wire signed [31:0] w_sys_tmp4585;
	wire signed [31:0] w_sys_tmp4586;
	wire signed [31:0] w_sys_tmp4587;
	wire        [31:0] w_sys_tmp4588;
	wire signed [31:0] w_sys_tmp4589;
	wire signed [31:0] w_sys_tmp4590;
	wire signed [31:0] w_sys_tmp4592;
	wire signed [31:0] w_sys_tmp4593;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 5'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 6'h1);
	assign w_fld_u_0_addr_0 = 15'sh0;
	assign w_fld_u_0_datain_0 = 32'h0;
	assign w_fld_u_0_r_w_0 = 1'h0;
	assign w_fld_u_0_ce_0 = w_sys_ce;
	assign w_fld_u_0_ce_1 = w_sys_ce;
	assign w_sub09_u_addr = ( (|r_sys_processing_methodID) ? r_sub09_u_addr : 13'sh0 ) ;
	assign w_sub09_u_datain = ( (|r_sys_processing_methodID) ? r_sub09_u_datain : 32'h0 ) ;
	assign w_sub09_u_r_w = ( (|r_sys_processing_methodID) ? r_sub09_u_r_w : 1'h0 ) ;
	assign w_sub09_result_addr = ( (|r_sys_processing_methodID) ? r_sub09_result_addr : 13'sh0 ) ;
	assign w_sub09_result_datain = ( (|r_sys_processing_methodID) ? r_sub09_result_datain : 32'h0 ) ;
	assign w_sub09_result_r_w = ( (|r_sys_processing_methodID) ? r_sub09_result_r_w : 1'h0 ) ;
	assign w_sub08_u_addr = ( (|r_sys_processing_methodID) ? r_sub08_u_addr : 13'sh0 ) ;
	assign w_sub08_u_datain = ( (|r_sys_processing_methodID) ? r_sub08_u_datain : 32'h0 ) ;
	assign w_sub08_u_r_w = ( (|r_sys_processing_methodID) ? r_sub08_u_r_w : 1'h0 ) ;
	assign w_sub08_result_addr = ( (|r_sys_processing_methodID) ? r_sub08_result_addr : 13'sh0 ) ;
	assign w_sub08_result_datain = ( (|r_sys_processing_methodID) ? r_sub08_result_datain : 32'h0 ) ;
	assign w_sub08_result_r_w = ( (|r_sys_processing_methodID) ? r_sub08_result_r_w : 1'h0 ) ;
	assign w_sub12_u_addr = ( (|r_sys_processing_methodID) ? r_sub12_u_addr : 13'sh0 ) ;
	assign w_sub12_u_datain = ( (|r_sys_processing_methodID) ? r_sub12_u_datain : 32'h0 ) ;
	assign w_sub12_u_r_w = ( (|r_sys_processing_methodID) ? r_sub12_u_r_w : 1'h0 ) ;
	assign w_sub12_result_addr = ( (|r_sys_processing_methodID) ? r_sub12_result_addr : 13'sh0 ) ;
	assign w_sub12_result_datain = ( (|r_sys_processing_methodID) ? r_sub12_result_datain : 32'h0 ) ;
	assign w_sub12_result_r_w = ( (|r_sys_processing_methodID) ? r_sub12_result_r_w : 1'h0 ) ;
	assign w_sub03_u_addr = ( (|r_sys_processing_methodID) ? r_sub03_u_addr : 13'sh0 ) ;
	assign w_sub03_u_datain = ( (|r_sys_processing_methodID) ? r_sub03_u_datain : 32'h0 ) ;
	assign w_sub03_u_r_w = ( (|r_sys_processing_methodID) ? r_sub03_u_r_w : 1'h0 ) ;
	assign w_sub03_result_addr = ( (|r_sys_processing_methodID) ? r_sub03_result_addr : 13'sh0 ) ;
	assign w_sub03_result_datain = ( (|r_sys_processing_methodID) ? r_sub03_result_datain : 32'h0 ) ;
	assign w_sub03_result_r_w = ( (|r_sys_processing_methodID) ? r_sub03_result_r_w : 1'h0 ) ;
	assign w_sub02_u_addr = ( (|r_sys_processing_methodID) ? r_sub02_u_addr : 13'sh0 ) ;
	assign w_sub02_u_datain = ( (|r_sys_processing_methodID) ? r_sub02_u_datain : 32'h0 ) ;
	assign w_sub02_u_r_w = ( (|r_sys_processing_methodID) ? r_sub02_u_r_w : 1'h0 ) ;
	assign w_sub02_result_addr = ( (|r_sys_processing_methodID) ? r_sub02_result_addr : 13'sh0 ) ;
	assign w_sub02_result_datain = ( (|r_sys_processing_methodID) ? r_sub02_result_datain : 32'h0 ) ;
	assign w_sub02_result_r_w = ( (|r_sys_processing_methodID) ? r_sub02_result_r_w : 1'h0 ) ;
	assign w_sub11_u_addr = ( (|r_sys_processing_methodID) ? r_sub11_u_addr : 13'sh0 ) ;
	assign w_sub11_u_datain = ( (|r_sys_processing_methodID) ? r_sub11_u_datain : 32'h0 ) ;
	assign w_sub11_u_r_w = ( (|r_sys_processing_methodID) ? r_sub11_u_r_w : 1'h0 ) ;
	assign w_sub11_result_addr = ( (|r_sys_processing_methodID) ? r_sub11_result_addr : 13'sh0 ) ;
	assign w_sub11_result_datain = ( (|r_sys_processing_methodID) ? r_sub11_result_datain : 32'h0 ) ;
	assign w_sub11_result_r_w = ( (|r_sys_processing_methodID) ? r_sub11_result_r_w : 1'h0 ) ;
	assign w_sub14_u_addr = ( (|r_sys_processing_methodID) ? r_sub14_u_addr : 13'sh0 ) ;
	assign w_sub14_u_datain = ( (|r_sys_processing_methodID) ? r_sub14_u_datain : 32'h0 ) ;
	assign w_sub14_u_r_w = ( (|r_sys_processing_methodID) ? r_sub14_u_r_w : 1'h0 ) ;
	assign w_sub14_result_addr = ( (|r_sys_processing_methodID) ? r_sub14_result_addr : 13'sh0 ) ;
	assign w_sub14_result_datain = ( (|r_sys_processing_methodID) ? r_sub14_result_datain : 32'h0 ) ;
	assign w_sub14_result_r_w = ( (|r_sys_processing_methodID) ? r_sub14_result_r_w : 1'h0 ) ;
	assign w_sub01_u_addr = ( (|r_sys_processing_methodID) ? r_sub01_u_addr : 13'sh0 ) ;
	assign w_sub01_u_datain = ( (|r_sys_processing_methodID) ? r_sub01_u_datain : 32'h0 ) ;
	assign w_sub01_u_r_w = ( (|r_sys_processing_methodID) ? r_sub01_u_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 13'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub13_u_addr = ( (|r_sys_processing_methodID) ? r_sub13_u_addr : 13'sh0 ) ;
	assign w_sub13_u_datain = ( (|r_sys_processing_methodID) ? r_sub13_u_datain : 32'h0 ) ;
	assign w_sub13_u_r_w = ( (|r_sys_processing_methodID) ? r_sub13_u_r_w : 1'h0 ) ;
	assign w_sub13_result_addr = ( (|r_sys_processing_methodID) ? r_sub13_result_addr : 13'sh0 ) ;
	assign w_sub13_result_datain = ( (|r_sys_processing_methodID) ? r_sub13_result_datain : 32'h0 ) ;
	assign w_sub13_result_r_w = ( (|r_sys_processing_methodID) ? r_sub13_result_r_w : 1'h0 ) ;
	assign w_sub00_u_addr = ( (|r_sys_processing_methodID) ? r_sub00_u_addr : 13'sh0 ) ;
	assign w_sub00_u_datain = ( (|r_sys_processing_methodID) ? r_sub00_u_datain : 32'h0 ) ;
	assign w_sub00_u_r_w = ( (|r_sys_processing_methodID) ? r_sub00_u_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 13'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sub07_u_addr = ( (|r_sys_processing_methodID) ? r_sub07_u_addr : 13'sh0 ) ;
	assign w_sub07_u_datain = ( (|r_sys_processing_methodID) ? r_sub07_u_datain : 32'h0 ) ;
	assign w_sub07_u_r_w = ( (|r_sys_processing_methodID) ? r_sub07_u_r_w : 1'h0 ) ;
	assign w_sub07_result_addr = ( (|r_sys_processing_methodID) ? r_sub07_result_addr : 13'sh0 ) ;
	assign w_sub07_result_datain = ( (|r_sys_processing_methodID) ? r_sub07_result_datain : 32'h0 ) ;
	assign w_sub07_result_r_w = ( (|r_sys_processing_methodID) ? r_sub07_result_r_w : 1'h0 ) ;
	assign w_sub06_u_addr = ( (|r_sys_processing_methodID) ? r_sub06_u_addr : 13'sh0 ) ;
	assign w_sub06_u_datain = ( (|r_sys_processing_methodID) ? r_sub06_u_datain : 32'h0 ) ;
	assign w_sub06_u_r_w = ( (|r_sys_processing_methodID) ? r_sub06_u_r_w : 1'h0 ) ;
	assign w_sub06_result_addr = ( (|r_sys_processing_methodID) ? r_sub06_result_addr : 13'sh0 ) ;
	assign w_sub06_result_datain = ( (|r_sys_processing_methodID) ? r_sub06_result_datain : 32'h0 ) ;
	assign w_sub06_result_r_w = ( (|r_sys_processing_methodID) ? r_sub06_result_r_w : 1'h0 ) ;
	assign w_sub15_u_addr = ( (|r_sys_processing_methodID) ? r_sub15_u_addr : 13'sh0 ) ;
	assign w_sub15_u_datain = ( (|r_sys_processing_methodID) ? r_sub15_u_datain : 32'h0 ) ;
	assign w_sub15_u_r_w = ( (|r_sys_processing_methodID) ? r_sub15_u_r_w : 1'h0 ) ;
	assign w_sub15_result_addr = ( (|r_sys_processing_methodID) ? r_sub15_result_addr : 13'sh0 ) ;
	assign w_sub15_result_datain = ( (|r_sys_processing_methodID) ? r_sub15_result_datain : 32'h0 ) ;
	assign w_sub15_result_r_w = ( (|r_sys_processing_methodID) ? r_sub15_result_r_w : 1'h0 ) ;
	assign w_sub05_u_addr = ( (|r_sys_processing_methodID) ? r_sub05_u_addr : 13'sh0 ) ;
	assign w_sub05_u_datain = ( (|r_sys_processing_methodID) ? r_sub05_u_datain : 32'h0 ) ;
	assign w_sub05_u_r_w = ( (|r_sys_processing_methodID) ? r_sub05_u_r_w : 1'h0 ) ;
	assign w_sub05_result_addr = ( (|r_sys_processing_methodID) ? r_sub05_result_addr : 13'sh0 ) ;
	assign w_sub05_result_datain = ( (|r_sys_processing_methodID) ? r_sub05_result_datain : 32'h0 ) ;
	assign w_sub05_result_r_w = ( (|r_sys_processing_methodID) ? r_sub05_result_r_w : 1'h0 ) ;
	assign w_sub04_u_addr = ( (|r_sys_processing_methodID) ? r_sub04_u_addr : 13'sh0 ) ;
	assign w_sub04_u_datain = ( (|r_sys_processing_methodID) ? r_sub04_u_datain : 32'h0 ) ;
	assign w_sub04_u_r_w = ( (|r_sys_processing_methodID) ? r_sub04_u_r_w : 1'h0 ) ;
	assign w_sub04_result_addr = ( (|r_sys_processing_methodID) ? r_sub04_result_addr : 13'sh0 ) ;
	assign w_sub04_result_datain = ( (|r_sys_processing_methodID) ? r_sub04_result_datain : 32'h0 ) ;
	assign w_sub04_result_r_w = ( (|r_sys_processing_methodID) ? r_sub04_result_r_w : 1'h0 ) ;
	assign w_sub10_u_addr = ( (|r_sys_processing_methodID) ? r_sub10_u_addr : 13'sh0 ) ;
	assign w_sub10_u_datain = ( (|r_sys_processing_methodID) ? r_sub10_u_datain : 32'h0 ) ;
	assign w_sub10_u_r_w = ( (|r_sys_processing_methodID) ? r_sub10_u_r_w : 1'h0 ) ;
	assign w_sub10_result_addr = ( (|r_sys_processing_methodID) ? r_sub10_result_addr : 13'sh0 ) ;
	assign w_sub10_result_datain = ( (|r_sys_processing_methodID) ? r_sub10_result_datain : 32'h0 ) ;
	assign w_sub10_result_r_w = ( (|r_sys_processing_methodID) ? r_sub10_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh00000081;
	assign w_sys_tmp3 = 32'sh00000002;
	assign w_sys_tmp4 = ( !w_sys_tmp5 );
	assign w_sys_tmp5 = (r_run_my_21 < r_run_k_17);
	assign w_sys_tmp6 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp7 = ( !w_sys_tmp8 );
	assign w_sys_tmp8 = (r_run_mx_20 < r_run_j_18);
	assign w_sys_tmp11 = (w_sys_tmp12 + r_run_k_17);
	assign w_sys_tmp12 = (r_run_j_18 * w_sys_tmp13);
	assign w_sys_tmp13 = 32'sh00000081;
	assign w_sys_tmp14 = 32'h0;
	assign w_sys_tmp15 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp52 = ( !w_sys_tmp53 );
	assign w_sys_tmp53 = (w_sys_tmp54 < r_run_k_17);
	assign w_sys_tmp54 = 32'sh00000021;
	assign w_sys_tmp55 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp56 = ( !w_sys_tmp57 );
	assign w_sys_tmp57 = (w_sys_tmp58 < r_run_j_18);
	assign w_sys_tmp58 = 32'sh00000021;
	assign w_sys_tmp61 = (w_sys_tmp62 + r_run_k_17);
	assign w_sys_tmp62 = (r_run_j_18 * w_sys_tmp63);
	assign w_sys_tmp63 = 32'sh00000081;
	assign w_sys_tmp64 = w_fld_u_0_dataout_1;
	assign w_sys_tmp65 = (w_sys_tmp66 + r_run_k_17);
	assign w_sys_tmp66 = (r_run_copy0_j_23 * w_sys_tmp63);
	assign w_sys_tmp68 = (r_run_copy0_j_23 + w_sys_intOne);
	assign w_sys_tmp69 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp130 = 32'sh00000020;
	assign w_sys_tmp131 = ( !w_sys_tmp132 );
	assign w_sys_tmp132 = (w_sys_tmp133 < r_run_j_18);
	assign w_sys_tmp133 = 32'sh00000041;
	assign w_sys_tmp136 = (w_sys_tmp137 + r_run_k_17);
	assign w_sys_tmp137 = (r_run_j_18 * w_sys_tmp138);
	assign w_sys_tmp138 = 32'sh00000081;
	assign w_sys_tmp139 = w_fld_u_0_dataout_1;
	assign w_sys_tmp140 = (w_sys_tmp141 + r_run_k_17);
	assign w_sys_tmp141 = (r_run_copy0_j_24 - w_sys_tmp142);
	assign w_sys_tmp142 = 32'sh00000f9f;
	assign w_sys_tmp143 = (r_run_copy0_j_24 + w_sys_intOne);
	assign w_sys_tmp144 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp205 = 32'sh00000040;
	assign w_sys_tmp206 = ( !w_sys_tmp207 );
	assign w_sys_tmp207 = (w_sys_tmp208 < r_run_j_18);
	assign w_sys_tmp208 = 32'sh00000061;
	assign w_sys_tmp211 = (w_sys_tmp212 + r_run_k_17);
	assign w_sys_tmp212 = (r_run_j_18 * w_sys_tmp213);
	assign w_sys_tmp213 = 32'sh00000081;
	assign w_sys_tmp214 = w_fld_u_0_dataout_1;
	assign w_sys_tmp215 = (w_sys_tmp216 + r_run_k_17);
	assign w_sys_tmp216 = (r_run_copy0_j_25 * w_sys_tmp213);
	assign w_sys_tmp218 = (r_run_copy0_j_25 + w_sys_intOne);
	assign w_sys_tmp219 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp280 = 32'sh00000060;
	assign w_sys_tmp281 = ( !w_sys_tmp282 );
	assign w_sys_tmp282 = (w_sys_tmp283 < r_run_j_18);
	assign w_sys_tmp283 = 32'sh00000081;
	assign w_sys_tmp286 = (w_sys_tmp287 + r_run_k_17);
	assign w_sys_tmp287 = (r_run_j_18 * w_sys_tmp288);
	assign w_sys_tmp288 = 32'sh00000081;
	assign w_sys_tmp289 = w_fld_u_0_dataout_1;
	assign w_sys_tmp290 = (w_sys_tmp291 + r_run_k_17);
	assign w_sys_tmp291 = (r_run_copy0_j_26 * w_sys_tmp288);
	assign w_sys_tmp293 = (r_run_copy0_j_26 + w_sys_intOne);
	assign w_sys_tmp294 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp355 = 32'sh00000020;
	assign w_sys_tmp356 = ( !w_sys_tmp357 );
	assign w_sys_tmp357 = (w_sys_tmp358 < r_run_k_17);
	assign w_sys_tmp358 = 32'sh00000041;
	assign w_sys_tmp359 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp360 = ( !w_sys_tmp361 );
	assign w_sys_tmp361 = (w_sys_tmp362 < r_run_j_18);
	assign w_sys_tmp362 = 32'sh00000021;
	assign w_sys_tmp365 = (w_sys_tmp366 + r_run_k_17);
	assign w_sys_tmp366 = (r_run_j_18 * w_sys_tmp367);
	assign w_sys_tmp367 = 32'sh00000081;
	assign w_sys_tmp368 = w_fld_u_0_dataout_1;
	assign w_sys_tmp369 = (w_sys_tmp370 + r_run_k_17);
	assign w_sys_tmp370 = (r_run_copy0_j_27 * w_sys_tmp367);
	assign w_sys_tmp372 = (r_run_copy0_j_27 + w_sys_intOne);
	assign w_sys_tmp373 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp434 = 32'sh00000020;
	assign w_sys_tmp435 = ( !w_sys_tmp436 );
	assign w_sys_tmp436 = (w_sys_tmp437 < r_run_j_18);
	assign w_sys_tmp437 = 32'sh00000041;
	assign w_sys_tmp440 = (w_sys_tmp441 + r_run_k_17);
	assign w_sys_tmp441 = (r_run_j_18 * w_sys_tmp442);
	assign w_sys_tmp442 = 32'sh00000081;
	assign w_sys_tmp443 = w_fld_u_0_dataout_1;
	assign w_sys_tmp444 = (w_sys_tmp445 + r_run_k_17);
	assign w_sys_tmp445 = (r_run_copy0_j_28 * w_sys_tmp442);
	assign w_sys_tmp447 = (r_run_copy0_j_28 + w_sys_intOne);
	assign w_sys_tmp448 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp509 = 32'sh00000040;
	assign w_sys_tmp510 = ( !w_sys_tmp511 );
	assign w_sys_tmp511 = (w_sys_tmp512 < r_run_j_18);
	assign w_sys_tmp512 = 32'sh00000061;
	assign w_sys_tmp515 = (w_sys_tmp516 + r_run_k_17);
	assign w_sys_tmp516 = (r_run_j_18 * w_sys_tmp517);
	assign w_sys_tmp517 = 32'sh00000081;
	assign w_sys_tmp518 = w_fld_u_0_dataout_1;
	assign w_sys_tmp519 = (w_sys_tmp520 + r_run_k_17);
	assign w_sys_tmp520 = (r_run_copy0_j_29 * w_sys_tmp517);
	assign w_sys_tmp522 = (r_run_copy0_j_29 + w_sys_intOne);
	assign w_sys_tmp523 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp584 = 32'sh00000060;
	assign w_sys_tmp585 = ( !w_sys_tmp586 );
	assign w_sys_tmp586 = (w_sys_tmp587 < r_run_j_18);
	assign w_sys_tmp587 = 32'sh00000081;
	assign w_sys_tmp590 = (w_sys_tmp591 + r_run_k_17);
	assign w_sys_tmp591 = (r_run_j_18 * w_sys_tmp592);
	assign w_sys_tmp592 = 32'sh00000081;
	assign w_sys_tmp593 = w_fld_u_0_dataout_1;
	assign w_sys_tmp594 = (w_sys_tmp595 + r_run_k_17);
	assign w_sys_tmp595 = (r_run_copy0_j_30 * w_sys_tmp592);
	assign w_sys_tmp597 = (r_run_copy0_j_30 + w_sys_intOne);
	assign w_sys_tmp598 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp659 = 32'sh00000040;
	assign w_sys_tmp660 = ( !w_sys_tmp661 );
	assign w_sys_tmp661 = (w_sys_tmp662 < r_run_k_17);
	assign w_sys_tmp662 = 32'sh00000061;
	assign w_sys_tmp663 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp664 = ( !w_sys_tmp665 );
	assign w_sys_tmp665 = (w_sys_tmp666 < r_run_j_18);
	assign w_sys_tmp666 = 32'sh00000021;
	assign w_sys_tmp669 = (w_sys_tmp670 + r_run_k_17);
	assign w_sys_tmp670 = (r_run_j_18 * w_sys_tmp671);
	assign w_sys_tmp671 = 32'sh00000081;
	assign w_sys_tmp672 = w_fld_u_0_dataout_1;
	assign w_sys_tmp673 = (w_sys_tmp674 + r_run_k_17);
	assign w_sys_tmp674 = (r_run_copy0_j_31 * w_sys_tmp671);
	assign w_sys_tmp676 = (r_run_copy0_j_31 + w_sys_intOne);
	assign w_sys_tmp677 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp738 = 32'sh00000020;
	assign w_sys_tmp739 = ( !w_sys_tmp740 );
	assign w_sys_tmp740 = (w_sys_tmp741 < r_run_j_18);
	assign w_sys_tmp741 = 32'sh00000041;
	assign w_sys_tmp744 = (w_sys_tmp745 + r_run_k_17);
	assign w_sys_tmp745 = (r_run_j_18 * w_sys_tmp746);
	assign w_sys_tmp746 = 32'sh00000081;
	assign w_sys_tmp747 = w_fld_u_0_dataout_1;
	assign w_sys_tmp748 = (w_sys_tmp749 + r_run_k_17);
	assign w_sys_tmp749 = (r_run_copy0_j_32 * w_sys_tmp746);
	assign w_sys_tmp751 = (r_run_copy0_j_32 + w_sys_intOne);
	assign w_sys_tmp752 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp813 = 32'sh00000040;
	assign w_sys_tmp814 = ( !w_sys_tmp815 );
	assign w_sys_tmp815 = (w_sys_tmp816 < r_run_j_18);
	assign w_sys_tmp816 = 32'sh00000061;
	assign w_sys_tmp819 = (w_sys_tmp820 + r_run_k_17);
	assign w_sys_tmp820 = (r_run_j_18 * w_sys_tmp821);
	assign w_sys_tmp821 = 32'sh00000081;
	assign w_sys_tmp822 = w_fld_u_0_dataout_1;
	assign w_sys_tmp823 = (w_sys_tmp824 + r_run_k_17);
	assign w_sys_tmp824 = (r_run_copy0_j_33 * w_sys_tmp821);
	assign w_sys_tmp826 = (r_run_copy0_j_33 + w_sys_intOne);
	assign w_sys_tmp827 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp888 = 32'sh00000060;
	assign w_sys_tmp889 = ( !w_sys_tmp890 );
	assign w_sys_tmp890 = (w_sys_tmp891 < r_run_j_18);
	assign w_sys_tmp891 = 32'sh00000081;
	assign w_sys_tmp894 = (w_sys_tmp895 + r_run_k_17);
	assign w_sys_tmp895 = (r_run_j_18 * w_sys_tmp896);
	assign w_sys_tmp896 = 32'sh00000081;
	assign w_sys_tmp897 = w_fld_u_0_dataout_1;
	assign w_sys_tmp898 = (w_sys_tmp899 + r_run_k_17);
	assign w_sys_tmp899 = (r_run_copy0_j_34 * w_sys_tmp896);
	assign w_sys_tmp901 = (r_run_copy0_j_34 + w_sys_intOne);
	assign w_sys_tmp902 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp963 = 32'sh00000060;
	assign w_sys_tmp964 = ( !w_sys_tmp965 );
	assign w_sys_tmp965 = (w_sys_tmp966 < r_run_k_17);
	assign w_sys_tmp966 = 32'sh00000081;
	assign w_sys_tmp967 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp968 = ( !w_sys_tmp969 );
	assign w_sys_tmp969 = (w_sys_tmp970 < r_run_j_18);
	assign w_sys_tmp970 = 32'sh00000021;
	assign w_sys_tmp973 = (w_sys_tmp974 + r_run_k_17);
	assign w_sys_tmp974 = (r_run_j_18 * w_sys_tmp975);
	assign w_sys_tmp975 = 32'sh00000081;
	assign w_sys_tmp976 = w_fld_u_0_dataout_1;
	assign w_sys_tmp977 = (w_sys_tmp978 + r_run_k_17);
	assign w_sys_tmp978 = (r_run_copy0_j_35 * w_sys_tmp975);
	assign w_sys_tmp980 = (r_run_copy0_j_35 + w_sys_intOne);
	assign w_sys_tmp981 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp1042 = 32'sh00000020;
	assign w_sys_tmp1043 = ( !w_sys_tmp1044 );
	assign w_sys_tmp1044 = (w_sys_tmp1045 < r_run_j_18);
	assign w_sys_tmp1045 = 32'sh00000041;
	assign w_sys_tmp1048 = (w_sys_tmp1049 + r_run_k_17);
	assign w_sys_tmp1049 = (r_run_j_18 * w_sys_tmp1050);
	assign w_sys_tmp1050 = 32'sh00000081;
	assign w_sys_tmp1051 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1052 = (w_sys_tmp1053 + r_run_k_17);
	assign w_sys_tmp1053 = (r_run_copy0_j_36 * w_sys_tmp1050);
	assign w_sys_tmp1055 = (r_run_copy0_j_36 + w_sys_intOne);
	assign w_sys_tmp1056 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp1117 = 32'sh00000040;
	assign w_sys_tmp1118 = ( !w_sys_tmp1119 );
	assign w_sys_tmp1119 = (w_sys_tmp1120 < r_run_j_18);
	assign w_sys_tmp1120 = 32'sh00000061;
	assign w_sys_tmp1123 = (w_sys_tmp1124 + r_run_k_17);
	assign w_sys_tmp1124 = (r_run_j_18 * w_sys_tmp1125);
	assign w_sys_tmp1125 = 32'sh00000081;
	assign w_sys_tmp1126 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1127 = (w_sys_tmp1128 + r_run_k_17);
	assign w_sys_tmp1128 = (r_run_copy0_j_37 * w_sys_tmp1125);
	assign w_sys_tmp1130 = (r_run_copy0_j_37 + w_sys_intOne);
	assign w_sys_tmp1131 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp1192 = 32'sh00000060;
	assign w_sys_tmp1193 = ( !w_sys_tmp1194 );
	assign w_sys_tmp1194 = (w_sys_tmp1195 < r_run_j_18);
	assign w_sys_tmp1195 = 32'sh00000081;
	assign w_sys_tmp1198 = (w_sys_tmp1199 + r_run_k_17);
	assign w_sys_tmp1199 = (r_run_j_18 * w_sys_tmp1200);
	assign w_sys_tmp1200 = 32'sh00000081;
	assign w_sys_tmp1201 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1202 = (w_sys_tmp1203 + r_run_k_17);
	assign w_sys_tmp1203 = (r_run_copy0_j_38 * w_sys_tmp1200);
	assign w_sys_tmp1205 = (r_run_copy0_j_38 + w_sys_intOne);
	assign w_sys_tmp1206 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp1267 = ( !w_sys_tmp1268 );
	assign w_sys_tmp1268 = (r_run_nlast_22 < r_run_n_19);
	assign w_sys_tmp1269 = (r_run_n_19 + w_sys_intOne);
	assign w_sys_tmp1270 = 32'sh00000002;
	assign w_sys_tmp1271 = ( !w_sys_tmp1272 );
	assign w_sys_tmp1272 = (w_sys_tmp1273 < r_run_k_17);
	assign w_sys_tmp1273 = 32'sh00000020;
	assign w_sys_tmp1276 = (w_sys_tmp1277 + r_run_k_17);
	assign w_sys_tmp1277 = 32'sh000010a1;
	assign w_sys_tmp1278 = w_sub04_result_dataout;
	assign w_sys_tmp1282 = (w_sys_tmp1283 + r_run_k_17);
	assign w_sys_tmp1283 = 32'sh00001020;
	assign w_sys_tmp1284 = w_sub00_result_dataout;
	assign w_sys_tmp1288 = (w_sys_tmp1289 + r_run_k_17);
	assign w_sys_tmp1289 = 32'sh000020c1;
	assign w_sys_tmp1293 = (w_sys_tmp1294 + r_run_k_17);
	assign w_sys_tmp1294 = 32'sh00002040;
	assign w_sys_tmp1299 = (w_sys_tmp1300 + r_run_k_17);
	assign w_sys_tmp1300 = 32'sh000030e1;
	assign w_sys_tmp1304 = (w_sys_tmp1305 + r_run_k_17);
	assign w_sys_tmp1305 = 32'sh00003060;
	assign w_sys_tmp1306 = w_sub08_result_dataout;
	assign w_sys_tmp1309 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp1310 = 32'sh00000021;
	assign w_sys_tmp1311 = ( !w_sys_tmp1312 );
	assign w_sys_tmp1312 = (w_sys_tmp1313 < r_run_k_17);
	assign w_sys_tmp1313 = 32'sh00000040;
	assign w_sys_tmp1316 = (w_sys_tmp1317 + r_run_k_17);
	assign w_sys_tmp1317 = 32'sh000010a1;
	assign w_sys_tmp1318 = w_sub05_result_dataout;
	assign w_sys_tmp1322 = (w_sys_tmp1323 + r_run_k_17);
	assign w_sys_tmp1323 = 32'sh00001020;
	assign w_sys_tmp1324 = w_sub01_result_dataout;
	assign w_sys_tmp1328 = (w_sys_tmp1329 + r_run_k_17);
	assign w_sys_tmp1329 = 32'sh000020c1;
	assign w_sys_tmp1333 = (w_sys_tmp1334 + r_run_k_17);
	assign w_sys_tmp1334 = 32'sh00002040;
	assign w_sys_tmp1339 = (w_sys_tmp1340 + r_run_k_17);
	assign w_sys_tmp1340 = 32'sh000030e1;
	assign w_sys_tmp1344 = (w_sys_tmp1345 + r_run_k_17);
	assign w_sys_tmp1345 = 32'sh00003060;
	assign w_sys_tmp1346 = w_sub09_result_dataout;
	assign w_sys_tmp1349 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp1350 = 32'sh00000041;
	assign w_sys_tmp1351 = ( !w_sys_tmp1352 );
	assign w_sys_tmp1352 = (w_sys_tmp1353 < r_run_k_17);
	assign w_sys_tmp1353 = 32'sh00000060;
	assign w_sys_tmp1356 = (w_sys_tmp1357 + r_run_k_17);
	assign w_sys_tmp1357 = 32'sh000010a1;
	assign w_sys_tmp1358 = w_sub06_result_dataout;
	assign w_sys_tmp1362 = (w_sys_tmp1363 + r_run_k_17);
	assign w_sys_tmp1363 = 32'sh00001020;
	assign w_sys_tmp1364 = w_sub02_result_dataout;
	assign w_sys_tmp1368 = (w_sys_tmp1369 + r_run_k_17);
	assign w_sys_tmp1369 = 32'sh000020c1;
	assign w_sys_tmp1373 = (w_sys_tmp1374 + r_run_k_17);
	assign w_sys_tmp1374 = 32'sh00002040;
	assign w_sys_tmp1379 = (w_sys_tmp1380 + r_run_k_17);
	assign w_sys_tmp1380 = 32'sh000030e1;
	assign w_sys_tmp1384 = (w_sys_tmp1385 + r_run_k_17);
	assign w_sys_tmp1385 = 32'sh00003060;
	assign w_sys_tmp1386 = w_sub10_result_dataout;
	assign w_sys_tmp1389 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp1390 = 32'sh00000061;
	assign w_sys_tmp1391 = ( !w_sys_tmp1392 );
	assign w_sys_tmp1392 = (w_sys_tmp1393 < r_run_k_17);
	assign w_sys_tmp1393 = 32'sh00000080;
	assign w_sys_tmp1396 = (w_sys_tmp1397 + r_run_k_17);
	assign w_sys_tmp1397 = 32'sh000010a1;
	assign w_sys_tmp1398 = w_sub07_result_dataout;
	assign w_sys_tmp1402 = (w_sys_tmp1403 + r_run_k_17);
	assign w_sys_tmp1403 = 32'sh00001020;
	assign w_sys_tmp1404 = w_sub03_result_dataout;
	assign w_sys_tmp1408 = (w_sys_tmp1409 + r_run_k_17);
	assign w_sys_tmp1409 = 32'sh000020c1;
	assign w_sys_tmp1413 = (w_sys_tmp1414 + r_run_k_17);
	assign w_sys_tmp1414 = 32'sh00002040;
	assign w_sys_tmp1419 = (w_sys_tmp1420 + r_run_k_17);
	assign w_sys_tmp1420 = 32'sh000030e1;
	assign w_sys_tmp1424 = (w_sys_tmp1425 + r_run_k_17);
	assign w_sys_tmp1425 = 32'sh00003060;
	assign w_sys_tmp1426 = w_sub11_result_dataout;
	assign w_sys_tmp1429 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp1430 = 32'sh00000002;
	assign w_sys_tmp1431 = ( !w_sys_tmp1432 );
	assign w_sys_tmp1432 = (w_sys_tmp1433 < r_run_j_18);
	assign w_sys_tmp1433 = 32'sh00000020;
	assign w_sys_tmp1436 = (w_sys_tmp1437 + w_sys_tmp1439);
	assign w_sys_tmp1437 = (r_run_j_18 * w_sys_tmp1438);
	assign w_sys_tmp1438 = 32'sh00000081;
	assign w_sys_tmp1439 = 32'sh00000021;
	assign w_sys_tmp1440 = w_sub01_result_dataout;
	assign w_sys_tmp1441 = (w_sys_tmp1442 + w_sys_tmp1439);
	assign w_sys_tmp1442 = (r_run_copy10_j_49 * w_sys_tmp1438);
	assign w_sys_tmp1446 = (w_sys_tmp1447 + w_sys_tmp1449);
	assign w_sys_tmp1447 = (r_run_copy9_j_48 * w_sys_tmp1438);
	assign w_sys_tmp1449 = 32'sh00000020;
	assign w_sys_tmp1450 = w_sub00_result_dataout;
	assign w_sys_tmp1451 = (w_sys_tmp1452 + w_sys_tmp1449);
	assign w_sys_tmp1452 = (r_run_copy8_j_47 * w_sys_tmp1438);
	assign w_sys_tmp1456 = (w_sys_tmp1457 + w_sys_tmp1459);
	assign w_sys_tmp1457 = (r_run_copy7_j_46 * w_sys_tmp1438);
	assign w_sys_tmp1459 = 32'sh00000041;
	assign w_sys_tmp1460 = (w_sys_tmp1461 + w_sys_tmp1459);
	assign w_sys_tmp1461 = (r_run_copy6_j_45 * w_sys_tmp1438);
	assign w_sys_tmp1465 = (w_sys_tmp1466 + w_sys_tmp1468);
	assign w_sys_tmp1466 = (r_run_copy5_j_44 * w_sys_tmp1438);
	assign w_sys_tmp1468 = 32'sh00000040;
	assign w_sys_tmp1470 = (w_sys_tmp1471 + w_sys_tmp1468);
	assign w_sys_tmp1471 = (r_run_copy4_j_43 * w_sys_tmp1438);
	assign w_sys_tmp1475 = (w_sys_tmp1476 + w_sys_tmp1478);
	assign w_sys_tmp1476 = (r_run_copy3_j_42 * w_sys_tmp1438);
	assign w_sys_tmp1478 = 32'sh00000061;
	assign w_sys_tmp1479 = (w_sys_tmp1480 + w_sys_tmp1478);
	assign w_sys_tmp1480 = (r_run_copy2_j_41 * w_sys_tmp1438);
	assign w_sys_tmp1484 = (w_sys_tmp1485 + w_sys_tmp1487);
	assign w_sys_tmp1485 = (r_run_copy1_j_40 * w_sys_tmp1438);
	assign w_sys_tmp1487 = 32'sh00000060;
	assign w_sys_tmp1488 = w_sub02_result_dataout;
	assign w_sys_tmp1489 = (w_sys_tmp1490 + w_sys_tmp1487);
	assign w_sys_tmp1490 = (r_run_copy0_j_39 * w_sys_tmp1438);
	assign w_sys_tmp1493 = (r_run_copy0_j_39 + w_sys_intOne);
	assign w_sys_tmp1494 = (r_run_copy1_j_40 + w_sys_intOne);
	assign w_sys_tmp1495 = (r_run_copy2_j_41 + w_sys_intOne);
	assign w_sys_tmp1496 = (r_run_copy3_j_42 + w_sys_intOne);
	assign w_sys_tmp1497 = (r_run_copy4_j_43 + w_sys_intOne);
	assign w_sys_tmp1498 = (r_run_copy5_j_44 + w_sys_intOne);
	assign w_sys_tmp1499 = (r_run_copy6_j_45 + w_sys_intOne);
	assign w_sys_tmp1500 = (r_run_copy7_j_46 + w_sys_intOne);
	assign w_sys_tmp1501 = (r_run_copy8_j_47 + w_sys_intOne);
	assign w_sys_tmp1502 = (r_run_copy9_j_48 + w_sys_intOne);
	assign w_sys_tmp1503 = (r_run_copy10_j_49 + w_sys_intOne);
	assign w_sys_tmp1504 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp1931 = 32'sh00000021;
	assign w_sys_tmp1932 = ( !w_sys_tmp1933 );
	assign w_sys_tmp1933 = (w_sys_tmp1934 < r_run_j_18);
	assign w_sys_tmp1934 = 32'sh00000040;
	assign w_sys_tmp1937 = (w_sys_tmp1938 + w_sys_tmp1940);
	assign w_sys_tmp1938 = (r_run_j_18 * w_sys_tmp1939);
	assign w_sys_tmp1939 = 32'sh00000081;
	assign w_sys_tmp1940 = 32'sh00000021;
	assign w_sys_tmp1941 = w_sub05_result_dataout;
	assign w_sys_tmp1942 = (w_sys_tmp1943 + w_sys_tmp1940);
	assign w_sys_tmp1943 = (r_run_copy10_j_60 * w_sys_tmp1939);
	assign w_sys_tmp1947 = (w_sys_tmp1948 + w_sys_tmp1950);
	assign w_sys_tmp1948 = (r_run_copy9_j_59 * w_sys_tmp1939);
	assign w_sys_tmp1950 = 32'sh00000020;
	assign w_sys_tmp1951 = w_sub04_result_dataout;
	assign w_sys_tmp1952 = (w_sys_tmp1953 + w_sys_tmp1950);
	assign w_sys_tmp1953 = (r_run_copy8_j_58 * w_sys_tmp1939);
	assign w_sys_tmp1957 = (w_sys_tmp1958 + w_sys_tmp1960);
	assign w_sys_tmp1958 = (r_run_copy7_j_57 * w_sys_tmp1939);
	assign w_sys_tmp1960 = 32'sh00000041;
	assign w_sys_tmp1961 = (w_sys_tmp1962 + w_sys_tmp1960);
	assign w_sys_tmp1962 = (r_run_copy6_j_56 * w_sys_tmp1939);
	assign w_sys_tmp1966 = (w_sys_tmp1967 + w_sys_tmp1969);
	assign w_sys_tmp1967 = (r_run_copy5_j_55 * w_sys_tmp1939);
	assign w_sys_tmp1969 = 32'sh00000040;
	assign w_sys_tmp1971 = (w_sys_tmp1972 + w_sys_tmp1969);
	assign w_sys_tmp1972 = (r_run_copy4_j_54 * w_sys_tmp1939);
	assign w_sys_tmp1976 = (w_sys_tmp1977 + w_sys_tmp1979);
	assign w_sys_tmp1977 = (r_run_copy3_j_53 * w_sys_tmp1939);
	assign w_sys_tmp1979 = 32'sh00000061;
	assign w_sys_tmp1980 = (w_sys_tmp1981 + w_sys_tmp1979);
	assign w_sys_tmp1981 = (r_run_copy2_j_52 * w_sys_tmp1939);
	assign w_sys_tmp1985 = (w_sys_tmp1986 + w_sys_tmp1988);
	assign w_sys_tmp1986 = (r_run_copy1_j_51 * w_sys_tmp1939);
	assign w_sys_tmp1988 = 32'sh00000060;
	assign w_sys_tmp1989 = w_sub06_result_dataout;
	assign w_sys_tmp1990 = (w_sys_tmp1991 + w_sys_tmp1988);
	assign w_sys_tmp1991 = (r_run_copy0_j_50 * w_sys_tmp1939);
	assign w_sys_tmp1994 = (r_run_copy0_j_50 + w_sys_intOne);
	assign w_sys_tmp1995 = (r_run_copy1_j_51 + w_sys_intOne);
	assign w_sys_tmp1996 = (r_run_copy2_j_52 + w_sys_intOne);
	assign w_sys_tmp1997 = (r_run_copy3_j_53 + w_sys_intOne);
	assign w_sys_tmp1998 = (r_run_copy4_j_54 + w_sys_intOne);
	assign w_sys_tmp1999 = (r_run_copy5_j_55 + w_sys_intOne);
	assign w_sys_tmp2000 = (r_run_copy6_j_56 + w_sys_intOne);
	assign w_sys_tmp2001 = (r_run_copy7_j_57 + w_sys_intOne);
	assign w_sys_tmp2002 = (r_run_copy8_j_58 + w_sys_intOne);
	assign w_sys_tmp2003 = (r_run_copy9_j_59 + w_sys_intOne);
	assign w_sys_tmp2004 = (r_run_copy10_j_60 + w_sys_intOne);
	assign w_sys_tmp2005 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp2432 = 32'sh00000041;
	assign w_sys_tmp2433 = ( !w_sys_tmp2434 );
	assign w_sys_tmp2434 = (w_sys_tmp2435 < r_run_j_18);
	assign w_sys_tmp2435 = 32'sh00000060;
	assign w_sys_tmp2438 = (w_sys_tmp2439 + w_sys_tmp2441);
	assign w_sys_tmp2439 = (r_run_j_18 * w_sys_tmp2440);
	assign w_sys_tmp2440 = 32'sh00000081;
	assign w_sys_tmp2441 = 32'sh00000021;
	assign w_sys_tmp2442 = w_sub09_result_dataout;
	assign w_sys_tmp2443 = (w_sys_tmp2444 + w_sys_tmp2441);
	assign w_sys_tmp2444 = (r_run_copy10_j_71 * w_sys_tmp2440);
	assign w_sys_tmp2448 = (w_sys_tmp2449 + w_sys_tmp2451);
	assign w_sys_tmp2449 = (r_run_copy9_j_70 * w_sys_tmp2440);
	assign w_sys_tmp2451 = 32'sh00000020;
	assign w_sys_tmp2452 = w_sub08_result_dataout;
	assign w_sys_tmp2453 = (w_sys_tmp2454 + w_sys_tmp2451);
	assign w_sys_tmp2454 = (r_run_copy8_j_69 * w_sys_tmp2440);
	assign w_sys_tmp2458 = (w_sys_tmp2459 + w_sys_tmp2461);
	assign w_sys_tmp2459 = (r_run_copy7_j_68 * w_sys_tmp2440);
	assign w_sys_tmp2461 = 32'sh00000041;
	assign w_sys_tmp2462 = (w_sys_tmp2463 + w_sys_tmp2461);
	assign w_sys_tmp2463 = (r_run_copy6_j_67 * w_sys_tmp2440);
	assign w_sys_tmp2467 = (w_sys_tmp2468 + w_sys_tmp2470);
	assign w_sys_tmp2468 = (r_run_copy5_j_66 * w_sys_tmp2440);
	assign w_sys_tmp2470 = 32'sh00000040;
	assign w_sys_tmp2472 = (w_sys_tmp2473 + w_sys_tmp2470);
	assign w_sys_tmp2473 = (r_run_copy4_j_65 * w_sys_tmp2440);
	assign w_sys_tmp2477 = (w_sys_tmp2478 + w_sys_tmp2480);
	assign w_sys_tmp2478 = (r_run_copy3_j_64 * w_sys_tmp2440);
	assign w_sys_tmp2480 = 32'sh00000061;
	assign w_sys_tmp2481 = (w_sys_tmp2482 + w_sys_tmp2480);
	assign w_sys_tmp2482 = (r_run_copy2_j_63 * w_sys_tmp2440);
	assign w_sys_tmp2486 = (w_sys_tmp2487 + w_sys_tmp2489);
	assign w_sys_tmp2487 = (r_run_copy1_j_62 * w_sys_tmp2440);
	assign w_sys_tmp2489 = 32'sh00000060;
	assign w_sys_tmp2490 = w_sub10_result_dataout;
	assign w_sys_tmp2491 = (w_sys_tmp2492 + w_sys_tmp2489);
	assign w_sys_tmp2492 = (r_run_copy0_j_61 * w_sys_tmp2440);
	assign w_sys_tmp2495 = (r_run_copy0_j_61 + w_sys_intOne);
	assign w_sys_tmp2496 = (r_run_copy1_j_62 + w_sys_intOne);
	assign w_sys_tmp2497 = (r_run_copy2_j_63 + w_sys_intOne);
	assign w_sys_tmp2498 = (r_run_copy3_j_64 + w_sys_intOne);
	assign w_sys_tmp2499 = (r_run_copy4_j_65 + w_sys_intOne);
	assign w_sys_tmp2500 = (r_run_copy5_j_66 + w_sys_intOne);
	assign w_sys_tmp2501 = (r_run_copy6_j_67 + w_sys_intOne);
	assign w_sys_tmp2502 = (r_run_copy7_j_68 + w_sys_intOne);
	assign w_sys_tmp2503 = (r_run_copy8_j_69 + w_sys_intOne);
	assign w_sys_tmp2504 = (r_run_copy9_j_70 + w_sys_intOne);
	assign w_sys_tmp2505 = (r_run_copy10_j_71 + w_sys_intOne);
	assign w_sys_tmp2506 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp2933 = 32'sh00000061;
	assign w_sys_tmp2934 = ( !w_sys_tmp2935 );
	assign w_sys_tmp2935 = (w_sys_tmp2936 < r_run_j_18);
	assign w_sys_tmp2936 = 32'sh00000080;
	assign w_sys_tmp2939 = (w_sys_tmp2940 + w_sys_tmp2942);
	assign w_sys_tmp2940 = (r_run_j_18 * w_sys_tmp2941);
	assign w_sys_tmp2941 = 32'sh00000081;
	assign w_sys_tmp2942 = 32'sh00000021;
	assign w_sys_tmp2943 = w_sub13_result_dataout;
	assign w_sys_tmp2944 = (w_sys_tmp2945 + w_sys_tmp2942);
	assign w_sys_tmp2945 = (r_run_copy10_j_82 * w_sys_tmp2941);
	assign w_sys_tmp2949 = (w_sys_tmp2950 + w_sys_tmp2952);
	assign w_sys_tmp2950 = (r_run_copy9_j_81 * w_sys_tmp2941);
	assign w_sys_tmp2952 = 32'sh00000020;
	assign w_sys_tmp2953 = w_sub12_result_dataout;
	assign w_sys_tmp2954 = (w_sys_tmp2955 + w_sys_tmp2952);
	assign w_sys_tmp2955 = (r_run_copy8_j_80 * w_sys_tmp2941);
	assign w_sys_tmp2959 = (w_sys_tmp2960 + w_sys_tmp2962);
	assign w_sys_tmp2960 = (r_run_copy7_j_79 * w_sys_tmp2941);
	assign w_sys_tmp2962 = 32'sh00000041;
	assign w_sys_tmp2963 = (w_sys_tmp2964 + w_sys_tmp2962);
	assign w_sys_tmp2964 = (r_run_copy6_j_78 * w_sys_tmp2941);
	assign w_sys_tmp2968 = (w_sys_tmp2969 + w_sys_tmp2971);
	assign w_sys_tmp2969 = (r_run_copy5_j_77 * w_sys_tmp2941);
	assign w_sys_tmp2971 = 32'sh00000040;
	assign w_sys_tmp2973 = (w_sys_tmp2974 + w_sys_tmp2971);
	assign w_sys_tmp2974 = (r_run_copy4_j_76 * w_sys_tmp2941);
	assign w_sys_tmp2978 = (w_sys_tmp2979 + w_sys_tmp2981);
	assign w_sys_tmp2979 = (r_run_copy3_j_75 * w_sys_tmp2941);
	assign w_sys_tmp2981 = 32'sh00000061;
	assign w_sys_tmp2982 = (w_sys_tmp2983 + w_sys_tmp2981);
	assign w_sys_tmp2983 = (r_run_copy2_j_74 * w_sys_tmp2941);
	assign w_sys_tmp2987 = (w_sys_tmp2988 + w_sys_tmp2990);
	assign w_sys_tmp2988 = (r_run_copy1_j_73 * w_sys_tmp2941);
	assign w_sys_tmp2990 = 32'sh00000060;
	assign w_sys_tmp2991 = w_sub14_result_dataout;
	assign w_sys_tmp2992 = (w_sys_tmp2993 + w_sys_tmp2990);
	assign w_sys_tmp2993 = (r_run_copy0_j_72 * w_sys_tmp2941);
	assign w_sys_tmp2996 = (r_run_copy0_j_72 + w_sys_intOne);
	assign w_sys_tmp2997 = (r_run_copy1_j_73 + w_sys_intOne);
	assign w_sys_tmp2998 = (r_run_copy2_j_74 + w_sys_intOne);
	assign w_sys_tmp2999 = (r_run_copy3_j_75 + w_sys_intOne);
	assign w_sys_tmp3000 = (r_run_copy4_j_76 + w_sys_intOne);
	assign w_sys_tmp3001 = (r_run_copy5_j_77 + w_sys_intOne);
	assign w_sys_tmp3002 = (r_run_copy6_j_78 + w_sys_intOne);
	assign w_sys_tmp3003 = (r_run_copy7_j_79 + w_sys_intOne);
	assign w_sys_tmp3004 = (r_run_copy8_j_80 + w_sys_intOne);
	assign w_sys_tmp3005 = (r_run_copy9_j_81 + w_sys_intOne);
	assign w_sys_tmp3006 = (r_run_copy10_j_82 + w_sys_intOne);
	assign w_sys_tmp3007 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp3434 = 32'sh00000002;
	assign w_sys_tmp3435 = ( !w_sys_tmp3436 );
	assign w_sys_tmp3436 = (w_sys_tmp3437 < r_run_k_17);
	assign w_sys_tmp3437 = 32'sh00000020;
	assign w_sys_tmp3438 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp3439 = 32'sh00000002;
	assign w_sys_tmp3440 = ( !w_sys_tmp3441 );
	assign w_sys_tmp3441 = (w_sys_tmp3442 < r_run_j_18);
	assign w_sys_tmp3442 = 32'sh00000020;
	assign w_sys_tmp3445 = (w_sys_tmp3446 + r_run_k_17);
	assign w_sys_tmp3446 = (r_run_j_18 * w_sys_tmp3447);
	assign w_sys_tmp3447 = 32'sh00000081;
	assign w_sys_tmp3448 = w_sub00_result_dataout;
	assign w_sys_tmp3449 = (w_sys_tmp3450 + r_run_k_17);
	assign w_sys_tmp3450 = (r_run_copy0_j_83 * w_sys_tmp3447);
	assign w_sys_tmp3452 = (r_run_copy0_j_83 + w_sys_intOne);
	assign w_sys_tmp3453 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp3514 = 32'sh00000021;
	assign w_sys_tmp3515 = ( !w_sys_tmp3516 );
	assign w_sys_tmp3516 = (w_sys_tmp3517 < r_run_j_18);
	assign w_sys_tmp3517 = 32'sh00000040;
	assign w_sys_tmp3520 = (w_sys_tmp3521 + r_run_k_17);
	assign w_sys_tmp3521 = (r_run_j_18 * w_sys_tmp3522);
	assign w_sys_tmp3522 = 32'sh00000081;
	assign w_sys_tmp3523 = w_sub01_result_dataout;
	assign w_sys_tmp3524 = (w_sys_tmp3525 + r_run_k_17);
	assign w_sys_tmp3525 = (r_run_copy0_j_84 * w_sys_tmp3522);
	assign w_sys_tmp3527 = (r_run_copy0_j_84 + w_sys_intOne);
	assign w_sys_tmp3528 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp3589 = 32'sh00000041;
	assign w_sys_tmp3590 = ( !w_sys_tmp3591 );
	assign w_sys_tmp3591 = (w_sys_tmp3592 < r_run_j_18);
	assign w_sys_tmp3592 = 32'sh00000060;
	assign w_sys_tmp3595 = (w_sys_tmp3596 + r_run_k_17);
	assign w_sys_tmp3596 = (r_run_j_18 * w_sys_tmp3597);
	assign w_sys_tmp3597 = 32'sh00000081;
	assign w_sys_tmp3598 = w_sub02_result_dataout;
	assign w_sys_tmp3599 = (w_sys_tmp3600 + r_run_k_17);
	assign w_sys_tmp3600 = (r_run_copy0_j_85 * w_sys_tmp3597);
	assign w_sys_tmp3602 = (r_run_copy0_j_85 + w_sys_intOne);
	assign w_sys_tmp3603 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp3664 = 32'sh00000061;
	assign w_sys_tmp3665 = ( !w_sys_tmp3666 );
	assign w_sys_tmp3666 = (w_sys_tmp3667 < r_run_j_18);
	assign w_sys_tmp3667 = 32'sh00000080;
	assign w_sys_tmp3670 = (w_sys_tmp3671 + r_run_k_17);
	assign w_sys_tmp3671 = (r_run_j_18 * w_sys_tmp3672);
	assign w_sys_tmp3672 = 32'sh00000081;
	assign w_sys_tmp3673 = w_sub03_result_dataout;
	assign w_sys_tmp3674 = (w_sys_tmp3675 + r_run_k_17);
	assign w_sys_tmp3675 = (r_run_copy0_j_86 * w_sys_tmp3672);
	assign w_sys_tmp3677 = (r_run_copy0_j_86 + w_sys_intOne);
	assign w_sys_tmp3678 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp3739 = 32'sh00000021;
	assign w_sys_tmp3740 = ( !w_sys_tmp3741 );
	assign w_sys_tmp3741 = (w_sys_tmp3742 < r_run_k_17);
	assign w_sys_tmp3742 = 32'sh00000040;
	assign w_sys_tmp3743 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp3744 = 32'sh00000002;
	assign w_sys_tmp3745 = ( !w_sys_tmp3746 );
	assign w_sys_tmp3746 = (w_sys_tmp3747 < r_run_j_18);
	assign w_sys_tmp3747 = 32'sh00000020;
	assign w_sys_tmp3750 = (w_sys_tmp3751 + r_run_k_17);
	assign w_sys_tmp3751 = (r_run_j_18 * w_sys_tmp3752);
	assign w_sys_tmp3752 = 32'sh00000081;
	assign w_sys_tmp3753 = w_sub04_result_dataout;
	assign w_sys_tmp3754 = (w_sys_tmp3755 + r_run_k_17);
	assign w_sys_tmp3755 = (r_run_copy0_j_87 * w_sys_tmp3752);
	assign w_sys_tmp3757 = (r_run_copy0_j_87 + w_sys_intOne);
	assign w_sys_tmp3758 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp3819 = 32'sh00000021;
	assign w_sys_tmp3820 = ( !w_sys_tmp3821 );
	assign w_sys_tmp3821 = (w_sys_tmp3822 < r_run_j_18);
	assign w_sys_tmp3822 = 32'sh00000040;
	assign w_sys_tmp3825 = (w_sys_tmp3826 + r_run_k_17);
	assign w_sys_tmp3826 = (r_run_j_18 * w_sys_tmp3827);
	assign w_sys_tmp3827 = 32'sh00000081;
	assign w_sys_tmp3828 = w_sub05_result_dataout;
	assign w_sys_tmp3829 = (w_sys_tmp3830 + r_run_k_17);
	assign w_sys_tmp3830 = (r_run_copy0_j_88 * w_sys_tmp3827);
	assign w_sys_tmp3832 = (r_run_copy0_j_88 + w_sys_intOne);
	assign w_sys_tmp3833 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp3894 = 32'sh00000041;
	assign w_sys_tmp3895 = ( !w_sys_tmp3896 );
	assign w_sys_tmp3896 = (w_sys_tmp3897 < r_run_j_18);
	assign w_sys_tmp3897 = 32'sh00000060;
	assign w_sys_tmp3900 = (w_sys_tmp3901 + r_run_k_17);
	assign w_sys_tmp3901 = (r_run_j_18 * w_sys_tmp3902);
	assign w_sys_tmp3902 = 32'sh00000081;
	assign w_sys_tmp3903 = w_sub06_result_dataout;
	assign w_sys_tmp3904 = (w_sys_tmp3905 + r_run_k_17);
	assign w_sys_tmp3905 = (r_run_copy0_j_89 * w_sys_tmp3902);
	assign w_sys_tmp3907 = (r_run_copy0_j_89 + w_sys_intOne);
	assign w_sys_tmp3908 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp3969 = 32'sh00000061;
	assign w_sys_tmp3970 = ( !w_sys_tmp3971 );
	assign w_sys_tmp3971 = (w_sys_tmp3972 < r_run_j_18);
	assign w_sys_tmp3972 = 32'sh00000080;
	assign w_sys_tmp3975 = (w_sys_tmp3976 + r_run_k_17);
	assign w_sys_tmp3976 = (r_run_j_18 * w_sys_tmp3977);
	assign w_sys_tmp3977 = 32'sh00000081;
	assign w_sys_tmp3978 = w_sub07_result_dataout;
	assign w_sys_tmp3979 = (w_sys_tmp3980 + r_run_k_17);
	assign w_sys_tmp3980 = (r_run_copy0_j_90 * w_sys_tmp3977);
	assign w_sys_tmp3982 = (r_run_copy0_j_90 + w_sys_intOne);
	assign w_sys_tmp3983 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp4044 = 32'sh00000041;
	assign w_sys_tmp4045 = ( !w_sys_tmp4046 );
	assign w_sys_tmp4046 = (w_sys_tmp4047 < r_run_k_17);
	assign w_sys_tmp4047 = 32'sh00000060;
	assign w_sys_tmp4048 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp4049 = 32'sh00000002;
	assign w_sys_tmp4050 = ( !w_sys_tmp4051 );
	assign w_sys_tmp4051 = (w_sys_tmp4052 < r_run_j_18);
	assign w_sys_tmp4052 = 32'sh00000020;
	assign w_sys_tmp4055 = (w_sys_tmp4056 + r_run_k_17);
	assign w_sys_tmp4056 = (r_run_j_18 * w_sys_tmp4057);
	assign w_sys_tmp4057 = 32'sh00000081;
	assign w_sys_tmp4058 = w_sub08_result_dataout;
	assign w_sys_tmp4059 = (w_sys_tmp4060 + r_run_k_17);
	assign w_sys_tmp4060 = (r_run_copy0_j_91 * w_sys_tmp4057);
	assign w_sys_tmp4062 = (r_run_copy0_j_91 + w_sys_intOne);
	assign w_sys_tmp4063 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp4124 = 32'sh00000021;
	assign w_sys_tmp4125 = ( !w_sys_tmp4126 );
	assign w_sys_tmp4126 = (w_sys_tmp4127 < r_run_j_18);
	assign w_sys_tmp4127 = 32'sh00000040;
	assign w_sys_tmp4130 = (w_sys_tmp4131 + r_run_k_17);
	assign w_sys_tmp4131 = (r_run_j_18 * w_sys_tmp4132);
	assign w_sys_tmp4132 = 32'sh00000081;
	assign w_sys_tmp4133 = w_sub09_result_dataout;
	assign w_sys_tmp4134 = (w_sys_tmp4135 + r_run_k_17);
	assign w_sys_tmp4135 = (r_run_copy0_j_92 * w_sys_tmp4132);
	assign w_sys_tmp4137 = (r_run_copy0_j_92 + w_sys_intOne);
	assign w_sys_tmp4138 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp4199 = 32'sh00000041;
	assign w_sys_tmp4200 = ( !w_sys_tmp4201 );
	assign w_sys_tmp4201 = (w_sys_tmp4202 < r_run_j_18);
	assign w_sys_tmp4202 = 32'sh00000060;
	assign w_sys_tmp4205 = (w_sys_tmp4206 + r_run_k_17);
	assign w_sys_tmp4206 = (r_run_j_18 * w_sys_tmp4207);
	assign w_sys_tmp4207 = 32'sh00000081;
	assign w_sys_tmp4208 = w_sub10_result_dataout;
	assign w_sys_tmp4209 = (w_sys_tmp4210 + r_run_k_17);
	assign w_sys_tmp4210 = (r_run_copy0_j_93 * w_sys_tmp4207);
	assign w_sys_tmp4212 = (r_run_copy0_j_93 + w_sys_intOne);
	assign w_sys_tmp4213 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp4274 = 32'sh00000061;
	assign w_sys_tmp4275 = ( !w_sys_tmp4276 );
	assign w_sys_tmp4276 = (w_sys_tmp4277 < r_run_j_18);
	assign w_sys_tmp4277 = 32'sh00000080;
	assign w_sys_tmp4280 = (w_sys_tmp4281 + r_run_k_17);
	assign w_sys_tmp4281 = (r_run_j_18 * w_sys_tmp4282);
	assign w_sys_tmp4282 = 32'sh00000081;
	assign w_sys_tmp4283 = w_sub11_result_dataout;
	assign w_sys_tmp4284 = (w_sys_tmp4285 + r_run_k_17);
	assign w_sys_tmp4285 = (r_run_copy0_j_94 * w_sys_tmp4282);
	assign w_sys_tmp4287 = (r_run_copy0_j_94 + w_sys_intOne);
	assign w_sys_tmp4288 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp4349 = 32'sh00000061;
	assign w_sys_tmp4350 = ( !w_sys_tmp4351 );
	assign w_sys_tmp4351 = (w_sys_tmp4352 < r_run_k_17);
	assign w_sys_tmp4352 = 32'sh00000080;
	assign w_sys_tmp4353 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp4354 = 32'sh00000002;
	assign w_sys_tmp4355 = ( !w_sys_tmp4356 );
	assign w_sys_tmp4356 = (w_sys_tmp4357 < r_run_j_18);
	assign w_sys_tmp4357 = 32'sh00000020;
	assign w_sys_tmp4360 = (w_sys_tmp4361 + r_run_k_17);
	assign w_sys_tmp4361 = (r_run_j_18 * w_sys_tmp4362);
	assign w_sys_tmp4362 = 32'sh00000081;
	assign w_sys_tmp4363 = w_sub12_result_dataout;
	assign w_sys_tmp4364 = (w_sys_tmp4365 + r_run_k_17);
	assign w_sys_tmp4365 = (r_run_copy0_j_95 * w_sys_tmp4362);
	assign w_sys_tmp4367 = (r_run_copy0_j_95 + w_sys_intOne);
	assign w_sys_tmp4368 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp4429 = 32'sh00000021;
	assign w_sys_tmp4430 = ( !w_sys_tmp4431 );
	assign w_sys_tmp4431 = (w_sys_tmp4432 < r_run_j_18);
	assign w_sys_tmp4432 = 32'sh00000040;
	assign w_sys_tmp4435 = (w_sys_tmp4436 + r_run_k_17);
	assign w_sys_tmp4436 = (r_run_j_18 * w_sys_tmp4437);
	assign w_sys_tmp4437 = 32'sh00000081;
	assign w_sys_tmp4438 = w_sub13_result_dataout;
	assign w_sys_tmp4439 = (w_sys_tmp4440 + r_run_k_17);
	assign w_sys_tmp4440 = (r_run_copy0_j_96 * w_sys_tmp4437);
	assign w_sys_tmp4442 = (r_run_copy0_j_96 + w_sys_intOne);
	assign w_sys_tmp4443 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp4504 = 32'sh00000041;
	assign w_sys_tmp4505 = ( !w_sys_tmp4506 );
	assign w_sys_tmp4506 = (w_sys_tmp4507 < r_run_j_18);
	assign w_sys_tmp4507 = 32'sh00000060;
	assign w_sys_tmp4510 = (w_sys_tmp4511 + r_run_k_17);
	assign w_sys_tmp4511 = (r_run_j_18 * w_sys_tmp4512);
	assign w_sys_tmp4512 = 32'sh00000081;
	assign w_sys_tmp4513 = w_sub14_result_dataout;
	assign w_sys_tmp4514 = (w_sys_tmp4515 + r_run_k_17);
	assign w_sys_tmp4515 = (r_run_copy0_j_97 * w_sys_tmp4512);
	assign w_sys_tmp4517 = (r_run_copy0_j_97 + w_sys_intOne);
	assign w_sys_tmp4518 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp4579 = 32'sh00000061;
	assign w_sys_tmp4580 = ( !w_sys_tmp4581 );
	assign w_sys_tmp4581 = (w_sys_tmp4582 < r_run_j_18);
	assign w_sys_tmp4582 = 32'sh00000080;
	assign w_sys_tmp4585 = (w_sys_tmp4586 + r_run_k_17);
	assign w_sys_tmp4586 = (r_run_j_18 * w_sys_tmp4587);
	assign w_sys_tmp4587 = 32'sh00000081;
	assign w_sys_tmp4588 = w_sub15_result_dataout;
	assign w_sys_tmp4589 = (w_sys_tmp4590 + r_run_k_17);
	assign w_sys_tmp4590 = (r_run_copy0_j_98 * w_sys_tmp4587);
	assign w_sys_tmp4592 = (r_run_copy0_j_98 + w_sys_intOne);
	assign w_sys_tmp4593 = (r_run_j_18 + w_sys_intOne);


	sub09
		sub09_inst(
			.i_fld_result_1_addr_0 (w_sub09_result_addr),
			.i_fld_result_1_datain_0 (w_sub09_result_datain),
			.o_fld_result_1_dataout_0 (w_sub09_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub09_result_r_w),
			.i_fld_u_0_addr_0 (w_sub09_u_addr),
			.i_fld_u_0_datain_0 (w_sub09_u_datain),
			.o_fld_u_0_dataout_0 (w_sub09_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub09_u_r_w),
			.o_run_busy (w_sub09_run_busy),
			.i_run_req (r_sub09_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub08
		sub08_inst(
			.i_fld_result_1_addr_0 (w_sub08_result_addr),
			.i_fld_result_1_datain_0 (w_sub08_result_datain),
			.o_fld_result_1_dataout_0 (w_sub08_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub08_result_r_w),
			.i_fld_u_0_addr_0 (w_sub08_u_addr),
			.i_fld_u_0_datain_0 (w_sub08_u_datain),
			.o_fld_u_0_dataout_0 (w_sub08_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub08_u_r_w),
			.o_run_busy (w_sub08_run_busy),
			.i_run_req (r_sub08_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub12
		sub12_inst(
			.i_fld_result_1_addr_0 (w_sub12_result_addr),
			.i_fld_result_1_datain_0 (w_sub12_result_datain),
			.o_fld_result_1_dataout_0 (w_sub12_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub12_result_r_w),
			.i_fld_u_0_addr_0 (w_sub12_u_addr),
			.i_fld_u_0_datain_0 (w_sub12_u_datain),
			.o_fld_u_0_dataout_0 (w_sub12_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub12_u_r_w),
			.o_run_busy (w_sub12_run_busy),
			.i_run_req (r_sub12_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub03
		sub03_inst(
			.i_fld_result_1_addr_0 (w_sub03_result_addr),
			.i_fld_result_1_datain_0 (w_sub03_result_datain),
			.o_fld_result_1_dataout_0 (w_sub03_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub03_result_r_w),
			.i_fld_u_0_addr_0 (w_sub03_u_addr),
			.i_fld_u_0_datain_0 (w_sub03_u_datain),
			.o_fld_u_0_dataout_0 (w_sub03_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub03_u_r_w),
			.o_run_busy (w_sub03_run_busy),
			.i_run_req (r_sub03_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub02
		sub02_inst(
			.i_fld_result_1_addr_0 (w_sub02_result_addr),
			.i_fld_result_1_datain_0 (w_sub02_result_datain),
			.o_fld_result_1_dataout_0 (w_sub02_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub02_result_r_w),
			.i_fld_u_0_addr_0 (w_sub02_u_addr),
			.i_fld_u_0_datain_0 (w_sub02_u_datain),
			.o_fld_u_0_dataout_0 (w_sub02_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub02_u_r_w),
			.o_run_busy (w_sub02_run_busy),
			.i_run_req (r_sub02_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub11
		sub11_inst(
			.i_fld_result_1_addr_0 (w_sub11_result_addr),
			.i_fld_result_1_datain_0 (w_sub11_result_datain),
			.o_fld_result_1_dataout_0 (w_sub11_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub11_result_r_w),
			.i_fld_u_0_addr_0 (w_sub11_u_addr),
			.i_fld_u_0_datain_0 (w_sub11_u_datain),
			.o_fld_u_0_dataout_0 (w_sub11_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub11_u_r_w),
			.o_run_busy (w_sub11_run_busy),
			.i_run_req (r_sub11_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub14
		sub14_inst(
			.i_fld_result_1_addr_0 (w_sub14_result_addr),
			.i_fld_result_1_datain_0 (w_sub14_result_datain),
			.o_fld_result_1_dataout_0 (w_sub14_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub14_result_r_w),
			.i_fld_u_0_addr_0 (w_sub14_u_addr),
			.i_fld_u_0_datain_0 (w_sub14_u_datain),
			.o_fld_u_0_dataout_0 (w_sub14_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub14_u_r_w),
			.o_run_busy (w_sub14_run_busy),
			.i_run_req (r_sub14_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub01
		sub01_inst(
			.i_fld_result_1_addr_0 (w_sub01_result_addr),
			.i_fld_result_1_datain_0 (w_sub01_result_datain),
			.o_fld_result_1_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub01_result_r_w),
			.i_fld_u_0_addr_0 (w_sub01_u_addr),
			.i_fld_u_0_datain_0 (w_sub01_u_datain),
			.o_fld_u_0_dataout_0 (w_sub01_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub01_u_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub13
		sub13_inst(
			.i_fld_result_1_addr_0 (w_sub13_result_addr),
			.i_fld_result_1_datain_0 (w_sub13_result_datain),
			.o_fld_result_1_dataout_0 (w_sub13_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub13_result_r_w),
			.i_fld_u_0_addr_0 (w_sub13_u_addr),
			.i_fld_u_0_datain_0 (w_sub13_u_datain),
			.o_fld_u_0_dataout_0 (w_sub13_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub13_u_r_w),
			.o_run_busy (w_sub13_run_busy),
			.i_run_req (r_sub13_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub00
		sub00_inst(
			.i_fld_result_1_addr_0 (w_sub00_result_addr),
			.i_fld_result_1_datain_0 (w_sub00_result_datain),
			.o_fld_result_1_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub00_result_r_w),
			.i_fld_u_0_addr_0 (w_sub00_u_addr),
			.i_fld_u_0_datain_0 (w_sub00_u_datain),
			.o_fld_u_0_dataout_0 (w_sub00_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub00_u_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub07
		sub07_inst(
			.i_fld_result_1_addr_0 (w_sub07_result_addr),
			.i_fld_result_1_datain_0 (w_sub07_result_datain),
			.o_fld_result_1_dataout_0 (w_sub07_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub07_result_r_w),
			.i_fld_u_0_addr_0 (w_sub07_u_addr),
			.i_fld_u_0_datain_0 (w_sub07_u_datain),
			.o_fld_u_0_dataout_0 (w_sub07_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub07_u_r_w),
			.o_run_busy (w_sub07_run_busy),
			.i_run_req (r_sub07_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub06
		sub06_inst(
			.i_fld_result_1_addr_0 (w_sub06_result_addr),
			.i_fld_result_1_datain_0 (w_sub06_result_datain),
			.o_fld_result_1_dataout_0 (w_sub06_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub06_result_r_w),
			.i_fld_u_0_addr_0 (w_sub06_u_addr),
			.i_fld_u_0_datain_0 (w_sub06_u_datain),
			.o_fld_u_0_dataout_0 (w_sub06_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub06_u_r_w),
			.o_run_busy (w_sub06_run_busy),
			.i_run_req (r_sub06_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub15
		sub15_inst(
			.i_fld_result_1_addr_0 (w_sub15_result_addr),
			.i_fld_result_1_datain_0 (w_sub15_result_datain),
			.o_fld_result_1_dataout_0 (w_sub15_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub15_result_r_w),
			.i_fld_u_0_addr_0 (w_sub15_u_addr),
			.i_fld_u_0_datain_0 (w_sub15_u_datain),
			.o_fld_u_0_dataout_0 (w_sub15_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub15_u_r_w),
			.o_run_busy (w_sub15_run_busy),
			.i_run_req (r_sub15_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub05
		sub05_inst(
			.i_fld_result_1_addr_0 (w_sub05_result_addr),
			.i_fld_result_1_datain_0 (w_sub05_result_datain),
			.o_fld_result_1_dataout_0 (w_sub05_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub05_result_r_w),
			.i_fld_u_0_addr_0 (w_sub05_u_addr),
			.i_fld_u_0_datain_0 (w_sub05_u_datain),
			.o_fld_u_0_dataout_0 (w_sub05_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub05_u_r_w),
			.o_run_busy (w_sub05_run_busy),
			.i_run_req (r_sub05_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub04
		sub04_inst(
			.i_fld_result_1_addr_0 (w_sub04_result_addr),
			.i_fld_result_1_datain_0 (w_sub04_result_datain),
			.o_fld_result_1_dataout_0 (w_sub04_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub04_result_r_w),
			.i_fld_u_0_addr_0 (w_sub04_u_addr),
			.i_fld_u_0_datain_0 (w_sub04_u_datain),
			.o_fld_u_0_dataout_0 (w_sub04_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub04_u_r_w),
			.o_run_busy (w_sub04_run_busy),
			.i_run_req (r_sub04_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub10
		sub10_inst(
			.i_fld_result_1_addr_0 (w_sub10_result_addr),
			.i_fld_result_1_datain_0 (w_sub10_result_datain),
			.o_fld_result_1_dataout_0 (w_sub10_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub10_result_r_w),
			.i_fld_u_0_addr_0 (w_sub10_u_addr),
			.i_fld_u_0_datain_0 (w_sub10_u_datain),
			.o_fld_u_0_dataout_0 (w_sub10_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub10_u_r_w),
			.o_run_busy (w_sub10_run_busy),
			.i_run_req (r_sub10_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_u_0(
			.clk (clock),
			.ce_0 (w_fld_u_0_ce_0),
			.addr_0 (w_fld_u_0_addr_0),
			.datain_0 (w_fld_u_0_datain_0),
			.dataout_0 (w_fld_u_0_dataout_0),
			.r_w_0 (w_fld_u_0_r_w_0),
			.ce_1 (w_fld_u_0_ce_1),
			.addr_1 (r_fld_u_0_addr_1),
			.datain_1 (r_fld_u_0_datain_1),
			.dataout_1 (w_fld_u_0_dataout_1),
			.r_w_1 (r_fld_u_0_r_w_1)
		);

	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						9'h12f: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 9'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h0: begin
							r_sys_run_phase <= 9'h2;
						end

						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h4;

									end
								end

							endcase
						end

						9'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h5;

									end
								end

							endcase
						end

						9'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4) ? 9'h9 : 9'hf);

									end
								end

							endcase
						end

						9'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h5;

									end
								end

							endcase
						end

						9'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'ha;

									end
								end

							endcase
						end

						9'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7) ? 9'hd : 9'h6);

									end
								end

							endcase
						end

						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sys_run_phase <= 9'ha;

									end
								end

							endcase
						end

						9'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h10;

									end
								end

							endcase
						end

						9'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp52) ? 9'h14 : 9'h2c);

									end
								end

							endcase
						end

						9'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h10;

									end
								end

							endcase
						end

						9'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h15;

									end
								end

							endcase
						end

						9'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp56) ? 9'h18 : 9'h1a);

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h15;

									end
								end

							endcase
						end

						9'h1a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h1b;

									end
								end

							endcase
						end

						9'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp131) ? 9'h1e : 9'h20);

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h1b;

									end
								end

							endcase
						end

						9'h20: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h21;

									end
								end

							endcase
						end

						9'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp206) ? 9'h24 : 9'h26);

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h21;

									end
								end

							endcase
						end

						9'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h27;

									end
								end

							endcase
						end

						9'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp281) ? 9'h2a : 9'h11);

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h27;

									end
								end

							endcase
						end

						9'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h2d;

									end
								end

							endcase
						end

						9'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp356) ? 9'h31 : 9'h49);

									end
								end

							endcase
						end

						9'h2e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h2d;

									end
								end

							endcase
						end

						9'h31: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h32;

									end
								end

							endcase
						end

						9'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp360) ? 9'h35 : 9'h37);

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h32;

									end
								end

							endcase
						end

						9'h37: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h38;

									end
								end

							endcase
						end

						9'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp435) ? 9'h3b : 9'h3d);

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h38;

									end
								end

							endcase
						end

						9'h3d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h3e;

									end
								end

							endcase
						end

						9'h3e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp510) ? 9'h41 : 9'h43);

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h3e;

									end
								end

							endcase
						end

						9'h43: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h44;

									end
								end

							endcase
						end

						9'h44: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp585) ? 9'h47 : 9'h2e);

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h44;

									end
								end

							endcase
						end

						9'h49: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h4a;

									end
								end

							endcase
						end

						9'h4a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp660) ? 9'h4e : 9'h66);

									end
								end

							endcase
						end

						9'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h4a;

									end
								end

							endcase
						end

						9'h4e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h4f;

									end
								end

							endcase
						end

						9'h4f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp664) ? 9'h52 : 9'h54);

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h4f;

									end
								end

							endcase
						end

						9'h54: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h55;

									end
								end

							endcase
						end

						9'h55: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp739) ? 9'h58 : 9'h5a);

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h55;

									end
								end

							endcase
						end

						9'h5a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h5b;

									end
								end

							endcase
						end

						9'h5b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp814) ? 9'h5e : 9'h60);

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h5b;

									end
								end

							endcase
						end

						9'h60: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h61;

									end
								end

							endcase
						end

						9'h61: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp889) ? 9'h64 : 9'h4b);

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h61;

									end
								end

							endcase
						end

						9'h66: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h67;

									end
								end

							endcase
						end

						9'h67: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp964) ? 9'h6b : 9'h83);

									end
								end

							endcase
						end

						9'h68: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h67;

									end
								end

							endcase
						end

						9'h6b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h6c;

									end
								end

							endcase
						end

						9'h6c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp968) ? 9'h6f : 9'h71);

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h6c;

									end
								end

							endcase
						end

						9'h71: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h72;

									end
								end

							endcase
						end

						9'h72: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1043) ? 9'h75 : 9'h77);

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h72;

									end
								end

							endcase
						end

						9'h77: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h78;

									end
								end

							endcase
						end

						9'h78: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1118) ? 9'h7b : 9'h7d);

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h78;

									end
								end

							endcase
						end

						9'h7d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h7e;

									end
								end

							endcase
						end

						9'h7e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1193) ? 9'h81 : 9'h68);

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h7e;

									end
								end

							endcase
						end

						9'h83: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h84;

									end
								end

							endcase
						end

						9'h84: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1267) ? 9'h87 : 9'hbb);

									end
								end

							endcase
						end

						9'h85: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h84;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h10: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_phase <= 9'h89;

									end
								end

							endcase
						end

						9'h89: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_phase <= 9'h8b;

									end
								end

							endcase
						end

						9'h8b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h8c;

									end
								end

							endcase
						end

						9'h8c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1271) ? 9'h8f : 9'h91);

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_phase <= 9'h8c;

									end
								end

							endcase
						end

						9'h91: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h92;

									end
								end

							endcase
						end

						9'h92: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1311) ? 9'h95 : 9'h97);

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_phase <= 9'h92;

									end
								end

							endcase
						end

						9'h97: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h98;

									end
								end

							endcase
						end

						9'h98: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1351) ? 9'h9b : 9'h9d);

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_phase <= 9'h98;

									end
								end

							endcase
						end

						9'h9d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h9e;

									end
								end

							endcase
						end

						9'h9e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1391) ? 9'ha1 : 9'ha3);

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_phase <= 9'h9e;

									end
								end

							endcase
						end

						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'ha4;

									end
								end

							endcase
						end

						9'ha4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1431) ? 9'ha7 : 9'ha9);

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 9'ha4;

									end
								end

							endcase
						end

						9'ha9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'haa;

									end
								end

							endcase
						end

						9'haa: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1932) ? 9'had : 9'haf);

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 9'haa;

									end
								end

							endcase
						end

						9'haf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hb0;

									end
								end

							endcase
						end

						9'hb0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2433) ? 9'hb3 : 9'hb5);

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 9'hb0;

									end
								end

							endcase
						end

						9'hb5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hb6;

									end
								end

							endcase
						end

						9'hb6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2934) ? 9'hb9 : 9'h85);

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 9'hb6;

									end
								end

							endcase
						end

						9'hbb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hbc;

									end
								end

							endcase
						end

						9'hbc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3435) ? 9'hc0 : 9'hd8);

									end
								end

							endcase
						end

						9'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hbc;

									end
								end

							endcase
						end

						9'hc0: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hc1;

									end
								end

							endcase
						end

						9'hc1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3440) ? 9'hc4 : 9'hc6);

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'hc1;

									end
								end

							endcase
						end

						9'hc6: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hc7;

									end
								end

							endcase
						end

						9'hc7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3515) ? 9'hca : 9'hcc);

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'hc7;

									end
								end

							endcase
						end

						9'hcc: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hcd;

									end
								end

							endcase
						end

						9'hcd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3590) ? 9'hd0 : 9'hd2);

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'hcd;

									end
								end

							endcase
						end

						9'hd2: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hd3;

									end
								end

							endcase
						end

						9'hd3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3665) ? 9'hd6 : 9'hbd);

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'hd3;

									end
								end

							endcase
						end

						9'hd8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hd9;

									end
								end

							endcase
						end

						9'hd9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3740) ? 9'hdd : 9'hf5);

									end
								end

							endcase
						end

						9'hda: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hd9;

									end
								end

							endcase
						end

						9'hdd: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hde;

									end
								end

							endcase
						end

						9'hde: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3745) ? 9'he1 : 9'he3);

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'hde;

									end
								end

							endcase
						end

						9'he3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'he4;

									end
								end

							endcase
						end

						9'he4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3820) ? 9'he7 : 9'he9);

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'he4;

									end
								end

							endcase
						end

						9'he9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hea;

									end
								end

							endcase
						end

						9'hea: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3895) ? 9'hed : 9'hef);

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'hea;

									end
								end

							endcase
						end

						9'hef: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hf0;

									end
								end

							endcase
						end

						9'hf0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3970) ? 9'hf3 : 9'hda);

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'hf0;

									end
								end

							endcase
						end

						9'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hf6;

									end
								end

							endcase
						end

						9'hf6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4045) ? 9'hfa : 9'h112);

									end
								end

							endcase
						end

						9'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hf6;

									end
								end

							endcase
						end

						9'hfa: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hfb;

									end
								end

							endcase
						end

						9'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4050) ? 9'hfe : 9'h100);

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'hfb;

									end
								end

							endcase
						end

						9'h100: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h101;

									end
								end

							endcase
						end

						9'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4125) ? 9'h104 : 9'h106);

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h101;

									end
								end

							endcase
						end

						9'h106: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h107;

									end
								end

							endcase
						end

						9'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4200) ? 9'h10a : 9'h10c);

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h107;

									end
								end

							endcase
						end

						9'h10c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h10d;

									end
								end

							endcase
						end

						9'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4275) ? 9'h110 : 9'hf7);

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h10d;

									end
								end

							endcase
						end

						9'h112: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h113;

									end
								end

							endcase
						end

						9'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4350) ? 9'h117 : 9'h12f);

									end
								end

							endcase
						end

						9'h114: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h113;

									end
								end

							endcase
						end

						9'h117: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h118;

									end
								end

							endcase
						end

						9'h118: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4355) ? 9'h11b : 9'h11d);

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h118;

									end
								end

							endcase
						end

						9'h11d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h11e;

									end
								end

							endcase
						end

						9'h11e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4430) ? 9'h121 : 9'h123);

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h11e;

									end
								end

							endcase
						end

						9'h123: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h124;

									end
								end

							endcase
						end

						9'h124: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4505) ? 9'h127 : 9'h129);

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h124;

									end
								end

							endcase
						end

						9'h129: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h12a;

									end
								end

							endcase
						end

						9'h12a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4580) ? 9'h12d : 9'h114);

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h12a;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sys_run_phase <= 9'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 5'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h2e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h31: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h37: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h3e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h43: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h44: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h49: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h4a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h4e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h4f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h54: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h55: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h5a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h5b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h60: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h61: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h66: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h67: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h68: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h6c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h72: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h78: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h7d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h7e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h83: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h84: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h85: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h89: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h8b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h8c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h91: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h92: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h97: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h98: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h9d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h9e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'haa: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'haf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hb0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hb5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hb6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hbb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hbc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hc0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hc1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hc6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hc7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hcc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hcd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hda: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hdd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hde: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'he3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'he4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'he9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hea: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hfa: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h100: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h106: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h10c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h112: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h114: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h117: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h118: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h11d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h11e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h123: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h124: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h129: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h12a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 6'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h5)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h2e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h31: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h37: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h3e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h43: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h44: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h49: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h4a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h4e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h4f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h54: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h55: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h5a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h5b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h60: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h61: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h66: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h67: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h68: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h6c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h72: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h78: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h7d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h7e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h83: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h84: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h85: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h89: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub00_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub01_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub02_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub03_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub04_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub05_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub06_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub07_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub08_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub09_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub10_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub11_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub12_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub13_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub14_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub15_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h8b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h8c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'hc)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h91: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h92: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'hc)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h97: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h98: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'hc)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h9d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h9e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'hc)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'ha3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'ha4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'ha9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'haa: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'haf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hb0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hb5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hb6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hbb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hbc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hc0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hc1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hc6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hc7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hcc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hcd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hd2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hd3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hd8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hd9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hda: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hdd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hde: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'he3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'he4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'he9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hea: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hf0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hf6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hfa: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h100: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h106: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h10c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h112: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h114: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h117: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h118: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h11d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h11e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h123: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h124: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h129: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h12a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						9'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						9'h12f: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp11[14:0] );

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp65[14:0] );

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp140[14:0] );

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp215[14:0] );

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp290[14:0] );

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp369[14:0] );

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp444[14:0] );

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp519[14:0] );

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp594[14:0] );

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp673[14:0] );

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp748[14:0] );

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp823[14:0] );

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp898[14:0] );

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp977[14:0] );

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1052[14:0] );

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1127[14:0] );

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1202[14:0] );

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3445[14:0] );

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3520[14:0] );

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3595[14:0] );

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3670[14:0] );

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3750[14:0] );

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3825[14:0] );

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3900[14:0] );

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3975[14:0] );

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4055[14:0] );

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4130[14:0] );

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4205[14:0] );

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4280[14:0] );

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4360[14:0] );

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4435[14:0] );

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4510[14:0] );

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4585[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp14;

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp3448;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp3523;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp3598;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp3673;

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp3753;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp3828;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp3903;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp3978;

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp4058;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp4133;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp4208;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp4283;

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp4363;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp4438;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp4513;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp4588;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h12f: begin
							r_fld_u_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_17 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_17 <= w_sys_tmp6;

									end
								end

							endcase
						end

						9'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_17 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_17 <= w_sys_tmp55;

									end
								end

							endcase
						end

						9'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_17 <= w_sys_tmp355;

									end
								end

							endcase
						end

						9'h2e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_17 <= w_sys_tmp359;

									end
								end

							endcase
						end

						9'h49: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_17 <= w_sys_tmp659;

									end
								end

							endcase
						end

						9'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_17 <= w_sys_tmp663;

									end
								end

							endcase
						end

						9'h66: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_17 <= w_sys_tmp963;

									end
								end

							endcase
						end

						9'h68: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_17 <= w_sys_tmp967;

									end
								end

							endcase
						end

						9'h8b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_17 <= w_sys_tmp1270;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_run_k_17 <= w_sys_tmp1309;

									end
								end

							endcase
						end

						9'h91: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_17 <= w_sys_tmp1310;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_run_k_17 <= w_sys_tmp1349;

									end
								end

							endcase
						end

						9'h97: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_17 <= w_sys_tmp1350;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_run_k_17 <= w_sys_tmp1389;

									end
								end

							endcase
						end

						9'h9d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_17 <= w_sys_tmp1390;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_run_k_17 <= w_sys_tmp1429;

									end
								end

							endcase
						end

						9'hbb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_17 <= w_sys_tmp3434;

									end
								end

							endcase
						end

						9'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_17 <= w_sys_tmp3438;

									end
								end

							endcase
						end

						9'hd8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_17 <= w_sys_tmp3739;

									end
								end

							endcase
						end

						9'hda: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_17 <= w_sys_tmp3743;

									end
								end

							endcase
						end

						9'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_17 <= w_sys_tmp4044;

									end
								end

							endcase
						end

						9'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_17 <= w_sys_tmp4048;

									end
								end

							endcase
						end

						9'h112: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_17 <= w_sys_tmp4349;

									end
								end

							endcase
						end

						9'h114: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_17 <= w_sys_tmp4353;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_18 <= w_sys_tmp15;

									end
								end

							endcase
						end

						9'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp69;

									end
								end

							endcase
						end

						9'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp130;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp144;

									end
								end

							endcase
						end

						9'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp205;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp219;

									end
								end

							endcase
						end

						9'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp280;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp294;

									end
								end

							endcase
						end

						9'h31: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp373;

									end
								end

							endcase
						end

						9'h37: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp434;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp448;

									end
								end

							endcase
						end

						9'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp509;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp523;

									end
								end

							endcase
						end

						9'h43: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp584;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp598;

									end
								end

							endcase
						end

						9'h4e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp677;

									end
								end

							endcase
						end

						9'h54: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp738;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp752;

									end
								end

							endcase
						end

						9'h5a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp813;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp827;

									end
								end

							endcase
						end

						9'h60: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp888;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp902;

									end
								end

							endcase
						end

						9'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp981;

									end
								end

							endcase
						end

						9'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp1042;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp1056;

									end
								end

							endcase
						end

						9'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp1117;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp1131;

									end
								end

							endcase
						end

						9'h7d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp1192;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp1206;

									end
								end

							endcase
						end

						9'ha3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp1430;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_18 <= w_sys_tmp1504;

									end
								end

							endcase
						end

						9'ha9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp1931;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_18 <= w_sys_tmp2005;

									end
								end

							endcase
						end

						9'haf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp2432;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_18 <= w_sys_tmp2506;

									end
								end

							endcase
						end

						9'hb5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp2933;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_18 <= w_sys_tmp3007;

									end
								end

							endcase
						end

						9'hc0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp3439;

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp3453;

									end
								end

							endcase
						end

						9'hc6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp3514;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp3528;

									end
								end

							endcase
						end

						9'hcc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp3589;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp3603;

									end
								end

							endcase
						end

						9'hd2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp3664;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp3678;

									end
								end

							endcase
						end

						9'hdd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp3744;

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp3758;

									end
								end

							endcase
						end

						9'he3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp3819;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp3833;

									end
								end

							endcase
						end

						9'he9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp3894;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp3908;

									end
								end

							endcase
						end

						9'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp3969;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp3983;

									end
								end

							endcase
						end

						9'hfa: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp4049;

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp4063;

									end
								end

							endcase
						end

						9'h100: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp4124;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp4138;

									end
								end

							endcase
						end

						9'h106: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp4199;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp4213;

									end
								end

							endcase
						end

						9'h10c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp4274;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp4288;

									end
								end

							endcase
						end

						9'h117: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp4354;

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp4368;

									end
								end

							endcase
						end

						9'h11d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp4429;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp4443;

									end
								end

							endcase
						end

						9'h123: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp4504;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp4518;

									end
								end

							endcase
						end

						9'h129: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_18 <= w_sys_tmp4579;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_18 <= w_sys_tmp4593;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h83: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_n_19 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h85: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_n_19 <= w_sys_tmp1269;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_mx_20 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_my_21 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_nlast_22 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_23 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_23 <= w_sys_tmp68;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_24 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_24 <= w_sys_tmp143;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h20: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_25 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_25 <= w_sys_tmp218;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_26 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_26 <= w_sys_tmp293;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h31: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_27 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_27 <= w_sys_tmp372;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h37: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_28 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_28 <= w_sys_tmp447;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_29 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_29 <= w_sys_tmp522;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h43: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_30 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_30 <= w_sys_tmp597;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h4e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_31 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_31 <= w_sys_tmp676;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h54: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_32 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_32 <= w_sys_tmp751;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_33 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_33 <= w_sys_tmp826;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h60: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_34 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_34 <= w_sys_tmp901;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_35 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_35 <= w_sys_tmp980;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h71: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_36 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_36 <= w_sys_tmp1055;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h77: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_37 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_37 <= w_sys_tmp1130;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_38 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_38 <= w_sys_tmp1205;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_39 <= r_run_j_18;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_39 <= w_sys_tmp1493;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_40 <= r_run_j_18;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_40 <= w_sys_tmp1494;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_41 <= r_run_j_18;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_41 <= w_sys_tmp1495;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_42 <= r_run_j_18;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_42 <= w_sys_tmp1496;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_43 <= r_run_j_18;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_43 <= w_sys_tmp1497;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_44 <= r_run_j_18;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_44 <= w_sys_tmp1498;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_45 <= r_run_j_18;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_45 <= w_sys_tmp1499;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_46 <= r_run_j_18;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_46 <= w_sys_tmp1500;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_47 <= r_run_j_18;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_47 <= w_sys_tmp1501;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_48 <= r_run_j_18;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_48 <= w_sys_tmp1502;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_49 <= r_run_j_18;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_49 <= w_sys_tmp1503;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_50 <= r_run_j_18;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_50 <= w_sys_tmp1994;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_51 <= r_run_j_18;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_51 <= w_sys_tmp1995;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_52 <= r_run_j_18;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_52 <= w_sys_tmp1996;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_53 <= r_run_j_18;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_53 <= w_sys_tmp1997;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_54 <= r_run_j_18;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_54 <= w_sys_tmp1998;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_55 <= r_run_j_18;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_55 <= w_sys_tmp1999;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_56 <= r_run_j_18;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_56 <= w_sys_tmp2000;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_57 <= r_run_j_18;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_57 <= w_sys_tmp2001;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_58 <= r_run_j_18;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_58 <= w_sys_tmp2002;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_59 <= r_run_j_18;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_59 <= w_sys_tmp2003;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_60 <= r_run_j_18;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_60 <= w_sys_tmp2004;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'haf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_61 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_61 <= w_sys_tmp2495;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'haf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_62 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_62 <= w_sys_tmp2496;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'haf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_63 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_63 <= w_sys_tmp2497;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'haf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_64 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_64 <= w_sys_tmp2498;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'haf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_65 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_65 <= w_sys_tmp2499;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'haf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_66 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_66 <= w_sys_tmp2500;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'haf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_67 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_67 <= w_sys_tmp2501;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'haf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_68 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_68 <= w_sys_tmp2502;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'haf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_69 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_69 <= w_sys_tmp2503;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'haf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_70 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_70 <= w_sys_tmp2504;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'haf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_71 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_71 <= w_sys_tmp2505;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hb5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_72 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_72 <= w_sys_tmp2996;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hb5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_73 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_73 <= w_sys_tmp2997;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hb5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_74 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_74 <= w_sys_tmp2998;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hb5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_75 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_75 <= w_sys_tmp2999;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hb5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_76 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_76 <= w_sys_tmp3000;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hb5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_77 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_77 <= w_sys_tmp3001;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hb5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_78 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_78 <= w_sys_tmp3002;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hb5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_79 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_79 <= w_sys_tmp3003;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hb5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_80 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_80 <= w_sys_tmp3004;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hb5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_81 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_81 <= w_sys_tmp3005;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hb5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_82 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_82 <= w_sys_tmp3006;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hc0: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_83 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_83 <= w_sys_tmp3452;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hc6: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_84 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_84 <= w_sys_tmp3527;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hcc: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_85 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_85 <= w_sys_tmp3602;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd2: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_86 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_86 <= w_sys_tmp3677;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hdd: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_87 <= r_run_j_18;

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_87 <= w_sys_tmp3757;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'he3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_88 <= r_run_j_18;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_88 <= w_sys_tmp3832;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'he9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_89 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_89 <= w_sys_tmp3907;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hef: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_90 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_90 <= w_sys_tmp3982;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hfa: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_91 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_91 <= w_sys_tmp4062;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h100: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_92 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_92 <= w_sys_tmp4137;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h106: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_93 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_93 <= w_sys_tmp4212;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h10c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_94 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_94 <= w_sys_tmp4287;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h117: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_95 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_95 <= w_sys_tmp4367;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h11d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_96 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_96 <= w_sys_tmp4442;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h123: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_97 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_97 <= w_sys_tmp4517;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h129: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_98 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_98 <= w_sys_tmp4592;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub09_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub09_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp744[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_u_datain <= w_sys_tmp747;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub09_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp1328[12:0] );

									end
									else
									if((r_sys_run_step==6'hb)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp1344[12:0] );

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp1339[12:0] );

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp1333[12:0] );

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp2448[12:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp2443[12:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp2458[12:0] );

									end
									else
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp2472[12:0] );

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4134[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9)) begin
										r_sub09_result_datain <= w_sys_tmp1318;

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_sub09_result_datain <= r_sys_tmp1_float;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub09_result_datain <= w_sys_tmp2452;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub09_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub09_result_datain <= w_sys_tmp2490;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha)) begin
										r_sub09_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub09_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub09_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub08_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub08_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp669[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_u_datain <= w_sys_tmp672;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub08_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1299[12:0] );

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1293[12:0] );

									end
									else
									if((r_sys_run_step==6'hb)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1304[12:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1288[12:0] );

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp2438[12:0] );

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp2453[12:0] );

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4059[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha)) begin
										r_sub08_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_sub08_result_datain <= w_sys_tmp1278;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub08_result_datain <= w_sys_tmp2442;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha)) begin
										r_sub08_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub08_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub08_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h10: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub12_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub12_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp973[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_u_datain <= w_sys_tmp976;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub12_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp1299[12:0] );

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp1304[12:0] );

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp2939[12:0] );

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp2954[12:0] );

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp4364[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub12_result_datain <= w_sys_tmp1306;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub12_result_datain <= w_sys_tmp2943;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_sub12_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub12_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub12_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp286[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_u_datain <= w_sys_tmp289;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub03_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1396[12:0] );

									end
									else
									if((r_sys_run_step==6'h3)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1402[12:0] );

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1479[12:0] );

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1484[12:0] );

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp3674[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub03_result_datain <= w_sys_tmp1398;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub03_result_datain <= w_sys_tmp1488;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub03_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub03_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub03_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h2: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp211[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_u_datain <= w_sys_tmp214;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub02_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1356[12:0] );

									end
									else
									if((r_sys_run_step==6'h3)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1362[12:0] );

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1460[12:0] );

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1475[12:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1465[12:0] );

									end
									else
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1489[12:0] );

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3599[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub02_result_datain <= w_sys_tmp1358;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub02_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub02_result_datain <= w_sys_tmp1440;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub02_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub02_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub02_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h9: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub11_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub11_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp894[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_u_datain <= w_sys_tmp897;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub11_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp1413[12:0] );

									end
									else
									if((r_sys_run_step==6'hb)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp1424[12:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp1408[12:0] );

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp1419[12:0] );

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp2481[12:0] );

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp2486[12:0] );

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp4284[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha)) begin
										r_sub11_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_sub11_result_datain <= w_sys_tmp1398;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub11_result_datain <= w_sys_tmp2490;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha)) begin
										r_sub11_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub11_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub11_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'hb: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub14_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub14_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp1123[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_u_datain <= w_sys_tmp1126;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub14_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp1379[12:0] );

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp1384[12:0] );

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp2992[12:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp2963[12:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp2968[12:0] );

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp2978[12:0] );

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp4514[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub14_result_datain <= w_sys_tmp1386;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub14_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub14_result_datain <= w_sys_tmp2943;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_sub14_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub14_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub14_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp136[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_u_datain <= w_sys_tmp139;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub01_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1316[12:0] );

									end
									else
									if((r_sys_run_step==6'h3)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1322[12:0] );

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1456[12:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1441[12:0] );

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1446[12:0] );

									end
									else
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1470[12:0] );

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3524[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub01_result_datain <= w_sys_tmp1318;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub01_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub01_result_datain <= w_sys_tmp1488;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub01_result_datain <= w_sys_tmp1450;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub01_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub01_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'ha: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub13_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub13_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp1048[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_u_datain <= w_sys_tmp1051;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub13_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp1344[12:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp1339[12:0] );

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp2973[12:0] );

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp2949[12:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp2944[12:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp2959[12:0] );

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp4439[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub13_result_datain <= w_sys_tmp1346;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub13_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub13_result_datain <= w_sys_tmp2991;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub13_result_datain <= w_sys_tmp2953;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_sub13_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub13_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub13_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp61[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_u_datain <= w_sys_tmp64;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub00_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1282[12:0] );

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1276[12:0] );

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1451[12:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1436[12:0] );

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3449[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub00_result_datain <= w_sys_tmp1278;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub00_result_datain <= w_sys_tmp1440;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub00_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub00_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub07_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub07_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp590[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_u_datain <= w_sys_tmp593;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub07_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1413[12:0] );

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1408[12:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1396[12:0] );

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1402[12:0] );

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1985[12:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1980[12:0] );

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp3979[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub07_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub07_result_datain <= w_sys_tmp1404;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub07_result_datain <= w_sys_tmp1989;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6)) begin
										r_sub07_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub07_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub07_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub06_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub06_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp515[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_u_datain <= w_sys_tmp518;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub06_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1356[12:0] );

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1368[12:0] );

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1362[12:0] );

									end
									else
									if((r_sys_run_step==6'h7)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1373[12:0] );

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1976[12:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1966[12:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1961[12:0] );

									end
									else
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1990[12:0] );

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp3904[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub06_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub06_result_datain <= w_sys_tmp1364;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub06_result_datain <= w_sys_tmp1941;

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub06_result_datain <= r_sys_tmp1_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6)) begin
										r_sub06_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub06_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub06_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub15_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub15_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp1198[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_u_datain <= w_sys_tmp1201;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub15_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp1424[12:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp1419[12:0] );

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp2987[12:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp2982[12:0] );

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp4589[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub15_result_datain <= w_sys_tmp1426;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub15_result_datain <= w_sys_tmp2991;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_sub15_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub15_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub15_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub05_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub05_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp440[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_u_datain <= w_sys_tmp443;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub05_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1328[12:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1316[12:0] );

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1322[12:0] );

									end
									else
									if((r_sys_run_step==6'h7)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1333[12:0] );

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1957[12:0] );

									end
									else
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1971[12:0] );

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1947[12:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1942[12:0] );

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp3829[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub05_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub05_result_datain <= w_sys_tmp1324;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub05_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub05_result_datain <= w_sys_tmp1951;

									end
									else
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub05_result_datain <= w_sys_tmp1989;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6)) begin
										r_sub05_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub05_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub05_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'he: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub04_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub04_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp365[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_u_datain <= w_sys_tmp368;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub04_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1293[12:0] );

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1288[12:0] );

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1282[12:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1276[12:0] );

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1952[12:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1937[12:0] );

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp3754[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5)) begin
										r_sub04_result_datain <= w_sys_tmp1284;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub04_result_datain <= r_sys_tmp0_float;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub04_result_datain <= w_sys_tmp1941;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6)) begin
										r_sub04_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub04_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub04_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub10_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub10_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp819[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_u_datain <= w_sys_tmp822;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub10_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp1379[12:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp1368[12:0] );

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp1373[12:0] );

									end
									else
									if((r_sys_run_step==6'hb)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp1384[12:0] );

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp2491[12:0] );

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp2477[12:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp2467[12:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp2462[12:0] );

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp4209[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9)) begin
										r_sub10_result_datain <= w_sys_tmp1358;

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_sub10_result_datain <= r_sys_tmp1_float;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub10_result_datain <= w_sys_tmp2442;

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub10_result_datain <= r_sys_tmp1_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha)) begin
										r_sub10_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub10_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub10_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp1_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp1_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp1_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp1_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
