/*
TimeStamp:	2017/1/5		15:47
*/


module ThreadTop(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_threadTopMain_req,	
	output                o_threadTopMain_busy,	
	output signed  [31:0] o_threadTopMain_return,	
	input  signed  [ 4:0] i_subB_arrayB_addr,	
	input  signed  [31:0] i_subB_arrayB_datain,	
	output signed  [31:0] o_subB_arrayB_dataout,	
	input                 i_subB_arrayB_r_w,	
	output signed  [31:0] o_subB_ret,	
	input  signed  [31:0] i_subB_numberB,	
	input  signed  [ 4:0] i_subA_arrayA_addr,	
	input  signed  [31:0] i_subA_arrayA_datain,	
	output signed  [31:0] o_subA_arrayA_dataout,	
	input                 i_subA_arrayA_r_w,	
	output signed  [31:0] o_subA_ret,	
	input  signed  [31:0] i_subA_numberA	
);

	reg                r_sys_threadTopSub_arbiter3;
	reg         [ 2:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg  signed [31:0] r_sys_threadTopMain_return;
	reg         [ 2:0] r_sys_threadTopMain_caller;
	reg                r_sys_threadTopMain_req;
	reg         [ 3:0] r_sys_threadTopMain_phase;
	reg         [ 2:0] r_sys_threadTopMain_stage;
	reg         [ 2:0] r_sys_threadTopMain_step;
	reg                r_sys_threadTopMain_busy;
	wire        [ 2:0] w_sys_threadTopMain_stage_p1;
	wire        [ 2:0] w_sys_threadTopMain_step_p1;
	reg         [ 2:0] r_sys_threadTopSub_caller;
	reg                r_sys_threadTopSub_req;
	reg         [ 4:0] r_sys_threadTopSub_phase;
	reg         [ 1:0] r_sys_threadTopSub_stage;
	reg         [ 2:0] r_sys_threadTopSub_step;
	reg                r_sys_threadTopSub_busy;
	wire        [ 1:0] w_sys_threadTopSub_stage_p1;
	wire        [ 2:0] w_sys_threadTopSub_step_p1;
	reg         [ 2:0] r_sys_setValueToChildArray_caller;
	reg                r_sys_setValueToChildArray_req;
	reg         [ 3:0] r_sys_setValueToChildArray_phase;
	reg         [ 1:0] r_sys_setValueToChildArray_stage;
	reg         [ 3:0] r_sys_setValueToChildArray_step;
	reg                r_sys_setValueToChildArray_busy;
	wire        [ 1:0] w_sys_setValueToChildArray_stage_p1;
	wire        [ 3:0] w_sys_setValueToChildArray_step_p1;
	wire signed [ 4:0] w_fld_topArray_2_addr_0;
	wire signed [31:0] w_fld_topArray_2_datain_0;
	wire signed [31:0] w_fld_topArray_2_dataout_0;
	wire               w_fld_topArray_2_r_w_0;
	wire               w_fld_topArray_2_ce_0;
	reg  signed [ 4:0] r_fld_topArray_2_addr_1;
	reg  signed [31:0] r_fld_topArray_2_datain_1;
	wire signed [31:0] w_fld_topArray_2_dataout_1;
	reg                r_fld_topArray_2_r_w_1;
	wire               w_fld_topArray_2_ce_1;
	reg  signed [31:0] r_fld_ret_3;
	reg  signed [31:0] r_fld_subRet_4;
	reg  signed [31:0] r_threadTopSub_topArray_5_addr;
	reg  signed [31:0] r_threadTopSub_topArray_5_datain;
	wire signed [31:0] w_threadTopSub_topArray_5_dataout;
	reg                r_threadTopSub_topArray_5_r_w;
	wire signed [31:0] w_threadTopSub_topArray_5_addr;
	wire signed [31:0] w_threadTopSub_topArray_5_datain;
	wire               w_threadTopSub_topArray_5_r_w;
	wire               w_threadTopSub_topArray_5_ce;
	wire               w_threadTopSub_topArray_5_cacheHit;
	reg  signed [31:0] r_threadTopSub_i_6;
	reg  signed [31:0] r_setValueToChildArray_i_7;
	reg  signed [31:0] r_setValueToChildArray_j_8;
	reg  signed [31:0] r_threadTopSub_copy0_i_9;
	reg  signed [31:0] r_setValueToChildArray_copy0_j_10;
	reg  signed [31:0] r_setValueToChildArray_copy1_j_11;
	reg  signed [31:0] r_setValueToChildArray_copy2_j_12;
	reg                r_subB_run_req;
	wire               w_subB_run_busy;
	reg                r_subB_getRet_req;
	wire               w_subB_getRet_busy;
	wire signed [31:0] w_subB_getRet_return;
	wire signed [ 4:0] w_subB_arrayB_addr;
	reg  signed [ 4:0] r_subB_arrayB_addr;
	wire signed [31:0] w_subB_arrayB_datain;
	reg  signed [31:0] r_subB_arrayB_datain;
	wire signed [31:0] w_subB_arrayB_dataout;
	wire               w_subB_arrayB_r_w;
	reg                r_subB_arrayB_r_w;
	reg                r_subA_run_req;
	wire               w_subA_run_busy;
	reg                r_subA_getRet_req;
	wire               w_subA_getRet_busy;
	wire signed [31:0] w_subA_getRet_return;
	wire signed [ 4:0] w_subA_arrayA_addr;
	reg  signed [ 4:0] r_subA_arrayA_addr;
	wire signed [31:0] w_subA_arrayA_datain;
	reg  signed [31:0] r_subA_arrayA_datain;
	wire signed [31:0] w_subA_arrayA_dataout;
	wire               w_subA_arrayA_r_w;
	reg                r_subA_arrayA_r_w;
	reg  signed [31:0] r_sys_tmp0_int;
	reg  signed [31:0] r_sys_tmp1_int;
	reg  signed [31:0] r_sys_tmp2_int;
	reg  signed [31:0] r_sys_tmp3_int;
	reg  signed [31:0] r_sys_tmp4_int;
	reg  signed [31:0] r_sys_tmp5_int;
	reg  signed [31:0] r_sys_tmp6_int;
	reg  signed [31:0] r_sys_tmp7_int;
	reg  signed [31:0] r_sys_tmp8_int;
	reg  signed [31:0] r_sys_tmp9_int;
	reg  signed [31:0] r_sys_tmp10_int;
	wire signed [31:0] w_sys_tmp1;
	wire signed [31:0] w_sys_tmp2;
	wire signed [31:0] w_sys_tmp3;
	wire               w_sys_tmp4;
	wire signed [31:0] w_sys_tmp5;
	wire signed [31:0] w_sys_tmp8;
	wire signed [31:0] w_sys_tmp9;
	wire               w_sys_tmp19;
	wire signed [31:0] w_sys_tmp20;
	wire signed [31:0] w_sys_tmp22;
	wire signed [31:0] w_sys_tmp23;
	wire signed [31:0] w_sys_tmp24;
	wire               w_sys_tmp34;
	wire signed [31:0] w_sys_tmp35;
	wire signed [31:0] w_sys_tmp36;
	wire               w_sys_tmp37;
	wire signed [31:0] w_sys_tmp38;
	wire signed [31:0] w_sys_tmp41;
	wire signed [31:0] w_sys_tmp42;
	wire signed [31:0] w_sys_tmp43;
	wire signed [31:0] w_sys_tmp44;
	wire signed [31:0] w_sys_tmp45;
	wire signed [31:0] w_sys_tmp46;
	wire signed [31:0] w_sys_tmp48;
	wire signed [31:0] w_sys_tmp50;
	wire signed [31:0] w_sys_tmp51;
	wire signed [31:0] w_sys_tmp54;
	wire signed [31:0] w_sys_tmp55;
	wire signed [31:0] w_sys_tmp56;
	wire signed [31:0] w_sys_tmp57;
	wire signed [31:0] w_sys_tmp58;
	wire signed [31:0] w_sys_tmp62;
	wire signed [31:0] w_sys_tmp63;
	wire signed [31:0] w_sys_tmp64;
	wire signed [31:0] w_sys_tmp69;
	wire signed [31:0] w_sys_tmp74;
	wire signed [31:0] w_sys_tmp122;
	wire signed [31:0] w_sys_tmp123;
	wire signed [31:0] w_sys_tmp124;
	wire signed [31:0] w_sys_tmp125;
	wire signed [31:0] w_sys_tmp126;
	wire signed [31:0] w_sys_tmp127;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce & w_threadTopSub_topArray_5_cacheHit;
	assign o_threadTopMain_busy = r_sys_threadTopMain_busy;
	assign o_threadTopMain_return = r_sys_threadTopMain_return;
	assign w_sys_threadTopMain_stage_p1 = (r_sys_threadTopMain_stage + 3'h1);
	assign w_sys_threadTopMain_step_p1 = (r_sys_threadTopMain_step + 3'h1);
	assign w_sys_threadTopSub_stage_p1 = (r_sys_threadTopSub_stage + 2'h1);
	assign w_sys_threadTopSub_step_p1 = (r_sys_threadTopSub_step + 3'h1);
	assign w_sys_setValueToChildArray_stage_p1 = (r_sys_setValueToChildArray_stage + 2'h1);
	assign w_sys_setValueToChildArray_step_p1 = (r_sys_setValueToChildArray_step + 4'h1);
	assign w_fld_topArray_2_addr_0 = ( r_sys_threadTopSub_arbiter3 ? $signed( w_threadTopSub_topArray_5_addr[4:0] ) : 5'sh0 ) ;
	assign w_fld_topArray_2_datain_0 = ( r_sys_threadTopSub_arbiter3 ? w_threadTopSub_topArray_5_datain : 32'sh0 ) ;
	assign w_fld_topArray_2_r_w_0 = ( r_sys_threadTopSub_arbiter3 ? w_threadTopSub_topArray_5_r_w : 1'h0 ) ;
	assign w_fld_topArray_2_ce_0 = w_sys_ce;
	assign w_fld_topArray_2_ce_1 = w_sys_ce;
	assign w_threadTopSub_topArray_5_dataout = ( r_sys_threadTopSub_arbiter3 ? w_fld_topArray_2_dataout_0 : 32'sh0 ) ;
	assign w_threadTopSub_topArray_5_addr = r_threadTopSub_topArray_5_addr;
	assign w_threadTopSub_topArray_5_datain = r_threadTopSub_topArray_5_datain;
	assign w_threadTopSub_topArray_5_r_w = r_threadTopSub_topArray_5_r_w;
	assign w_threadTopSub_topArray_5_ce = w_sys_ce;
	assign w_threadTopSub_topArray_5_cacheHit = ( r_sys_threadTopSub_arbiter3 ? w_sys_boolTrue : w_sys_boolTrue ) ;
	assign w_subB_arrayB_addr = ( (|r_sys_processing_methodID) ? r_subB_arrayB_addr : i_subB_arrayB_addr ) ;
	assign w_subB_arrayB_datain = ( (|r_sys_processing_methodID) ? r_subB_arrayB_datain : i_subB_arrayB_datain ) ;
	assign o_subB_arrayB_dataout = w_subB_arrayB_dataout;
	assign w_subB_arrayB_r_w = ( (|r_sys_processing_methodID) ? r_subB_arrayB_r_w : i_subB_arrayB_r_w ) ;
	assign w_subA_arrayA_addr = ( (|r_sys_processing_methodID) ? r_subA_arrayA_addr : i_subA_arrayA_addr ) ;
	assign w_subA_arrayA_datain = ( (|r_sys_processing_methodID) ? r_subA_arrayA_datain : i_subA_arrayA_datain ) ;
	assign o_subA_arrayA_dataout = w_subA_arrayA_dataout;
	assign w_subA_arrayA_r_w = ( (|r_sys_processing_methodID) ? r_subA_arrayA_r_w : i_subA_arrayA_r_w ) ;
	assign w_sys_tmp1 = (r_fld_ret_3 + r_fld_subRet_4);
	assign w_sys_tmp2 = (r_fld_ret_3 + r_fld_subRet_4);
	assign w_sys_tmp3 = r_fld_ret_3;
	assign w_sys_tmp4 = (r_threadTopSub_i_6 < w_sys_tmp5);
	assign w_sys_tmp5 = 32'sh00000020;
	assign w_sys_tmp8 = (r_threadTopSub_copy0_i_9 + w_sys_intOne);
	assign w_sys_tmp9 = (r_threadTopSub_i_6 + w_sys_intOne);
	assign w_sys_tmp19 = (r_threadTopSub_i_6 < w_sys_tmp20);
	assign w_sys_tmp20 = 32'sh00000020;
	assign w_sys_tmp22 = (r_fld_ret_3 + w_sys_tmp23);
	assign w_sys_tmp23 = w_threadTopSub_topArray_5_dataout;
	assign w_sys_tmp24 = (r_threadTopSub_i_6 + w_sys_intOne);
	assign w_sys_tmp34 = (r_setValueToChildArray_i_7 < w_sys_tmp35);
	assign w_sys_tmp35 = 32'sh00000004;
	assign w_sys_tmp36 = (r_setValueToChildArray_i_7 + w_sys_intOne);
	assign w_sys_tmp37 = (r_setValueToChildArray_j_8 < w_sys_tmp38);
	assign w_sys_tmp38 = 32'sh00000008;
	assign w_sys_tmp41 = (w_sys_tmp42 + r_setValueToChildArray_j_8);
	assign w_sys_tmp42 = (w_sys_tmp43 * r_setValueToChildArray_i_7);
	assign w_sys_tmp43 = 32'sh00000008;
	assign w_sys_tmp44 = (w_sys_tmp45 * w_sys_tmp46);
	assign w_sys_tmp45 = (r_setValueToChildArray_i_7 + r_setValueToChildArray_copy2_j_12);
	assign w_sys_tmp46 = 32'sh0000000f;
	assign w_sys_tmp48 = (r_setValueToChildArray_i_7 * w_sys_tmp43);
	assign w_sys_tmp50 = (w_sys_tmp51 * w_sys_tmp54);
	assign w_sys_tmp51 = w_subA_arrayA_dataout;
	assign w_sys_tmp54 = 32'sh00000022;
	assign w_sys_tmp55 = (r_setValueToChildArray_copy0_j_10 + w_sys_intOne);
	assign w_sys_tmp56 = (r_setValueToChildArray_copy1_j_11 + w_sys_intOne);
	assign w_sys_tmp57 = (r_setValueToChildArray_copy2_j_12 + w_sys_intOne);
	assign w_sys_tmp58 = (r_setValueToChildArray_j_8 + w_sys_intOne);
	assign w_sys_tmp62 = w_sys_tmp58;
	assign w_sys_tmp63 = (r_setValueToChildArray_i_7 + w_sys_tmp64);
	assign w_sys_tmp64 = w_sys_tmp57;
	assign w_sys_tmp69 = w_sys_tmp56;
	assign w_sys_tmp74 = w_sys_tmp55;
	assign w_sys_tmp122 = (w_sys_tmp48 + r_setValueToChildArray_copy1_j_11);
	assign w_sys_tmp123 = (w_sys_tmp42 + r_setValueToChildArray_copy0_j_10);
	assign w_sys_tmp124 = (w_sys_tmp42 + w_sys_tmp62);
	assign w_sys_tmp125 = (w_sys_tmp63 * w_sys_tmp46);
	assign w_sys_tmp126 = (w_sys_tmp48 + w_sys_tmp69);
	assign w_sys_tmp127 = (w_sys_tmp42 + w_sys_tmp74);


	ThreadSubB
		subB_inst(
			.i_fld_arrayB_0_addr_0 (w_subB_arrayB_addr),
			.i_fld_arrayB_0_datain_0 (w_subB_arrayB_datain),
			.o_fld_arrayB_0_dataout_0 (w_subB_arrayB_dataout),
			.i_fld_arrayB_0_r_w_0 (w_subB_arrayB_r_w),
			.i_fld_numberB_2 (i_subB_numberB),
			.o_fld_ret_1 (o_subB_ret),
			.o_getRet_busy (w_subB_getRet_busy),
			.i_getRet_req (r_subB_getRet_req),
			.o_getRet_return (w_subB_getRet_return),
			.o_run_busy (w_subB_run_busy),
			.i_run_req (r_subB_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	ThreadSubA
		subA_inst(
			.i_fld_arrayA_0_addr_0 (w_subA_arrayA_addr),
			.i_fld_arrayA_0_datain_0 (w_subA_arrayA_datain),
			.o_fld_arrayA_0_dataout_0 (w_subA_arrayA_dataout),
			.i_fld_arrayA_0_r_w_0 (w_subA_arrayA_r_w),
			.i_fld_numberA_2 (i_subA_numberA),
			.o_fld_ret_1 (o_subA_ret),
			.o_getRet_busy (w_subA_getRet_busy),
			.i_getRet_req (r_subA_getRet_req),
			.o_getRet_return (w_subA_getRet_return),
			.o_run_busy (w_subA_run_busy),
			.i_run_req (r_subA_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(5), .WORDS(32) )
		dpram_topArray_2(
			.clk (clock),
			.ce_0 (w_fld_topArray_2_ce_0),
			.addr_0 (w_fld_topArray_2_addr_0),
			.datain_0 (w_fld_topArray_2_datain_0),
			.dataout_0 (w_fld_topArray_2_dataout_0),
			.r_w_0 (w_fld_topArray_2_r_w_0),
			.ce_1 (w_fld_topArray_2_ce_1),
			.addr_1 (r_fld_topArray_2_addr_1),
			.datain_1 (r_fld_topArray_2_datain_1),
			.dataout_1 (w_fld_topArray_2_dataout_1),
			.r_w_1 (r_fld_topArray_2_r_w_1)
		);

	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_threadTopSub_arbiter3 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_threadTopMain_phase) 
						4'h2: begin

							case(r_sys_threadTopMain_stage) 
								3'h3: begin
									if((r_sys_threadTopMain_step==3'h1)) begin
										r_sys_threadTopSub_arbiter3 <= w_sys_boolFalse;

									end
									else
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_sys_threadTopSub_arbiter3 <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 3'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h0: begin
					r_sys_processing_methodID <= ((i_threadTopMain_req) ? 3'h1 : r_sys_processing_methodID);
				end

				3'h1: begin

					case(r_sys_threadTopMain_phase) 
						4'h2: begin

							case(r_sys_threadTopMain_stage) 
								3'h0: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_sys_processing_methodID <= 3'h3;

									end
								end

								3'h3: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_sys_processing_methodID <= 3'h2;

									end
								end

							endcase
						end

						4'h9: begin
							r_sys_processing_methodID <= r_sys_threadTopMain_caller;
						end

					endcase
				end

				3'h2: begin

					case(r_sys_threadTopSub_phase) 
						5'h10: begin
							r_sys_processing_methodID <= r_sys_threadTopSub_caller;
						end

					endcase
				end

				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'he: begin
							r_sys_processing_methodID <= r_sys_setValueToChildArray_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_threadTopMain_return <= 32'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_threadTopMain_phase) 
						4'h6: begin
							r_sys_threadTopMain_return <= w_sys_tmp3;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_threadTopMain_caller <= 3'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_threadTopMain_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_threadTopMain_phase <= 4'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_threadTopMain_phase) 
						4'h0: begin
							r_sys_threadTopMain_phase <= 4'h2;
						end

						4'h2: begin

							case(r_sys_threadTopMain_stage) 
								3'h3: begin
									if((r_sys_threadTopMain_step==3'h1)) begin
										r_sys_threadTopMain_phase <= 4'h4;

									end
								end

							endcase
						end

						4'h4: begin

							case(r_sys_threadTopMain_stage) 
								3'h1: begin
									if((r_sys_threadTopMain_step==3'h1)) begin
										r_sys_threadTopMain_phase <= 4'h5;

									end
								end

							endcase
						end

						4'h5: begin

							case(r_sys_threadTopMain_stage) 
								3'h3: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_sys_threadTopMain_phase <= 4'h7;

									end
								end

							endcase
						end

						4'h6: begin
							r_sys_threadTopMain_phase <= 4'h9;
						end

						4'h7: begin

							case(r_sys_threadTopMain_stage) 
								3'h0: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_sys_threadTopMain_phase <= 4'h6;

									end
								end

							endcase
						end

						4'h9: begin
							r_sys_threadTopMain_phase <= 4'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_threadTopMain_stage <= 3'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_threadTopMain_phase) 
						4'h2: begin

							case(r_sys_threadTopMain_stage) 
								3'h0: begin
									if((r_sys_threadTopMain_step==3'h1)) begin
										r_sys_threadTopMain_stage <= w_sys_threadTopMain_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_threadTopMain_step==3'h1)) begin
										r_sys_threadTopMain_stage <= w_sys_threadTopMain_stage_p1;

									end
								end

								3'h2: begin
									if((r_sys_threadTopMain_step==3'h1)) begin
										r_sys_threadTopMain_stage <= w_sys_threadTopMain_stage_p1;

									end
								end

								3'h3: begin
									if((r_sys_threadTopMain_step==3'h1)) begin
										r_sys_threadTopMain_stage <= 3'h0;

									end
								end

							endcase
						end

						4'h4: begin

							case(r_sys_threadTopMain_stage) 
								3'h0: begin
									if((r_sys_threadTopMain_step==3'h1)) begin
										r_sys_threadTopMain_stage <= w_sys_threadTopMain_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_threadTopMain_step==3'h1)) begin
										r_sys_threadTopMain_stage <= 3'h0;

									end
								end

							endcase
						end

						4'h5: begin

							case(r_sys_threadTopMain_stage) 
								3'h0: begin
									if((r_sys_threadTopMain_step==3'h3)) begin
										r_sys_threadTopMain_stage <= w_sys_threadTopMain_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_sys_threadTopMain_stage <= w_sys_threadTopMain_stage_p1;

									end
								end

								3'h2: begin
									if((r_sys_threadTopMain_step==3'h3)) begin
										r_sys_threadTopMain_stage <= w_sys_threadTopMain_stage_p1;

									end
								end

								3'h3: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_sys_threadTopMain_stage <= 3'h0;

									end
								end

							endcase
						end

						4'h7: begin

							case(r_sys_threadTopMain_stage) 
								3'h0: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_sys_threadTopMain_stage <= 3'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_threadTopMain_step <= 3'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_threadTopMain_phase) 
						4'h2: begin

							case(r_sys_threadTopMain_stage) 
								3'h0: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_sys_threadTopMain_step <= w_sys_threadTopMain_step_p1;

									end
									else
									if((r_sys_threadTopMain_step==3'h1)) begin
										r_sys_threadTopMain_step <= 3'h0;

									end
								end

								3'h1: begin
									if((r_sys_threadTopMain_step==3'h1)) begin
										r_sys_threadTopMain_step <= 3'h0;

									end
									else
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_sys_threadTopMain_step <= w_sys_threadTopMain_step_p1;

									end
								end

								3'h2: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_sys_threadTopMain_step <= w_sys_threadTopMain_step_p1;

									end
									else
									if((r_sys_threadTopMain_step==3'h1)) begin
										r_sys_threadTopMain_step <= 3'h0;

									end
								end

								3'h3: begin
									if((r_sys_threadTopMain_step==3'h1)) begin
										r_sys_threadTopMain_step <= 3'h0;

									end
									else
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_sys_threadTopMain_step <= w_sys_threadTopMain_step_p1;

									end
								end

							endcase
						end

						4'h4: begin

							case(r_sys_threadTopMain_stage) 
								3'h0: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_sys_threadTopMain_step <= ((w_subA_run_busy) ? r_sys_threadTopMain_step : w_sys_threadTopMain_step_p1);

									end
									else
									if((r_sys_threadTopMain_step==3'h1)) begin
										r_sys_threadTopMain_step <= 3'h0;

									end
								end

								3'h1: begin
									if((r_sys_threadTopMain_step==3'h1)) begin
										r_sys_threadTopMain_step <= 3'h0;

									end
									else
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_sys_threadTopMain_step <= ((w_subB_run_busy) ? r_sys_threadTopMain_step : w_sys_threadTopMain_step_p1);

									end
								end

							endcase
						end

						4'h5: begin

							case(r_sys_threadTopMain_stage) 
								3'h0: begin
									if((r_sys_threadTopMain_step==3'h3)) begin
										r_sys_threadTopMain_step <= 3'h0;

									end
									else
									if((r_sys_threadTopMain_step==3'h0) || (r_sys_threadTopMain_step==3'h1)) begin
										r_sys_threadTopMain_step <= w_sys_threadTopMain_step_p1;

									end
									else
									if((r_sys_threadTopMain_step==3'h2)) begin
										r_sys_threadTopMain_step <= ((w_subA_getRet_busy) ? r_sys_threadTopMain_step : w_sys_threadTopMain_step_p1);

									end
								end

								3'h1: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_sys_threadTopMain_step <= 3'h0;

									end
								end

								3'h2: begin
									if((r_sys_threadTopMain_step==3'h3)) begin
										r_sys_threadTopMain_step <= 3'h0;

									end
									else
									if((r_sys_threadTopMain_step==3'h0) || (r_sys_threadTopMain_step==3'h1)) begin
										r_sys_threadTopMain_step <= w_sys_threadTopMain_step_p1;

									end
									else
									if((r_sys_threadTopMain_step==3'h2)) begin
										r_sys_threadTopMain_step <= ((w_subB_getRet_busy) ? r_sys_threadTopMain_step : w_sys_threadTopMain_step_p1);

									end
								end

								3'h3: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_sys_threadTopMain_step <= 3'h0;

									end
								end

							endcase
						end

						4'h7: begin

							case(r_sys_threadTopMain_stage) 
								3'h0: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_sys_threadTopMain_step <= 3'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_threadTopMain_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h0: begin
					r_sys_threadTopMain_busy <= ((i_threadTopMain_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				3'h1: begin

					case(r_sys_threadTopMain_phase) 
						4'h0: begin
							r_sys_threadTopMain_busy <= w_sys_boolTrue;
						end

						4'h9: begin
							r_sys_threadTopMain_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_threadTopSub_caller <= 3'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_threadTopMain_phase) 
						4'h2: begin

							case(r_sys_threadTopMain_stage) 
								3'h3: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_sys_threadTopSub_caller <= r_sys_processing_methodID;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_threadTopSub_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_threadTopSub_phase <= 5'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_threadTopSub_phase) 
						5'h0: begin
							r_sys_threadTopSub_phase <= 5'h2;
						end

						5'h2: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((r_sys_threadTopSub_step==3'h0)) begin
										r_sys_threadTopSub_phase <= 5'h4;

									end
								end

							endcase
						end

						5'h4: begin

							case(r_sys_threadTopSub_stage) 
								2'h1: begin
									if((r_sys_threadTopSub_step==3'h0)) begin
										r_sys_threadTopSub_phase <= 5'h5;

									end
								end

							endcase
						end

						5'h5: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((r_sys_threadTopSub_step==3'h0)) begin
										r_sys_threadTopSub_phase <= ((w_sys_tmp4) ? 5'h8 : 5'ha);

									end
								end

							endcase
						end

						5'h8: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((r_sys_threadTopSub_step==3'h3)) begin
										r_sys_threadTopSub_phase <= 5'h5;

									end
								end

							endcase
						end

						5'ha: begin

							case(r_sys_threadTopSub_stage) 
								2'h1: begin
									if((r_sys_threadTopSub_step==3'h0)) begin
										r_sys_threadTopSub_phase <= 5'hb;

									end
								end

							endcase
						end

						5'hb: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((r_sys_threadTopSub_step==3'h0)) begin
										r_sys_threadTopSub_phase <= ((w_sys_tmp19) ? 5'he : 5'h10);

									end
								end

							endcase
						end

						5'he: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((r_sys_threadTopSub_step==3'h5)) begin
										r_sys_threadTopSub_phase <= 5'hb;

									end
								end

							endcase
						end

						5'h10: begin
							r_sys_threadTopSub_phase <= 5'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_threadTopSub_stage <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_threadTopSub_phase) 
						5'h2: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((r_sys_threadTopSub_step==3'h0)) begin
										r_sys_threadTopSub_stage <= 2'h0;

									end
								end

							endcase
						end

						5'h4: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((r_sys_threadTopSub_step==3'h0)) begin
										r_sys_threadTopSub_stage <= w_sys_threadTopSub_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_threadTopSub_step==3'h0)) begin
										r_sys_threadTopSub_stage <= 2'h0;

									end
								end

							endcase
						end

						5'h5: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((r_sys_threadTopSub_step==3'h0)) begin
										r_sys_threadTopSub_stage <= 2'h0;

									end
								end

							endcase
						end

						5'h8: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((r_sys_threadTopSub_step==3'h3)) begin
										r_sys_threadTopSub_stage <= 2'h0;

									end
								end

							endcase
						end

						5'ha: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((r_sys_threadTopSub_step==3'h0)) begin
										r_sys_threadTopSub_stage <= w_sys_threadTopSub_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_threadTopSub_step==3'h0)) begin
										r_sys_threadTopSub_stage <= 2'h0;

									end
								end

							endcase
						end

						5'hb: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((r_sys_threadTopSub_step==3'h0)) begin
										r_sys_threadTopSub_stage <= 2'h0;

									end
								end

							endcase
						end

						5'he: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((r_sys_threadTopSub_step==3'h5)) begin
										r_sys_threadTopSub_stage <= 2'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_threadTopSub_step <= 3'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_threadTopSub_phase) 
						5'h2: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((r_sys_threadTopSub_step==3'h0)) begin
										r_sys_threadTopSub_step <= 3'h0;

									end
								end

							endcase
						end

						5'h4: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((r_sys_threadTopSub_step==3'h0)) begin
										r_sys_threadTopSub_step <= 3'h0;

									end
								end

								2'h1: begin
									if((r_sys_threadTopSub_step==3'h0)) begin
										r_sys_threadTopSub_step <= 3'h0;

									end
								end

							endcase
						end

						5'h5: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((r_sys_threadTopSub_step==3'h0)) begin
										r_sys_threadTopSub_step <= 3'h0;

									end
								end

							endcase
						end

						5'h8: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((r_sys_threadTopSub_step==3'h3)) begin
										r_sys_threadTopSub_step <= 3'h0;

									end
									else
									if((r_sys_threadTopSub_step==3'h0) || (r_sys_threadTopSub_step==3'h1) || (r_sys_threadTopSub_step==3'h2)) begin
										r_sys_threadTopSub_step <= w_sys_threadTopSub_step_p1;

									end
								end

							endcase
						end

						5'ha: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((r_sys_threadTopSub_step==3'h0)) begin
										r_sys_threadTopSub_step <= 3'h0;

									end
								end

								2'h1: begin
									if((r_sys_threadTopSub_step==3'h0)) begin
										r_sys_threadTopSub_step <= 3'h0;

									end
								end

							endcase
						end

						5'hb: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((r_sys_threadTopSub_step==3'h0)) begin
										r_sys_threadTopSub_step <= 3'h0;

									end
								end

							endcase
						end

						5'he: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((r_sys_threadTopSub_step==3'h5)) begin
										r_sys_threadTopSub_step <= 3'h0;

									end
									else
									if((3'h0<=r_sys_threadTopSub_step && r_sys_threadTopSub_step<=3'h4)) begin
										r_sys_threadTopSub_step <= w_sys_threadTopSub_step_p1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_threadTopSub_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_threadTopSub_phase) 
						5'h0: begin
							r_sys_threadTopSub_busy <= w_sys_boolTrue;
						end

						5'h10: begin
							r_sys_threadTopSub_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_setValueToChildArray_caller <= 3'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_threadTopMain_phase) 
						4'h2: begin

							case(r_sys_threadTopMain_stage) 
								3'h0: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_sys_setValueToChildArray_caller <= r_sys_processing_methodID;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_setValueToChildArray_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_setValueToChildArray_phase <= 4'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h0: begin
							r_sys_setValueToChildArray_phase <= 4'h3;
						end

						4'h3: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_sys_setValueToChildArray_phase <= 4'h4;

									end
								end

							endcase
						end

						4'h4: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_sys_setValueToChildArray_phase <= ((w_sys_tmp34) ? 4'h8 : 4'he);

									end
								end

							endcase
						end

						4'h5: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_sys_setValueToChildArray_phase <= 4'h4;

									end
								end

							endcase
						end

						4'h8: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h1: begin
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_sys_setValueToChildArray_phase <= 4'h9;

									end
								end

							endcase
						end

						4'h9: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_sys_setValueToChildArray_phase <= ((w_sys_tmp37) ? 4'hc : 4'h5);

									end
								end

							endcase
						end

						4'hc: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h9)) begin
										r_sys_setValueToChildArray_phase <= 4'h9;

									end
								end

							endcase
						end

						4'he: begin
							r_sys_setValueToChildArray_phase <= 4'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_setValueToChildArray_stage <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h3: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_sys_setValueToChildArray_stage <= 2'h0;

									end
								end

							endcase
						end

						4'h4: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_sys_setValueToChildArray_stage <= 2'h0;

									end
								end

							endcase
						end

						4'h5: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_sys_setValueToChildArray_stage <= 2'h0;

									end
								end

							endcase
						end

						4'h8: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_sys_setValueToChildArray_stage <= w_sys_setValueToChildArray_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_sys_setValueToChildArray_stage <= 2'h0;

									end
								end

							endcase
						end

						4'h9: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_sys_setValueToChildArray_stage <= 2'h0;

									end
								end

							endcase
						end

						4'hc: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h9)) begin
										r_sys_setValueToChildArray_stage <= 2'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_setValueToChildArray_step <= 4'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h3: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_sys_setValueToChildArray_step <= 4'h0;

									end
								end

							endcase
						end

						4'h4: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_sys_setValueToChildArray_step <= 4'h0;

									end
								end

							endcase
						end

						4'h5: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_sys_setValueToChildArray_step <= 4'h0;

									end
								end

							endcase
						end

						4'h8: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_sys_setValueToChildArray_step <= 4'h0;

									end
								end

								2'h1: begin
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_sys_setValueToChildArray_step <= 4'h0;

									end
								end

							endcase
						end

						4'h9: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_sys_setValueToChildArray_step <= 4'h0;

									end
								end

							endcase
						end

						4'hc: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((4'h0<=r_sys_setValueToChildArray_step && r_sys_setValueToChildArray_step<=4'h8)) begin
										r_sys_setValueToChildArray_step <= w_sys_setValueToChildArray_step_p1;

									end
									else
									if((r_sys_setValueToChildArray_step==4'h9)) begin
										r_sys_setValueToChildArray_step <= 4'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_setValueToChildArray_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h0: begin
							r_sys_setValueToChildArray_busy <= w_sys_boolTrue;
						end

						4'he: begin
							r_sys_setValueToChildArray_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_topArray_2_addr_1 <= 5'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_topArray_2_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_threadTopMain_phase) 
						4'h9: begin
							r_fld_topArray_2_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

				3'h2: begin

					case(r_sys_threadTopSub_phase) 
						5'h10: begin
							r_fld_topArray_2_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'he: begin
							r_fld_topArray_2_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_ret_3 <= w_sys_intZero;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_threadTopMain_phase) 
						4'h5: begin

							case(r_sys_threadTopMain_stage) 
								3'h1: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_fld_ret_3 <= w_sys_tmp1;

									end
								end

								3'h3: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_fld_ret_3 <= w_sys_tmp2;

									end
								end

							endcase
						end

					endcase
				end

				3'h2: begin

					case(r_sys_threadTopSub_phase) 
						5'he: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((3'h2<=r_sys_threadTopSub_step && r_sys_threadTopSub_step<=3'h5)) begin
										r_fld_ret_3 <= w_sys_tmp22;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_subRet_4 <= w_sys_intZero;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_threadTopMain_phase) 
						4'h5: begin

							case(r_sys_threadTopMain_stage) 
								3'h0: begin
									if((r_sys_threadTopMain_step==3'h3)) begin
										r_fld_subRet_4 <= w_subA_getRet_return;

									end
								end

								3'h2: begin
									if((r_sys_threadTopMain_step==3'h3)) begin
										r_fld_subRet_4 <= w_subB_getRet_return;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_threadTopSub_topArray_5_addr <= 32'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_threadTopSub_phase) 
						5'h8: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((r_sys_threadTopSub_step==3'h1) || (r_sys_threadTopSub_step==3'h2) || (r_sys_threadTopSub_step==3'h3)) begin
										r_threadTopSub_topArray_5_addr <= r_sys_tmp1_int;

									end
									else
									if((r_sys_threadTopSub_step==3'h0)) begin
										r_threadTopSub_topArray_5_addr <= r_threadTopSub_i_6;

									end
								end

							endcase
						end

						5'he: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((r_sys_threadTopSub_step==3'h0)) begin
										r_threadTopSub_topArray_5_addr <= r_threadTopSub_i_6;

									end
									else
									if((r_sys_threadTopSub_step==3'h1) || (r_sys_threadTopSub_step==3'h2) || (r_sys_threadTopSub_step==3'h3)) begin
										r_threadTopSub_topArray_5_addr <= r_sys_tmp0_int;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_threadTopSub_phase) 
						5'h8: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((r_sys_threadTopSub_step==3'h0)) begin
										r_threadTopSub_topArray_5_datain <= r_threadTopSub_copy0_i_9;

									end
									else
									if((r_sys_threadTopSub_step==3'h1) || (r_sys_threadTopSub_step==3'h2) || (r_sys_threadTopSub_step==3'h3)) begin
										r_threadTopSub_topArray_5_datain <= r_sys_tmp0_int;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_threadTopSub_topArray_5_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_threadTopMain_phase) 
						4'h9: begin
							r_threadTopSub_topArray_5_r_w <= w_sys_boolFalse;
						end

					endcase
				end

				3'h2: begin

					case(r_sys_threadTopSub_phase) 
						5'h8: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((3'h0<=r_sys_threadTopSub_step && r_sys_threadTopSub_step<=3'h3)) begin
										r_threadTopSub_topArray_5_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						5'he: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((3'h0<=r_sys_threadTopSub_step && r_sys_threadTopSub_step<=3'h3)) begin
										r_threadTopSub_topArray_5_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						5'h10: begin
							r_threadTopSub_topArray_5_r_w <= w_sys_boolFalse;
						end

					endcase
				end

				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'he: begin
							r_threadTopSub_topArray_5_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_threadTopSub_phase) 
						5'h4: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((r_sys_threadTopSub_step==3'h0)) begin
										r_threadTopSub_i_6 <= w_sys_intZero;

									end
								end

							endcase
						end

						5'h8: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((3'h0<=r_sys_threadTopSub_step && r_sys_threadTopSub_step<=3'h3)) begin
										r_threadTopSub_i_6 <= w_sys_tmp9;

									end
								end

							endcase
						end

						5'ha: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((r_sys_threadTopSub_step==3'h0)) begin
										r_threadTopSub_i_6 <= w_sys_intZero;

									end
								end

							endcase
						end

						5'he: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((3'h0<=r_sys_threadTopSub_step && r_sys_threadTopSub_step<=3'h3)) begin
										r_threadTopSub_i_6 <= w_sys_tmp24;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h3: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_setValueToChildArray_i_7 <= w_sys_intZero;

									end
								end

							endcase
						end

						4'h5: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_setValueToChildArray_i_7 <= w_sys_tmp36;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h8: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_setValueToChildArray_j_8 <= w_sys_intZero;

									end
								end

							endcase
						end

						4'hc: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((4'h0<=r_sys_setValueToChildArray_step && r_sys_setValueToChildArray_step<=4'h3)) begin
										r_setValueToChildArray_j_8 <= w_sys_tmp58;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_threadTopSub_phase) 
						5'h4: begin

							case(r_sys_threadTopSub_stage) 
								2'h1: begin
									if((r_sys_threadTopSub_step==3'h0)) begin
										r_threadTopSub_copy0_i_9 <= r_threadTopSub_i_6;

									end
								end

							endcase
						end

						5'h8: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((3'h0<=r_sys_threadTopSub_step && r_sys_threadTopSub_step<=3'h3)) begin
										r_threadTopSub_copy0_i_9 <= w_sys_tmp8;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h8: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h1: begin
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_setValueToChildArray_copy0_j_10 <= r_setValueToChildArray_j_8;

									end
								end

							endcase
						end

						4'hc: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((4'h0<=r_sys_setValueToChildArray_step && r_sys_setValueToChildArray_step<=4'h3)) begin
										r_setValueToChildArray_copy0_j_10 <= w_sys_tmp55;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h8: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h1: begin
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_setValueToChildArray_copy1_j_11 <= r_setValueToChildArray_j_8;

									end
								end

							endcase
						end

						4'hc: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((4'h0<=r_sys_setValueToChildArray_step && r_sys_setValueToChildArray_step<=4'h3)) begin
										r_setValueToChildArray_copy1_j_11 <= w_sys_tmp56;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h8: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h1: begin
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_setValueToChildArray_copy2_j_12 <= r_setValueToChildArray_j_8;

									end
								end

							endcase
						end

						4'hc: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((4'h0<=r_sys_setValueToChildArray_step && r_sys_setValueToChildArray_step<=4'h3)) begin
										r_setValueToChildArray_copy2_j_12 <= w_sys_tmp57;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_subB_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_threadTopMain_phase) 
						4'h2: begin

							case(r_sys_threadTopMain_stage) 
								3'h2: begin
									if((r_sys_threadTopMain_step==3'h1)) begin
										r_subB_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_subB_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_subB_getRet_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_threadTopMain_phase) 
						4'h5: begin

							case(r_sys_threadTopMain_stage) 
								3'h2: begin
									if((r_sys_threadTopMain_step==3'h1)) begin
										r_subB_getRet_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_subB_getRet_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_subB_arrayB_addr <= 5'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'hc: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h9)) begin
										r_subB_arrayB_addr <= $signed( r_sys_tmp1_int[4:0] );

									end
									else
									if((r_sys_setValueToChildArray_step==4'h7)) begin
										r_subB_arrayB_addr <= $signed( r_sys_tmp4_int[4:0] );

									end
									else
									if((r_sys_setValueToChildArray_step==4'h3)) begin
										r_subB_arrayB_addr <= $signed( r_sys_tmp5_int[4:0] );

									end
									else
									if((r_sys_setValueToChildArray_step==4'h5)) begin
										r_subB_arrayB_addr <= $signed( r_sys_tmp6_int[4:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'hc: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h3) || (r_sys_setValueToChildArray_step==4'h5) || (r_sys_setValueToChildArray_step==4'h7) || (r_sys_setValueToChildArray_step==4'h9)) begin
										r_subB_arrayB_datain <= w_sys_tmp50;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_subB_arrayB_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_threadTopMain_phase) 
						4'h2: begin

							case(r_sys_threadTopMain_stage) 
								3'h0: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_subB_arrayB_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_subB_arrayB_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_subB_arrayB_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_subB_arrayB_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						4'h5: begin

							case(r_sys_threadTopMain_stage) 
								3'h0: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_subB_arrayB_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_subB_arrayB_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						4'h9: begin
							r_subB_arrayB_r_w <= w_sys_boolFalse;
						end

					endcase
				end

				3'h2: begin

					case(r_sys_threadTopSub_phase) 
						5'h10: begin
							r_subB_arrayB_r_w <= w_sys_boolFalse;
						end

					endcase
				end

				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'hc: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h3) || (r_sys_setValueToChildArray_step==4'h5) || (r_sys_setValueToChildArray_step==4'h7) || (r_sys_setValueToChildArray_step==4'h9)) begin
										r_subB_arrayB_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						4'he: begin
							r_subB_arrayB_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_subA_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_threadTopMain_phase) 
						4'h2: begin

							case(r_sys_threadTopMain_stage) 
								3'h1: begin
									if((r_sys_threadTopMain_step==3'h1)) begin
										r_subA_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_subA_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_subA_getRet_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_threadTopMain_phase) 
						4'h5: begin

							case(r_sys_threadTopMain_stage) 
								3'h0: begin
									if((r_sys_threadTopMain_step==3'h1)) begin
										r_subA_getRet_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_subA_getRet_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_subA_arrayA_addr <= 5'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'hc: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h2) || (r_sys_setValueToChildArray_step==4'h6)) begin
										r_subA_arrayA_addr <= $signed( r_sys_tmp9_int[4:0] );

									end
									else
									if((r_sys_setValueToChildArray_step==4'h1) || (r_sys_setValueToChildArray_step==4'h5)) begin
										r_subA_arrayA_addr <= $signed( r_sys_tmp8_int[4:0] );

									end
									else
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_subA_arrayA_addr <= $signed( w_sys_tmp41[4:0] );

									end
									else
									if((r_sys_setValueToChildArray_step==4'h4)) begin
										r_subA_arrayA_addr <= $signed( r_sys_tmp3_int[4:0] );

									end
									else
									if((r_sys_setValueToChildArray_step==4'h7)) begin
										r_subA_arrayA_addr <= $signed( r_sys_tmp0_int[4:0] );

									end
									else
									if((r_sys_setValueToChildArray_step==4'h3)) begin
										r_subA_arrayA_addr <= $signed( r_sys_tmp7_int[4:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'hc: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h2) || (r_sys_setValueToChildArray_step==4'h6)) begin
										r_subA_arrayA_datain <= r_sys_tmp10_int;

									end
									else
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_subA_arrayA_datain <= w_sys_tmp44;

									end
									else
									if((r_sys_setValueToChildArray_step==4'h4)) begin
										r_subA_arrayA_datain <= r_sys_tmp2_int;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_subA_arrayA_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_threadTopMain_phase) 
						4'h2: begin

							case(r_sys_threadTopMain_stage) 
								3'h0: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_subA_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_subA_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_subA_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_subA_arrayA_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						4'h5: begin

							case(r_sys_threadTopMain_stage) 
								3'h0: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_subA_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_threadTopMain_step==3'h0)) begin
										r_subA_arrayA_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						4'h9: begin
							r_subA_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

				3'h2: begin

					case(r_sys_threadTopSub_phase) 
						5'h10: begin
							r_subA_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'hc: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h1) || (r_sys_setValueToChildArray_step==4'h3) || (r_sys_setValueToChildArray_step==4'h5) || (r_sys_setValueToChildArray_step==4'h7)) begin
										r_subA_arrayA_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_setValueToChildArray_step==4'h0) || (r_sys_setValueToChildArray_step==4'h2) || (r_sys_setValueToChildArray_step==4'h4) || (r_sys_setValueToChildArray_step==4'h6)) begin
										r_subA_arrayA_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						4'he: begin
							r_subA_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_threadTopSub_phase) 
						5'h8: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((r_sys_threadTopSub_step==3'h0) || (r_sys_threadTopSub_step==3'h1) || (r_sys_threadTopSub_step==3'h2)) begin
										r_sys_tmp0_int <= w_sys_tmp8;

									end
								end

							endcase
						end

						5'he: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((r_sys_threadTopSub_step==3'h0) || (r_sys_threadTopSub_step==3'h1) || (r_sys_threadTopSub_step==3'h2)) begin
										r_sys_tmp0_int <= w_sys_tmp24;

									end
								end

							endcase
						end

					endcase
				end

				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'hc: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h2)) begin
										r_sys_tmp0_int <= w_sys_tmp127;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_threadTopSub_phase) 
						5'h8: begin

							case(r_sys_threadTopSub_stage) 
								2'h0: begin
									if((r_sys_threadTopSub_step==3'h0) || (r_sys_threadTopSub_step==3'h1) || (r_sys_threadTopSub_step==3'h2)) begin
										r_sys_tmp1_int <= w_sys_tmp9;

									end
								end

							endcase
						end

					endcase
				end

				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'hc: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h2)) begin
										r_sys_tmp1_int <= w_sys_tmp126;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'hc: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h1)) begin
										r_sys_tmp2_int <= w_sys_tmp125;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'hc: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h1)) begin
										r_sys_tmp3_int <= w_sys_tmp124;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'hc: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h1)) begin
										r_sys_tmp4_int <= w_sys_tmp126;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'hc: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_sys_tmp5_int <= w_sys_tmp122;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'hc: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_sys_tmp6_int <= w_sys_tmp126;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'hc: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_sys_tmp7_int <= w_sys_tmp127;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'hc: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h0)) begin
										r_sys_tmp8_int <= w_sys_tmp123;

									end
									else
									if((r_sys_setValueToChildArray_step==4'h1)) begin
										r_sys_tmp8_int <= w_sys_tmp127;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'hc: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h0) || (r_sys_setValueToChildArray_step==4'h2)) begin
										r_sys_tmp9_int <= w_sys_tmp124;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_setValueToChildArray_phase) 
						4'hc: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==4'h0) || (r_sys_setValueToChildArray_step==4'h2)) begin
										r_sys_tmp10_int <= w_sys_tmp125;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
