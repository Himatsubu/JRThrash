/*
TimeStamp:	2016/11/11		13:0
*/


module P3_2dim(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy,	
	output signed  [31:0] o_run_return	
);

	reg         [31:0] r_ip_AddFloat_portA_0;
	reg         [31:0] r_ip_AddFloat_portB_0;
	wire        [31:0] w_ip_AddFloat_result_0;
	reg         [31:0] r_ip_MultFloat_multiplicand_0;
	reg         [31:0] r_ip_MultFloat_multiplier_0;
	wire        [31:0] w_ip_MultFloat_product_0;
	reg  signed [31:0] r_ip_FixedToFloat_fixed_0;
	wire        [31:0] w_ip_FixedToFloat_floating_0;
	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [31:0] r_sys_run_return;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 9:0] r_sys_run_phase;
	reg         [ 5:0] r_sys_run_stage;
	reg         [ 5:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 5:0] w_sys_run_stage_p1;
	wire        [ 5:0] w_sys_run_step_p1;
	wire signed [14:0] w_fld_T_0_addr_0;
	wire        [31:0] w_fld_T_0_datain_0;
	wire        [31:0] w_fld_T_0_dataout_0;
	wire               w_fld_T_0_r_w_0;
	wire               w_fld_T_0_ce_0;
	reg  signed [14:0] r_fld_T_0_addr_1;
	reg         [31:0] r_fld_T_0_datain_1;
	wire        [31:0] w_fld_T_0_dataout_1;
	reg                r_fld_T_0_r_w_1;
	wire               w_fld_T_0_ce_1;
	wire signed [14:0] w_fld_TT_1_addr_0;
	wire        [31:0] w_fld_TT_1_datain_0;
	wire        [31:0] w_fld_TT_1_dataout_0;
	wire               w_fld_TT_1_r_w_0;
	wire               w_fld_TT_1_ce_0;
	reg  signed [14:0] r_fld_TT_1_addr_1;
	reg         [31:0] r_fld_TT_1_datain_1;
	wire        [31:0] w_fld_TT_1_dataout_1;
	reg                r_fld_TT_1_r_w_1;
	wire               w_fld_TT_1_ce_1;
	wire signed [14:0] w_fld_U_2_addr_0;
	wire        [31:0] w_fld_U_2_datain_0;
	wire        [31:0] w_fld_U_2_dataout_0;
	wire               w_fld_U_2_r_w_0;
	wire               w_fld_U_2_ce_0;
	reg  signed [14:0] r_fld_U_2_addr_1;
	reg         [31:0] r_fld_U_2_datain_1;
	wire        [31:0] w_fld_U_2_dataout_1;
	reg                r_fld_U_2_r_w_1;
	wire               w_fld_U_2_ce_1;
	reg  signed [31:0] r_run_k_35;
	reg  signed [31:0] r_run_j_36;
	reg  signed [31:0] r_run_n_37;
	reg  signed [31:0] r_run_mx_38;
	reg  signed [31:0] r_run_my_39;
	reg         [31:0] r_run_dt_40;
	reg         [31:0] r_run_dx_41;
	reg         [31:0] r_run_dy_42;
	reg         [31:0] r_run_r1_43;
	reg         [31:0] r_run_r2_44;
	reg         [31:0] r_run_r3_45;
	reg         [31:0] r_run_r4_46;
	reg         [31:0] r_run_YY_47;
	reg  signed [31:0] r_run_kx_48;
	reg  signed [31:0] r_run_ky_49;
	reg  signed [31:0] r_run_nlast_50;
	reg  signed [31:0] r_run_tmpj_51;
	reg  signed [31:0] r_run_copy0_j_52;
	reg  signed [31:0] r_run_copy1_j_53;
	reg  signed [31:0] r_run_copy0_j_54;
	reg  signed [31:0] r_run_copy0_j_55;
	reg  signed [31:0] r_run_copy1_j_56;
	reg  signed [31:0] r_run_copy2_j_57;
	reg  signed [31:0] r_run_copy0_j_58;
	reg  signed [31:0] r_run_copy1_j_59;
	reg  signed [31:0] r_run_copy2_j_60;
	reg  signed [31:0] r_run_copy0_j_61;
	reg  signed [31:0] r_run_copy1_j_62;
	reg  signed [31:0] r_run_copy2_j_63;
	reg  signed [31:0] r_run_copy0_j_64;
	reg  signed [31:0] r_run_copy1_j_65;
	reg  signed [31:0] r_run_copy2_j_66;
	reg  signed [31:0] r_run_copy0_j_67;
	reg  signed [31:0] r_run_copy1_j_68;
	reg  signed [31:0] r_run_copy2_j_69;
	reg  signed [31:0] r_run_copy0_j_70;
	reg  signed [31:0] r_run_copy1_j_71;
	reg  signed [31:0] r_run_copy2_j_72;
	reg  signed [31:0] r_run_copy0_j_73;
	reg  signed [31:0] r_run_copy1_j_74;
	reg  signed [31:0] r_run_copy2_j_75;
	reg  signed [31:0] r_run_copy0_j_76;
	reg  signed [31:0] r_run_copy1_j_77;
	reg  signed [31:0] r_run_copy2_j_78;
	reg  signed [31:0] r_run_copy0_j_79;
	reg  signed [31:0] r_run_copy1_j_80;
	reg  signed [31:0] r_run_copy2_j_81;
	reg  signed [31:0] r_run_copy0_j_82;
	reg  signed [31:0] r_run_copy1_j_83;
	reg  signed [31:0] r_run_copy2_j_84;
	reg  signed [31:0] r_run_copy0_j_85;
	reg  signed [31:0] r_run_copy1_j_86;
	reg  signed [31:0] r_run_copy2_j_87;
	reg  signed [31:0] r_run_copy0_j_88;
	reg  signed [31:0] r_run_copy1_j_89;
	reg  signed [31:0] r_run_copy2_j_90;
	reg  signed [31:0] r_run_copy0_j_91;
	reg  signed [31:0] r_run_copy1_j_92;
	reg  signed [31:0] r_run_copy2_j_93;
	reg  signed [31:0] r_run_copy0_j_94;
	reg  signed [31:0] r_run_copy1_j_95;
	reg  signed [31:0] r_run_copy2_j_96;
	reg  signed [31:0] r_run_copy0_j_97;
	reg  signed [31:0] r_run_copy1_j_98;
	reg  signed [31:0] r_run_copy2_j_99;
	reg  signed [31:0] r_run_copy0_j_100;
	reg  signed [31:0] r_run_copy1_j_101;
	reg  signed [31:0] r_run_copy2_j_102;
	reg  signed [31:0] r_run_copy0_j_103;
	reg  signed [31:0] r_run_copy1_j_104;
	reg  signed [31:0] r_run_copy2_j_105;
	reg  signed [31:0] r_run_copy0_j_106;
	reg  signed [31:0] r_run_copy1_j_107;
	reg  signed [31:0] r_run_copy2_j_108;
	reg  signed [31:0] r_run_copy0_j_109;
	reg  signed [31:0] r_run_copy1_j_110;
	reg  signed [31:0] r_run_copy2_j_111;
	reg  signed [31:0] r_run_copy0_j_112;
	reg  signed [31:0] r_run_copy1_j_113;
	reg  signed [31:0] r_run_copy2_j_114;
	reg  signed [31:0] r_run_copy0_j_115;
	reg  signed [31:0] r_run_copy1_j_116;
	reg  signed [31:0] r_run_copy2_j_117;
	reg  signed [31:0] r_run_copy0_j_118;
	reg  signed [31:0] r_run_copy1_j_119;
	reg  signed [31:0] r_run_copy2_j_120;
	reg  signed [31:0] r_run_copy0_j_121;
	reg  signed [31:0] r_run_copy1_j_122;
	reg  signed [31:0] r_run_copy2_j_123;
	reg  signed [31:0] r_run_copy0_j_124;
	reg  signed [31:0] r_run_copy1_j_125;
	reg  signed [31:0] r_run_copy2_j_126;
	reg  signed [31:0] r_run_copy0_j_127;
	reg  signed [31:0] r_run_copy1_j_128;
	reg  signed [31:0] r_run_copy2_j_129;
	reg  signed [31:0] r_run_copy0_j_130;
	reg  signed [31:0] r_run_copy1_j_131;
	reg  signed [31:0] r_run_copy2_j_132;
	reg  signed [31:0] r_run_copy0_j_133;
	reg  signed [31:0] r_run_copy1_j_134;
	reg  signed [31:0] r_run_copy2_j_135;
	reg  signed [31:0] r_run_copy0_j_136;
	reg  signed [31:0] r_run_copy1_j_137;
	reg  signed [31:0] r_run_copy2_j_138;
	reg  signed [31:0] r_run_copy0_j_139;
	reg  signed [31:0] r_run_copy1_j_140;
	reg  signed [31:0] r_run_copy2_j_141;
	reg  signed [31:0] r_run_copy0_j_142;
	reg  signed [31:0] r_run_copy1_j_143;
	reg  signed [31:0] r_run_copy2_j_144;
	reg  signed [31:0] r_run_copy0_j_145;
	reg  signed [31:0] r_run_copy1_j_146;
	reg  signed [31:0] r_run_copy2_j_147;
	reg  signed [31:0] r_run_copy0_j_148;
	reg  signed [31:0] r_run_copy1_j_149;
	reg  signed [31:0] r_run_copy2_j_150;
	reg  signed [31:0] r_run_copy0_j_151;
	reg  signed [31:0] r_run_copy1_j_152;
	reg  signed [31:0] r_run_copy2_j_153;
	reg  signed [31:0] r_run_copy3_j_154;
	reg  signed [31:0] r_run_copy4_j_155;
	reg  signed [31:0] r_run_copy5_j_156;
	reg  signed [31:0] r_run_copy6_j_157;
	reg  signed [31:0] r_run_copy7_j_158;
	reg  signed [31:0] r_run_copy8_j_159;
	reg  signed [31:0] r_run_copy9_j_160;
	reg  signed [31:0] r_run_copy10_j_161;
	reg  signed [31:0] r_run_copy0_j_162;
	reg  signed [31:0] r_run_copy1_j_163;
	reg  signed [31:0] r_run_copy2_j_164;
	reg  signed [31:0] r_run_copy3_j_165;
	reg  signed [31:0] r_run_copy4_j_166;
	reg  signed [31:0] r_run_copy5_j_167;
	reg  signed [31:0] r_run_copy6_j_168;
	reg  signed [31:0] r_run_copy7_j_169;
	reg  signed [31:0] r_run_copy8_j_170;
	reg  signed [31:0] r_run_copy9_j_171;
	reg  signed [31:0] r_run_copy10_j_172;
	reg  signed [31:0] r_run_copy0_j_173;
	reg  signed [31:0] r_run_copy1_j_174;
	reg  signed [31:0] r_run_copy2_j_175;
	reg  signed [31:0] r_run_copy3_j_176;
	reg  signed [31:0] r_run_copy4_j_177;
	reg  signed [31:0] r_run_copy5_j_178;
	reg  signed [31:0] r_run_copy6_j_179;
	reg  signed [31:0] r_run_copy7_j_180;
	reg  signed [31:0] r_run_copy8_j_181;
	reg  signed [31:0] r_run_copy9_j_182;
	reg  signed [31:0] r_run_copy10_j_183;
	reg  signed [31:0] r_run_copy0_j_184;
	reg  signed [31:0] r_run_copy1_j_185;
	reg  signed [31:0] r_run_copy2_j_186;
	reg  signed [31:0] r_run_copy3_j_187;
	reg  signed [31:0] r_run_copy4_j_188;
	reg  signed [31:0] r_run_copy5_j_189;
	reg  signed [31:0] r_run_copy6_j_190;
	reg  signed [31:0] r_run_copy7_j_191;
	reg  signed [31:0] r_run_copy8_j_192;
	reg  signed [31:0] r_run_copy9_j_193;
	reg  signed [31:0] r_run_copy10_j_194;
	reg  signed [31:0] r_run_copy0_j_195;
	reg  signed [31:0] r_run_copy1_j_196;
	reg  signed [31:0] r_run_copy2_j_197;
	reg  signed [31:0] r_run_copy3_j_198;
	reg  signed [31:0] r_run_copy4_j_199;
	reg  signed [31:0] r_run_copy5_j_200;
	reg  signed [31:0] r_run_copy6_j_201;
	reg  signed [31:0] r_run_copy7_j_202;
	reg  signed [31:0] r_run_copy8_j_203;
	reg  signed [31:0] r_run_copy9_j_204;
	reg  signed [31:0] r_run_copy10_j_205;
	reg  signed [31:0] r_run_copy0_j_206;
	reg  signed [31:0] r_run_copy1_j_207;
	reg  signed [31:0] r_run_copy2_j_208;
	reg  signed [31:0] r_run_copy3_j_209;
	reg  signed [31:0] r_run_copy4_j_210;
	reg  signed [31:0] r_run_copy5_j_211;
	reg  signed [31:0] r_run_copy6_j_212;
	reg  signed [31:0] r_run_copy7_j_213;
	reg  signed [31:0] r_run_copy8_j_214;
	reg  signed [31:0] r_run_copy9_j_215;
	reg  signed [31:0] r_run_copy10_j_216;
	reg  signed [31:0] r_run_copy0_j_217;
	reg  signed [31:0] r_run_copy1_j_218;
	reg  signed [31:0] r_run_copy2_j_219;
	reg  signed [31:0] r_run_copy3_j_220;
	reg  signed [31:0] r_run_copy4_j_221;
	reg  signed [31:0] r_run_copy5_j_222;
	reg  signed [31:0] r_run_copy6_j_223;
	reg  signed [31:0] r_run_copy7_j_224;
	reg  signed [31:0] r_run_copy8_j_225;
	reg  signed [31:0] r_run_copy9_j_226;
	reg  signed [31:0] r_run_copy10_j_227;
	reg  signed [31:0] r_run_copy0_j_228;
	reg  signed [31:0] r_run_copy1_j_229;
	reg  signed [31:0] r_run_copy2_j_230;
	reg  signed [31:0] r_run_copy3_j_231;
	reg  signed [31:0] r_run_copy4_j_232;
	reg  signed [31:0] r_run_copy5_j_233;
	reg  signed [31:0] r_run_copy6_j_234;
	reg  signed [31:0] r_run_copy7_j_235;
	reg  signed [31:0] r_run_copy8_j_236;
	reg  signed [31:0] r_run_copy9_j_237;
	reg  signed [31:0] r_run_copy10_j_238;
	reg  signed [31:0] r_run_copy0_j_239;
	reg  signed [31:0] r_run_copy0_j_240;
	reg  signed [31:0] r_run_copy1_j_241;
	reg  signed [31:0] r_run_copy0_j_242;
	reg  signed [31:0] r_run_copy1_j_243;
	reg  signed [31:0] r_run_copy0_j_244;
	reg  signed [31:0] r_run_copy1_j_245;
	reg  signed [31:0] r_run_copy0_j_246;
	reg  signed [31:0] r_run_copy1_j_247;
	reg  signed [31:0] r_run_copy0_j_248;
	reg  signed [31:0] r_run_copy1_j_249;
	reg  signed [31:0] r_run_copy0_j_250;
	reg  signed [31:0] r_run_copy1_j_251;
	reg  signed [31:0] r_run_copy0_j_252;
	reg  signed [31:0] r_run_copy1_j_253;
	reg  signed [31:0] r_run_copy0_j_254;
	reg  signed [31:0] r_run_copy0_j_255;
	reg  signed [31:0] r_run_copy1_j_256;
	reg  signed [31:0] r_run_copy0_j_257;
	reg  signed [31:0] r_run_copy1_j_258;
	reg  signed [31:0] r_run_copy0_j_259;
	reg  signed [31:0] r_run_copy1_j_260;
	reg  signed [31:0] r_run_copy0_j_261;
	reg  signed [31:0] r_run_copy1_j_262;
	reg  signed [31:0] r_run_copy0_j_263;
	reg  signed [31:0] r_run_copy1_j_264;
	reg  signed [31:0] r_run_copy0_j_265;
	reg  signed [31:0] r_run_copy1_j_266;
	reg  signed [31:0] r_run_copy0_j_267;
	reg  signed [31:0] r_run_copy1_j_268;
	reg  signed [31:0] r_run_copy0_j_269;
	reg  signed [31:0] r_run_copy0_j_270;
	reg  signed [31:0] r_run_copy1_j_271;
	reg  signed [31:0] r_run_copy0_j_272;
	reg  signed [31:0] r_run_copy1_j_273;
	reg  signed [31:0] r_run_copy0_j_274;
	reg  signed [31:0] r_run_copy1_j_275;
	reg  signed [31:0] r_run_copy0_j_276;
	reg  signed [31:0] r_run_copy1_j_277;
	reg  signed [31:0] r_run_copy0_j_278;
	reg  signed [31:0] r_run_copy1_j_279;
	reg  signed [31:0] r_run_copy0_j_280;
	reg  signed [31:0] r_run_copy1_j_281;
	reg  signed [31:0] r_run_copy0_j_282;
	reg  signed [31:0] r_run_copy1_j_283;
	reg  signed [31:0] r_run_copy0_j_284;
	reg  signed [31:0] r_run_copy0_j_285;
	reg  signed [31:0] r_run_copy1_j_286;
	reg  signed [31:0] r_run_copy0_j_287;
	reg  signed [31:0] r_run_copy1_j_288;
	reg  signed [31:0] r_run_copy0_j_289;
	reg  signed [31:0] r_run_copy1_j_290;
	reg  signed [31:0] r_run_copy0_j_291;
	reg  signed [31:0] r_run_copy1_j_292;
	reg  signed [31:0] r_run_copy0_j_293;
	reg  signed [31:0] r_run_copy1_j_294;
	reg  signed [31:0] r_run_copy0_j_295;
	reg  signed [31:0] r_run_copy1_j_296;
	reg  signed [31:0] r_run_copy0_j_297;
	reg  signed [31:0] r_run_copy1_j_298;
	reg                r_sub19_run_req;
	wire               w_sub19_run_busy;
	wire signed [11:0] w_sub19_T_addr;
	reg  signed [11:0] r_sub19_T_addr;
	wire        [31:0] w_sub19_T_datain;
	reg         [31:0] r_sub19_T_datain;
	wire        [31:0] w_sub19_T_dataout;
	wire               w_sub19_T_r_w;
	reg                r_sub19_T_r_w;
	wire signed [11:0] w_sub19_U_addr;
	reg  signed [11:0] r_sub19_U_addr;
	wire        [31:0] w_sub19_U_datain;
	reg         [31:0] r_sub19_U_datain;
	wire        [31:0] w_sub19_U_dataout;
	wire               w_sub19_U_r_w;
	reg                r_sub19_U_r_w;
	wire signed [11:0] w_sub19_result_addr;
	reg  signed [11:0] r_sub19_result_addr;
	wire        [31:0] w_sub19_result_datain;
	reg         [31:0] r_sub19_result_datain;
	wire        [31:0] w_sub19_result_dataout;
	wire               w_sub19_result_r_w;
	reg                r_sub19_result_r_w;
	reg                r_sub12_run_req;
	wire               w_sub12_run_busy;
	wire signed [11:0] w_sub12_T_addr;
	reg  signed [11:0] r_sub12_T_addr;
	wire        [31:0] w_sub12_T_datain;
	reg         [31:0] r_sub12_T_datain;
	wire        [31:0] w_sub12_T_dataout;
	wire               w_sub12_T_r_w;
	reg                r_sub12_T_r_w;
	wire signed [11:0] w_sub12_U_addr;
	reg  signed [11:0] r_sub12_U_addr;
	wire        [31:0] w_sub12_U_datain;
	reg         [31:0] r_sub12_U_datain;
	wire        [31:0] w_sub12_U_dataout;
	wire               w_sub12_U_r_w;
	reg                r_sub12_U_r_w;
	wire signed [11:0] w_sub12_result_addr;
	reg  signed [11:0] r_sub12_result_addr;
	wire        [31:0] w_sub12_result_datain;
	reg         [31:0] r_sub12_result_datain;
	wire        [31:0] w_sub12_result_dataout;
	wire               w_sub12_result_r_w;
	reg                r_sub12_result_r_w;
	reg                r_sub11_run_req;
	wire               w_sub11_run_busy;
	wire signed [11:0] w_sub11_T_addr;
	reg  signed [11:0] r_sub11_T_addr;
	wire        [31:0] w_sub11_T_datain;
	reg         [31:0] r_sub11_T_datain;
	wire        [31:0] w_sub11_T_dataout;
	wire               w_sub11_T_r_w;
	reg                r_sub11_T_r_w;
	wire signed [11:0] w_sub11_V_addr;
	reg  signed [11:0] r_sub11_V_addr;
	wire        [31:0] w_sub11_V_datain;
	reg         [31:0] r_sub11_V_datain;
	wire        [31:0] w_sub11_V_dataout;
	wire               w_sub11_V_r_w;
	reg                r_sub11_V_r_w;
	wire signed [11:0] w_sub11_U_addr;
	reg  signed [11:0] r_sub11_U_addr;
	wire        [31:0] w_sub11_U_datain;
	reg         [31:0] r_sub11_U_datain;
	wire        [31:0] w_sub11_U_dataout;
	wire               w_sub11_U_r_w;
	reg                r_sub11_U_r_w;
	wire signed [11:0] w_sub11_result_addr;
	reg  signed [11:0] r_sub11_result_addr;
	wire        [31:0] w_sub11_result_datain;
	reg         [31:0] r_sub11_result_datain;
	wire        [31:0] w_sub11_result_dataout;
	wire               w_sub11_result_r_w;
	reg                r_sub11_result_r_w;
	reg                r_sub14_run_req;
	wire               w_sub14_run_busy;
	wire signed [11:0] w_sub14_T_addr;
	reg  signed [11:0] r_sub14_T_addr;
	wire        [31:0] w_sub14_T_datain;
	reg         [31:0] r_sub14_T_datain;
	wire        [31:0] w_sub14_T_dataout;
	wire               w_sub14_T_r_w;
	reg                r_sub14_T_r_w;
	wire signed [11:0] w_sub14_U_addr;
	reg  signed [11:0] r_sub14_U_addr;
	wire        [31:0] w_sub14_U_datain;
	reg         [31:0] r_sub14_U_datain;
	wire        [31:0] w_sub14_U_dataout;
	wire               w_sub14_U_r_w;
	reg                r_sub14_U_r_w;
	wire signed [11:0] w_sub14_result_addr;
	reg  signed [11:0] r_sub14_result_addr;
	wire        [31:0] w_sub14_result_datain;
	reg         [31:0] r_sub14_result_datain;
	wire        [31:0] w_sub14_result_dataout;
	wire               w_sub14_result_r_w;
	reg                r_sub14_result_r_w;
	reg                r_sub13_run_req;
	wire               w_sub13_run_busy;
	wire signed [11:0] w_sub13_T_addr;
	reg  signed [11:0] r_sub13_T_addr;
	wire        [31:0] w_sub13_T_datain;
	reg         [31:0] r_sub13_T_datain;
	wire        [31:0] w_sub13_T_dataout;
	wire               w_sub13_T_r_w;
	reg                r_sub13_T_r_w;
	wire signed [11:0] w_sub13_U_addr;
	reg  signed [11:0] r_sub13_U_addr;
	wire        [31:0] w_sub13_U_datain;
	reg         [31:0] r_sub13_U_datain;
	wire        [31:0] w_sub13_U_dataout;
	wire               w_sub13_U_r_w;
	reg                r_sub13_U_r_w;
	wire signed [11:0] w_sub13_result_addr;
	reg  signed [11:0] r_sub13_result_addr;
	wire        [31:0] w_sub13_result_datain;
	reg         [31:0] r_sub13_result_datain;
	wire        [31:0] w_sub13_result_dataout;
	wire               w_sub13_result_r_w;
	reg                r_sub13_result_r_w;
	reg                r_sub16_run_req;
	wire               w_sub16_run_busy;
	wire signed [11:0] w_sub16_T_addr;
	reg  signed [11:0] r_sub16_T_addr;
	wire        [31:0] w_sub16_T_datain;
	reg         [31:0] r_sub16_T_datain;
	wire        [31:0] w_sub16_T_dataout;
	wire               w_sub16_T_r_w;
	reg                r_sub16_T_r_w;
	wire signed [11:0] w_sub16_U_addr;
	reg  signed [11:0] r_sub16_U_addr;
	wire        [31:0] w_sub16_U_datain;
	reg         [31:0] r_sub16_U_datain;
	wire        [31:0] w_sub16_U_dataout;
	wire               w_sub16_U_r_w;
	reg                r_sub16_U_r_w;
	wire signed [11:0] w_sub16_result_addr;
	reg  signed [11:0] r_sub16_result_addr;
	wire        [31:0] w_sub16_result_datain;
	reg         [31:0] r_sub16_result_datain;
	wire        [31:0] w_sub16_result_dataout;
	wire               w_sub16_result_r_w;
	reg                r_sub16_result_r_w;
	reg                r_sub15_run_req;
	wire               w_sub15_run_busy;
	wire signed [11:0] w_sub15_T_addr;
	reg  signed [11:0] r_sub15_T_addr;
	wire        [31:0] w_sub15_T_datain;
	reg         [31:0] r_sub15_T_datain;
	wire        [31:0] w_sub15_T_dataout;
	wire               w_sub15_T_r_w;
	reg                r_sub15_T_r_w;
	wire signed [11:0] w_sub15_U_addr;
	reg  signed [11:0] r_sub15_U_addr;
	wire        [31:0] w_sub15_U_datain;
	reg         [31:0] r_sub15_U_datain;
	wire        [31:0] w_sub15_U_dataout;
	wire               w_sub15_U_r_w;
	reg                r_sub15_U_r_w;
	wire signed [11:0] w_sub15_result_addr;
	reg  signed [11:0] r_sub15_result_addr;
	wire        [31:0] w_sub15_result_datain;
	reg         [31:0] r_sub15_result_datain;
	wire        [31:0] w_sub15_result_dataout;
	wire               w_sub15_result_r_w;
	reg                r_sub15_result_r_w;
	reg                r_sub18_run_req;
	wire               w_sub18_run_busy;
	wire signed [11:0] w_sub18_T_addr;
	reg  signed [11:0] r_sub18_T_addr;
	wire        [31:0] w_sub18_T_datain;
	reg         [31:0] r_sub18_T_datain;
	wire        [31:0] w_sub18_T_dataout;
	wire               w_sub18_T_r_w;
	reg                r_sub18_T_r_w;
	wire signed [11:0] w_sub18_U_addr;
	reg  signed [11:0] r_sub18_U_addr;
	wire        [31:0] w_sub18_U_datain;
	reg         [31:0] r_sub18_U_datain;
	wire        [31:0] w_sub18_U_dataout;
	wire               w_sub18_U_r_w;
	reg                r_sub18_U_r_w;
	wire signed [11:0] w_sub18_result_addr;
	reg  signed [11:0] r_sub18_result_addr;
	wire        [31:0] w_sub18_result_datain;
	reg         [31:0] r_sub18_result_datain;
	wire        [31:0] w_sub18_result_dataout;
	wire               w_sub18_result_r_w;
	reg                r_sub18_result_r_w;
	reg                r_sub17_run_req;
	wire               w_sub17_run_busy;
	wire signed [11:0] w_sub17_T_addr;
	reg  signed [11:0] r_sub17_T_addr;
	wire        [31:0] w_sub17_T_datain;
	reg         [31:0] r_sub17_T_datain;
	wire        [31:0] w_sub17_T_dataout;
	wire               w_sub17_T_r_w;
	reg                r_sub17_T_r_w;
	wire signed [11:0] w_sub17_U_addr;
	reg  signed [11:0] r_sub17_U_addr;
	wire        [31:0] w_sub17_U_datain;
	reg         [31:0] r_sub17_U_datain;
	wire        [31:0] w_sub17_U_dataout;
	wire               w_sub17_U_r_w;
	reg                r_sub17_U_r_w;
	wire signed [11:0] w_sub17_result_addr;
	reg  signed [11:0] r_sub17_result_addr;
	wire        [31:0] w_sub17_result_datain;
	reg         [31:0] r_sub17_result_datain;
	wire        [31:0] w_sub17_result_dataout;
	wire               w_sub17_result_r_w;
	reg                r_sub17_result_r_w;
	reg                r_sub20_run_req;
	wire               w_sub20_run_busy;
	wire signed [11:0] w_sub20_T_addr;
	reg  signed [11:0] r_sub20_T_addr;
	wire        [31:0] w_sub20_T_datain;
	reg         [31:0] r_sub20_T_datain;
	wire        [31:0] w_sub20_T_dataout;
	wire               w_sub20_T_r_w;
	reg                r_sub20_T_r_w;
	wire signed [11:0] w_sub20_U_addr;
	reg  signed [11:0] r_sub20_U_addr;
	wire        [31:0] w_sub20_U_datain;
	reg         [31:0] r_sub20_U_datain;
	wire        [31:0] w_sub20_U_dataout;
	wire               w_sub20_U_r_w;
	reg                r_sub20_U_r_w;
	wire signed [11:0] w_sub20_result_addr;
	reg  signed [11:0] r_sub20_result_addr;
	wire        [31:0] w_sub20_result_datain;
	reg         [31:0] r_sub20_result_datain;
	wire        [31:0] w_sub20_result_dataout;
	wire               w_sub20_result_r_w;
	reg                r_sub20_result_r_w;
	reg                r_sub21_run_req;
	wire               w_sub21_run_busy;
	wire signed [11:0] w_sub21_T_addr;
	reg  signed [11:0] r_sub21_T_addr;
	wire        [31:0] w_sub21_T_datain;
	reg         [31:0] r_sub21_T_datain;
	wire        [31:0] w_sub21_T_dataout;
	wire               w_sub21_T_r_w;
	reg                r_sub21_T_r_w;
	wire signed [11:0] w_sub21_U_addr;
	reg  signed [11:0] r_sub21_U_addr;
	wire        [31:0] w_sub21_U_datain;
	reg         [31:0] r_sub21_U_datain;
	wire        [31:0] w_sub21_U_dataout;
	wire               w_sub21_U_r_w;
	reg                r_sub21_U_r_w;
	wire signed [11:0] w_sub21_result_addr;
	reg  signed [11:0] r_sub21_result_addr;
	wire        [31:0] w_sub21_result_datain;
	reg         [31:0] r_sub21_result_datain;
	wire        [31:0] w_sub21_result_dataout;
	wire               w_sub21_result_r_w;
	reg                r_sub21_result_r_w;
	reg                r_sub28_run_req;
	wire               w_sub28_run_busy;
	wire signed [11:0] w_sub28_T_addr;
	reg  signed [11:0] r_sub28_T_addr;
	wire        [31:0] w_sub28_T_datain;
	reg         [31:0] r_sub28_T_datain;
	wire        [31:0] w_sub28_T_dataout;
	wire               w_sub28_T_r_w;
	reg                r_sub28_T_r_w;
	wire signed [11:0] w_sub28_U_addr;
	reg  signed [11:0] r_sub28_U_addr;
	wire        [31:0] w_sub28_U_datain;
	reg         [31:0] r_sub28_U_datain;
	wire        [31:0] w_sub28_U_dataout;
	wire               w_sub28_U_r_w;
	reg                r_sub28_U_r_w;
	wire signed [11:0] w_sub28_result_addr;
	reg  signed [11:0] r_sub28_result_addr;
	wire        [31:0] w_sub28_result_datain;
	reg         [31:0] r_sub28_result_datain;
	wire        [31:0] w_sub28_result_dataout;
	wire               w_sub28_result_r_w;
	reg                r_sub28_result_r_w;
	reg                r_sub29_run_req;
	wire               w_sub29_run_busy;
	wire signed [11:0] w_sub29_T_addr;
	reg  signed [11:0] r_sub29_T_addr;
	wire        [31:0] w_sub29_T_datain;
	reg         [31:0] r_sub29_T_datain;
	wire        [31:0] w_sub29_T_dataout;
	wire               w_sub29_T_r_w;
	reg                r_sub29_T_r_w;
	wire signed [11:0] w_sub29_U_addr;
	reg  signed [11:0] r_sub29_U_addr;
	wire        [31:0] w_sub29_U_datain;
	reg         [31:0] r_sub29_U_datain;
	wire        [31:0] w_sub29_U_dataout;
	wire               w_sub29_U_r_w;
	reg                r_sub29_U_r_w;
	wire signed [11:0] w_sub29_result_addr;
	reg  signed [11:0] r_sub29_result_addr;
	wire        [31:0] w_sub29_result_datain;
	reg         [31:0] r_sub29_result_datain;
	wire        [31:0] w_sub29_result_dataout;
	wire               w_sub29_result_r_w;
	reg                r_sub29_result_r_w;
	reg                r_sub26_run_req;
	wire               w_sub26_run_busy;
	wire signed [11:0] w_sub26_T_addr;
	reg  signed [11:0] r_sub26_T_addr;
	wire        [31:0] w_sub26_T_datain;
	reg         [31:0] r_sub26_T_datain;
	wire        [31:0] w_sub26_T_dataout;
	wire               w_sub26_T_r_w;
	reg                r_sub26_T_r_w;
	wire signed [11:0] w_sub26_U_addr;
	reg  signed [11:0] r_sub26_U_addr;
	wire        [31:0] w_sub26_U_datain;
	reg         [31:0] r_sub26_U_datain;
	wire        [31:0] w_sub26_U_dataout;
	wire               w_sub26_U_r_w;
	reg                r_sub26_U_r_w;
	wire signed [11:0] w_sub26_result_addr;
	reg  signed [11:0] r_sub26_result_addr;
	wire        [31:0] w_sub26_result_datain;
	reg         [31:0] r_sub26_result_datain;
	wire        [31:0] w_sub26_result_dataout;
	wire               w_sub26_result_r_w;
	reg                r_sub26_result_r_w;
	reg                r_sub09_run_req;
	wire               w_sub09_run_busy;
	wire signed [11:0] w_sub09_T_addr;
	reg  signed [11:0] r_sub09_T_addr;
	wire        [31:0] w_sub09_T_datain;
	reg         [31:0] r_sub09_T_datain;
	wire        [31:0] w_sub09_T_dataout;
	wire               w_sub09_T_r_w;
	reg                r_sub09_T_r_w;
	wire signed [11:0] w_sub09_U_addr;
	reg  signed [11:0] r_sub09_U_addr;
	wire        [31:0] w_sub09_U_datain;
	reg         [31:0] r_sub09_U_datain;
	wire        [31:0] w_sub09_U_dataout;
	wire               w_sub09_U_r_w;
	reg                r_sub09_U_r_w;
	wire signed [11:0] w_sub09_result_addr;
	reg  signed [11:0] r_sub09_result_addr;
	wire        [31:0] w_sub09_result_datain;
	reg         [31:0] r_sub09_result_datain;
	wire        [31:0] w_sub09_result_dataout;
	wire               w_sub09_result_r_w;
	reg                r_sub09_result_r_w;
	reg                r_sub27_run_req;
	wire               w_sub27_run_busy;
	wire signed [11:0] w_sub27_T_addr;
	reg  signed [11:0] r_sub27_T_addr;
	wire        [31:0] w_sub27_T_datain;
	reg         [31:0] r_sub27_T_datain;
	wire        [31:0] w_sub27_T_dataout;
	wire               w_sub27_T_r_w;
	reg                r_sub27_T_r_w;
	wire signed [11:0] w_sub27_U_addr;
	reg  signed [11:0] r_sub27_U_addr;
	wire        [31:0] w_sub27_U_datain;
	reg         [31:0] r_sub27_U_datain;
	wire        [31:0] w_sub27_U_dataout;
	wire               w_sub27_U_r_w;
	reg                r_sub27_U_r_w;
	wire signed [11:0] w_sub27_result_addr;
	reg  signed [11:0] r_sub27_result_addr;
	wire        [31:0] w_sub27_result_datain;
	reg         [31:0] r_sub27_result_datain;
	wire        [31:0] w_sub27_result_dataout;
	wire               w_sub27_result_r_w;
	reg                r_sub27_result_r_w;
	reg                r_sub08_run_req;
	wire               w_sub08_run_busy;
	wire signed [11:0] w_sub08_T_addr;
	reg  signed [11:0] r_sub08_T_addr;
	wire        [31:0] w_sub08_T_datain;
	reg         [31:0] r_sub08_T_datain;
	wire        [31:0] w_sub08_T_dataout;
	wire               w_sub08_T_r_w;
	reg                r_sub08_T_r_w;
	wire signed [11:0] w_sub08_U_addr;
	reg  signed [11:0] r_sub08_U_addr;
	wire        [31:0] w_sub08_U_datain;
	reg         [31:0] r_sub08_U_datain;
	wire        [31:0] w_sub08_U_dataout;
	wire               w_sub08_U_r_w;
	reg                r_sub08_U_r_w;
	wire signed [11:0] w_sub08_result_addr;
	reg  signed [11:0] r_sub08_result_addr;
	wire        [31:0] w_sub08_result_datain;
	reg         [31:0] r_sub08_result_datain;
	wire        [31:0] w_sub08_result_dataout;
	wire               w_sub08_result_r_w;
	reg                r_sub08_result_r_w;
	reg                r_sub24_run_req;
	wire               w_sub24_run_busy;
	wire signed [11:0] w_sub24_T_addr;
	reg  signed [11:0] r_sub24_T_addr;
	wire        [31:0] w_sub24_T_datain;
	reg         [31:0] r_sub24_T_datain;
	wire        [31:0] w_sub24_T_dataout;
	wire               w_sub24_T_r_w;
	reg                r_sub24_T_r_w;
	wire signed [11:0] w_sub24_U_addr;
	reg  signed [11:0] r_sub24_U_addr;
	wire        [31:0] w_sub24_U_datain;
	reg         [31:0] r_sub24_U_datain;
	wire        [31:0] w_sub24_U_dataout;
	wire               w_sub24_U_r_w;
	reg                r_sub24_U_r_w;
	wire signed [11:0] w_sub24_result_addr;
	reg  signed [11:0] r_sub24_result_addr;
	wire        [31:0] w_sub24_result_datain;
	reg         [31:0] r_sub24_result_datain;
	wire        [31:0] w_sub24_result_dataout;
	wire               w_sub24_result_r_w;
	reg                r_sub24_result_r_w;
	reg                r_sub25_run_req;
	wire               w_sub25_run_busy;
	wire signed [11:0] w_sub25_T_addr;
	reg  signed [11:0] r_sub25_T_addr;
	wire        [31:0] w_sub25_T_datain;
	reg         [31:0] r_sub25_T_datain;
	wire        [31:0] w_sub25_T_dataout;
	wire               w_sub25_T_r_w;
	reg                r_sub25_T_r_w;
	wire signed [11:0] w_sub25_U_addr;
	reg  signed [11:0] r_sub25_U_addr;
	wire        [31:0] w_sub25_U_datain;
	reg         [31:0] r_sub25_U_datain;
	wire        [31:0] w_sub25_U_dataout;
	wire               w_sub25_U_r_w;
	reg                r_sub25_U_r_w;
	wire signed [11:0] w_sub25_result_addr;
	reg  signed [11:0] r_sub25_result_addr;
	wire        [31:0] w_sub25_result_datain;
	reg         [31:0] r_sub25_result_datain;
	wire        [31:0] w_sub25_result_dataout;
	wire               w_sub25_result_r_w;
	reg                r_sub25_result_r_w;
	reg                r_sub22_run_req;
	wire               w_sub22_run_busy;
	wire signed [11:0] w_sub22_T_addr;
	reg  signed [11:0] r_sub22_T_addr;
	wire        [31:0] w_sub22_T_datain;
	reg         [31:0] r_sub22_T_datain;
	wire        [31:0] w_sub22_T_dataout;
	wire               w_sub22_T_r_w;
	reg                r_sub22_T_r_w;
	wire signed [11:0] w_sub22_U_addr;
	reg  signed [11:0] r_sub22_U_addr;
	wire        [31:0] w_sub22_U_datain;
	reg         [31:0] r_sub22_U_datain;
	wire        [31:0] w_sub22_U_dataout;
	wire               w_sub22_U_r_w;
	reg                r_sub22_U_r_w;
	wire signed [11:0] w_sub22_result_addr;
	reg  signed [11:0] r_sub22_result_addr;
	wire        [31:0] w_sub22_result_datain;
	reg         [31:0] r_sub22_result_datain;
	wire        [31:0] w_sub22_result_dataout;
	wire               w_sub22_result_r_w;
	reg                r_sub22_result_r_w;
	reg                r_sub23_run_req;
	wire               w_sub23_run_busy;
	wire signed [11:0] w_sub23_T_addr;
	reg  signed [11:0] r_sub23_T_addr;
	wire        [31:0] w_sub23_T_datain;
	reg         [31:0] r_sub23_T_datain;
	wire        [31:0] w_sub23_T_dataout;
	wire               w_sub23_T_r_w;
	reg                r_sub23_T_r_w;
	wire signed [11:0] w_sub23_U_addr;
	reg  signed [11:0] r_sub23_U_addr;
	wire        [31:0] w_sub23_U_datain;
	reg         [31:0] r_sub23_U_datain;
	wire        [31:0] w_sub23_U_dataout;
	wire               w_sub23_U_r_w;
	reg                r_sub23_U_r_w;
	wire signed [11:0] w_sub23_result_addr;
	reg  signed [11:0] r_sub23_result_addr;
	wire        [31:0] w_sub23_result_datain;
	reg         [31:0] r_sub23_result_datain;
	wire        [31:0] w_sub23_result_dataout;
	wire               w_sub23_result_r_w;
	reg                r_sub23_result_r_w;
	reg                r_sub03_run_req;
	wire               w_sub03_run_busy;
	wire signed [11:0] w_sub03_T_addr;
	reg  signed [11:0] r_sub03_T_addr;
	wire        [31:0] w_sub03_T_datain;
	reg         [31:0] r_sub03_T_datain;
	wire        [31:0] w_sub03_T_dataout;
	wire               w_sub03_T_r_w;
	reg                r_sub03_T_r_w;
	wire signed [11:0] w_sub03_U_addr;
	reg  signed [11:0] r_sub03_U_addr;
	wire        [31:0] w_sub03_U_datain;
	reg         [31:0] r_sub03_U_datain;
	wire        [31:0] w_sub03_U_dataout;
	wire               w_sub03_U_r_w;
	reg                r_sub03_U_r_w;
	wire signed [11:0] w_sub03_result_addr;
	reg  signed [11:0] r_sub03_result_addr;
	wire        [31:0] w_sub03_result_datain;
	reg         [31:0] r_sub03_result_datain;
	wire        [31:0] w_sub03_result_dataout;
	wire               w_sub03_result_r_w;
	reg                r_sub03_result_r_w;
	reg                r_sub02_run_req;
	wire               w_sub02_run_busy;
	wire signed [11:0] w_sub02_T_addr;
	reg  signed [11:0] r_sub02_T_addr;
	wire        [31:0] w_sub02_T_datain;
	reg         [31:0] r_sub02_T_datain;
	wire        [31:0] w_sub02_T_dataout;
	wire               w_sub02_T_r_w;
	reg                r_sub02_T_r_w;
	wire signed [11:0] w_sub02_U_addr;
	reg  signed [11:0] r_sub02_U_addr;
	wire        [31:0] w_sub02_U_datain;
	reg         [31:0] r_sub02_U_datain;
	wire        [31:0] w_sub02_U_dataout;
	wire               w_sub02_U_r_w;
	reg                r_sub02_U_r_w;
	wire signed [11:0] w_sub02_result_addr;
	reg  signed [11:0] r_sub02_result_addr;
	wire        [31:0] w_sub02_result_datain;
	reg         [31:0] r_sub02_result_datain;
	wire        [31:0] w_sub02_result_dataout;
	wire               w_sub02_result_r_w;
	reg                r_sub02_result_r_w;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [11:0] w_sub01_T_addr;
	reg  signed [11:0] r_sub01_T_addr;
	wire        [31:0] w_sub01_T_datain;
	reg         [31:0] r_sub01_T_datain;
	wire        [31:0] w_sub01_T_dataout;
	wire               w_sub01_T_r_w;
	reg                r_sub01_T_r_w;
	wire signed [11:0] w_sub01_U_addr;
	reg  signed [11:0] r_sub01_U_addr;
	wire        [31:0] w_sub01_U_datain;
	reg         [31:0] r_sub01_U_datain;
	wire        [31:0] w_sub01_U_dataout;
	wire               w_sub01_U_r_w;
	reg                r_sub01_U_r_w;
	wire signed [11:0] w_sub01_result_addr;
	reg  signed [11:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [11:0] w_sub00_T_addr;
	reg  signed [11:0] r_sub00_T_addr;
	wire        [31:0] w_sub00_T_datain;
	reg         [31:0] r_sub00_T_datain;
	wire        [31:0] w_sub00_T_dataout;
	wire               w_sub00_T_r_w;
	reg                r_sub00_T_r_w;
	wire signed [11:0] w_sub00_U_addr;
	reg  signed [11:0] r_sub00_U_addr;
	wire        [31:0] w_sub00_U_datain;
	reg         [31:0] r_sub00_U_datain;
	wire        [31:0] w_sub00_U_dataout;
	wire               w_sub00_U_r_w;
	reg                r_sub00_U_r_w;
	wire signed [11:0] w_sub00_result_addr;
	reg  signed [11:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	reg                r_sub07_run_req;
	wire               w_sub07_run_busy;
	wire signed [11:0] w_sub07_T_addr;
	reg  signed [11:0] r_sub07_T_addr;
	wire        [31:0] w_sub07_T_datain;
	reg         [31:0] r_sub07_T_datain;
	wire        [31:0] w_sub07_T_dataout;
	wire               w_sub07_T_r_w;
	reg                r_sub07_T_r_w;
	wire signed [11:0] w_sub07_U_addr;
	reg  signed [11:0] r_sub07_U_addr;
	wire        [31:0] w_sub07_U_datain;
	reg         [31:0] r_sub07_U_datain;
	wire        [31:0] w_sub07_U_dataout;
	wire               w_sub07_U_r_w;
	reg                r_sub07_U_r_w;
	wire signed [11:0] w_sub07_result_addr;
	reg  signed [11:0] r_sub07_result_addr;
	wire        [31:0] w_sub07_result_datain;
	reg         [31:0] r_sub07_result_datain;
	wire        [31:0] w_sub07_result_dataout;
	wire               w_sub07_result_r_w;
	reg                r_sub07_result_r_w;
	reg                r_sub06_run_req;
	wire               w_sub06_run_busy;
	wire signed [11:0] w_sub06_T_addr;
	reg  signed [11:0] r_sub06_T_addr;
	wire        [31:0] w_sub06_T_datain;
	reg         [31:0] r_sub06_T_datain;
	wire        [31:0] w_sub06_T_dataout;
	wire               w_sub06_T_r_w;
	reg                r_sub06_T_r_w;
	wire signed [11:0] w_sub06_U_addr;
	reg  signed [11:0] r_sub06_U_addr;
	wire        [31:0] w_sub06_U_datain;
	reg         [31:0] r_sub06_U_datain;
	wire        [31:0] w_sub06_U_dataout;
	wire               w_sub06_U_r_w;
	reg                r_sub06_U_r_w;
	wire signed [11:0] w_sub06_result_addr;
	reg  signed [11:0] r_sub06_result_addr;
	wire        [31:0] w_sub06_result_datain;
	reg         [31:0] r_sub06_result_datain;
	wire        [31:0] w_sub06_result_dataout;
	wire               w_sub06_result_r_w;
	reg                r_sub06_result_r_w;
	reg                r_sub05_run_req;
	wire               w_sub05_run_busy;
	wire signed [11:0] w_sub05_T_addr;
	reg  signed [11:0] r_sub05_T_addr;
	wire        [31:0] w_sub05_T_datain;
	reg         [31:0] r_sub05_T_datain;
	wire        [31:0] w_sub05_T_dataout;
	wire               w_sub05_T_r_w;
	reg                r_sub05_T_r_w;
	wire signed [11:0] w_sub05_U_addr;
	reg  signed [11:0] r_sub05_U_addr;
	wire        [31:0] w_sub05_U_datain;
	reg         [31:0] r_sub05_U_datain;
	wire        [31:0] w_sub05_U_dataout;
	wire               w_sub05_U_r_w;
	reg                r_sub05_U_r_w;
	wire signed [11:0] w_sub05_result_addr;
	reg  signed [11:0] r_sub05_result_addr;
	wire        [31:0] w_sub05_result_datain;
	reg         [31:0] r_sub05_result_datain;
	wire        [31:0] w_sub05_result_dataout;
	wire               w_sub05_result_r_w;
	reg                r_sub05_result_r_w;
	reg                r_sub04_run_req;
	wire               w_sub04_run_busy;
	wire signed [11:0] w_sub04_T_addr;
	reg  signed [11:0] r_sub04_T_addr;
	wire        [31:0] w_sub04_T_datain;
	reg         [31:0] r_sub04_T_datain;
	wire        [31:0] w_sub04_T_dataout;
	wire               w_sub04_T_r_w;
	reg                r_sub04_T_r_w;
	wire signed [11:0] w_sub04_U_addr;
	reg  signed [11:0] r_sub04_U_addr;
	wire        [31:0] w_sub04_U_datain;
	reg         [31:0] r_sub04_U_datain;
	wire        [31:0] w_sub04_U_dataout;
	wire               w_sub04_U_r_w;
	reg                r_sub04_U_r_w;
	wire signed [11:0] w_sub04_result_addr;
	reg  signed [11:0] r_sub04_result_addr;
	wire        [31:0] w_sub04_result_datain;
	reg         [31:0] r_sub04_result_datain;
	wire        [31:0] w_sub04_result_dataout;
	wire               w_sub04_result_r_w;
	reg                r_sub04_result_r_w;
	reg                r_sub10_run_req;
	wire               w_sub10_run_busy;
	wire signed [11:0] w_sub10_T_addr;
	reg  signed [11:0] r_sub10_T_addr;
	wire        [31:0] w_sub10_T_datain;
	reg         [31:0] r_sub10_T_datain;
	wire        [31:0] w_sub10_T_dataout;
	wire               w_sub10_T_r_w;
	reg                r_sub10_T_r_w;
	wire signed [11:0] w_sub10_U_addr;
	reg  signed [11:0] r_sub10_U_addr;
	wire        [31:0] w_sub10_U_datain;
	reg         [31:0] r_sub10_U_datain;
	wire        [31:0] w_sub10_U_dataout;
	wire               w_sub10_U_r_w;
	reg                r_sub10_U_r_w;
	wire signed [11:0] w_sub10_result_addr;
	reg  signed [11:0] r_sub10_result_addr;
	wire        [31:0] w_sub10_result_datain;
	reg         [31:0] r_sub10_result_datain;
	wire        [31:0] w_sub10_result_dataout;
	wire               w_sub10_result_r_w;
	reg                r_sub10_result_r_w;
	reg                r_sub31_run_req;
	wire               w_sub31_run_busy;
	wire signed [11:0] w_sub31_T_addr;
	reg  signed [11:0] r_sub31_T_addr;
	wire        [31:0] w_sub31_T_datain;
	reg         [31:0] r_sub31_T_datain;
	wire        [31:0] w_sub31_T_dataout;
	wire               w_sub31_T_r_w;
	reg                r_sub31_T_r_w;
	wire signed [11:0] w_sub31_U_addr;
	reg  signed [11:0] r_sub31_U_addr;
	wire        [31:0] w_sub31_U_datain;
	reg         [31:0] r_sub31_U_datain;
	wire        [31:0] w_sub31_U_dataout;
	wire               w_sub31_U_r_w;
	reg                r_sub31_U_r_w;
	wire signed [11:0] w_sub31_result_addr;
	reg  signed [11:0] r_sub31_result_addr;
	wire        [31:0] w_sub31_result_datain;
	reg         [31:0] r_sub31_result_datain;
	wire        [31:0] w_sub31_result_dataout;
	wire               w_sub31_result_r_w;
	reg                r_sub31_result_r_w;
	reg                r_sub30_run_req;
	wire               w_sub30_run_busy;
	wire signed [11:0] w_sub30_T_addr;
	reg  signed [11:0] r_sub30_T_addr;
	wire        [31:0] w_sub30_T_datain;
	reg         [31:0] r_sub30_T_datain;
	wire        [31:0] w_sub30_T_dataout;
	wire               w_sub30_T_r_w;
	reg                r_sub30_T_r_w;
	wire signed [11:0] w_sub30_U_addr;
	reg  signed [11:0] r_sub30_U_addr;
	wire        [31:0] w_sub30_U_datain;
	reg         [31:0] r_sub30_U_datain;
	wire        [31:0] w_sub30_U_dataout;
	wire               w_sub30_U_r_w;
	reg                r_sub30_U_r_w;
	wire signed [11:0] w_sub30_result_addr;
	reg  signed [11:0] r_sub30_result_addr;
	wire        [31:0] w_sub30_result_datain;
	reg         [31:0] r_sub30_result_datain;
	wire        [31:0] w_sub30_result_dataout;
	wire               w_sub30_result_r_w;
	reg                r_sub30_result_r_w;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg         [31:0] r_sys_tmp4_float;
	reg         [31:0] r_sys_tmp5_float;
	reg         [31:0] r_sys_tmp6_float;
	reg         [31:0] r_sys_tmp7_float;
	wire signed [31:0] w_sys_tmp1;
	wire signed [31:0] w_sys_tmp3;
	wire        [31:0] w_sys_tmp5;
	wire        [31:0] w_sys_tmp6;
	wire        [31:0] w_sys_tmp7;
	wire        [31:0] w_sys_tmp8;
	wire        [31:0] w_sys_tmp9;
	wire        [31:0] w_sys_tmp10;
	wire        [31:0] w_sys_tmp11;
	wire               w_sys_tmp12;
	wire               w_sys_tmp13;
	wire signed [31:0] w_sys_tmp14;
	wire               w_sys_tmp15;
	wire               w_sys_tmp16;
	wire        [31:0] w_sys_tmp18;
	wire        [31:0] w_sys_tmp19;
	wire signed [31:0] w_sys_tmp20;
	wire signed [31:0] w_sys_tmp22;
	wire signed [31:0] w_sys_tmp23;
	wire signed [31:0] w_sys_tmp24;
	wire        [31:0] w_sys_tmp25;
	wire signed [31:0] w_sys_tmp27;
	wire signed [31:0] w_sys_tmp28;
	wire signed [31:0] w_sys_tmp32;
	wire signed [31:0] w_sys_tmp33;
	wire        [31:0] w_sys_tmp36;
	wire        [31:0] w_sys_tmp37;
	wire        [31:0] w_sys_tmp38;
	wire signed [31:0] w_sys_tmp40;
	wire signed [31:0] w_sys_tmp41;
	wire signed [31:0] w_sys_tmp42;
	wire        [31:0] w_sys_tmp110;
	wire               w_sys_tmp184;
	wire               w_sys_tmp185;
	wire signed [31:0] w_sys_tmp186;
	wire signed [31:0] w_sys_tmp189;
	wire signed [31:0] w_sys_tmp190;
	wire        [31:0] w_sys_tmp191;
	wire signed [31:0] w_sys_tmp193;
	wire signed [31:0] w_sys_tmp194;
	wire        [31:0] w_sys_tmp196;
	wire signed [31:0] w_sys_tmp197;
	wire signed [31:0] w_sys_tmp198;
	wire signed [31:0] w_sys_tmp199;
	wire signed [31:0] w_sys_tmp201;
	wire               w_sys_tmp202;
	wire               w_sys_tmp203;
	wire signed [31:0] w_sys_tmp204;
	wire signed [31:0] w_sys_tmp207;
	wire signed [31:0] w_sys_tmp208;
	wire signed [31:0] w_sys_tmp209;
	wire        [31:0] w_sys_tmp210;
	wire signed [31:0] w_sys_tmp212;
	wire signed [31:0] w_sys_tmp213;
	wire signed [31:0] w_sys_tmp216;
	wire signed [31:0] w_sys_tmp217;
	wire signed [31:0] w_sys_tmp290;
	wire signed [31:0] w_sys_tmp291;
	wire               w_sys_tmp292;
	wire               w_sys_tmp293;
	wire signed [31:0] w_sys_tmp294;
	wire signed [31:0] w_sys_tmp295;
	wire signed [31:0] w_sys_tmp298;
	wire signed [31:0] w_sys_tmp299;
	wire signed [31:0] w_sys_tmp300;
	wire        [31:0] w_sys_tmp301;
	wire signed [31:0] w_sys_tmp302;
	wire               w_sys_tmp339;
	wire               w_sys_tmp340;
	wire signed [31:0] w_sys_tmp341;
	wire signed [31:0] w_sys_tmp342;
	wire               w_sys_tmp343;
	wire               w_sys_tmp344;
	wire signed [31:0] w_sys_tmp345;
	wire signed [31:0] w_sys_tmp348;
	wire signed [31:0] w_sys_tmp349;
	wire signed [31:0] w_sys_tmp350;
	wire        [31:0] w_sys_tmp351;
	wire signed [31:0] w_sys_tmp352;
	wire signed [31:0] w_sys_tmp353;
	wire signed [31:0] w_sys_tmp356;
	wire signed [31:0] w_sys_tmp357;
	wire        [31:0] w_sys_tmp359;
	wire signed [31:0] w_sys_tmp360;
	wire signed [31:0] w_sys_tmp361;
	wire signed [31:0] w_sys_tmp363;
	wire signed [31:0] w_sys_tmp364;
	wire signed [31:0] w_sys_tmp365;
	wire signed [31:0] w_sys_tmp366;
	wire signed [31:0] w_sys_tmp487;
	wire               w_sys_tmp488;
	wire               w_sys_tmp489;
	wire signed [31:0] w_sys_tmp490;
	wire signed [31:0] w_sys_tmp493;
	wire signed [31:0] w_sys_tmp494;
	wire signed [31:0] w_sys_tmp495;
	wire        [31:0] w_sys_tmp496;
	wire signed [31:0] w_sys_tmp497;
	wire signed [31:0] w_sys_tmp498;
	wire signed [31:0] w_sys_tmp501;
	wire signed [31:0] w_sys_tmp502;
	wire        [31:0] w_sys_tmp504;
	wire signed [31:0] w_sys_tmp505;
	wire signed [31:0] w_sys_tmp506;
	wire signed [31:0] w_sys_tmp508;
	wire signed [31:0] w_sys_tmp509;
	wire signed [31:0] w_sys_tmp510;
	wire signed [31:0] w_sys_tmp511;
	wire signed [31:0] w_sys_tmp632;
	wire               w_sys_tmp633;
	wire               w_sys_tmp634;
	wire signed [31:0] w_sys_tmp635;
	wire signed [31:0] w_sys_tmp638;
	wire signed [31:0] w_sys_tmp639;
	wire signed [31:0] w_sys_tmp640;
	wire        [31:0] w_sys_tmp641;
	wire signed [31:0] w_sys_tmp642;
	wire signed [31:0] w_sys_tmp643;
	wire signed [31:0] w_sys_tmp646;
	wire signed [31:0] w_sys_tmp647;
	wire        [31:0] w_sys_tmp649;
	wire signed [31:0] w_sys_tmp650;
	wire signed [31:0] w_sys_tmp651;
	wire signed [31:0] w_sys_tmp653;
	wire signed [31:0] w_sys_tmp654;
	wire signed [31:0] w_sys_tmp655;
	wire signed [31:0] w_sys_tmp656;
	wire signed [31:0] w_sys_tmp777;
	wire               w_sys_tmp778;
	wire               w_sys_tmp779;
	wire signed [31:0] w_sys_tmp780;
	wire signed [31:0] w_sys_tmp783;
	wire signed [31:0] w_sys_tmp784;
	wire signed [31:0] w_sys_tmp785;
	wire        [31:0] w_sys_tmp786;
	wire signed [31:0] w_sys_tmp787;
	wire signed [31:0] w_sys_tmp788;
	wire signed [31:0] w_sys_tmp791;
	wire signed [31:0] w_sys_tmp792;
	wire        [31:0] w_sys_tmp794;
	wire signed [31:0] w_sys_tmp795;
	wire signed [31:0] w_sys_tmp796;
	wire signed [31:0] w_sys_tmp798;
	wire signed [31:0] w_sys_tmp799;
	wire signed [31:0] w_sys_tmp800;
	wire signed [31:0] w_sys_tmp801;
	wire signed [31:0] w_sys_tmp922;
	wire               w_sys_tmp923;
	wire               w_sys_tmp924;
	wire signed [31:0] w_sys_tmp925;
	wire signed [31:0] w_sys_tmp928;
	wire signed [31:0] w_sys_tmp929;
	wire signed [31:0] w_sys_tmp930;
	wire        [31:0] w_sys_tmp931;
	wire signed [31:0] w_sys_tmp932;
	wire signed [31:0] w_sys_tmp933;
	wire signed [31:0] w_sys_tmp936;
	wire signed [31:0] w_sys_tmp937;
	wire        [31:0] w_sys_tmp939;
	wire signed [31:0] w_sys_tmp940;
	wire signed [31:0] w_sys_tmp941;
	wire signed [31:0] w_sys_tmp943;
	wire signed [31:0] w_sys_tmp944;
	wire signed [31:0] w_sys_tmp945;
	wire signed [31:0] w_sys_tmp946;
	wire signed [31:0] w_sys_tmp1067;
	wire               w_sys_tmp1068;
	wire               w_sys_tmp1069;
	wire signed [31:0] w_sys_tmp1070;
	wire signed [31:0] w_sys_tmp1073;
	wire signed [31:0] w_sys_tmp1074;
	wire signed [31:0] w_sys_tmp1075;
	wire        [31:0] w_sys_tmp1076;
	wire signed [31:0] w_sys_tmp1077;
	wire signed [31:0] w_sys_tmp1078;
	wire signed [31:0] w_sys_tmp1081;
	wire signed [31:0] w_sys_tmp1082;
	wire        [31:0] w_sys_tmp1084;
	wire signed [31:0] w_sys_tmp1085;
	wire signed [31:0] w_sys_tmp1086;
	wire signed [31:0] w_sys_tmp1088;
	wire signed [31:0] w_sys_tmp1089;
	wire signed [31:0] w_sys_tmp1090;
	wire signed [31:0] w_sys_tmp1091;
	wire signed [31:0] w_sys_tmp1212;
	wire               w_sys_tmp1213;
	wire               w_sys_tmp1214;
	wire signed [31:0] w_sys_tmp1215;
	wire signed [31:0] w_sys_tmp1218;
	wire signed [31:0] w_sys_tmp1219;
	wire signed [31:0] w_sys_tmp1220;
	wire        [31:0] w_sys_tmp1221;
	wire signed [31:0] w_sys_tmp1222;
	wire signed [31:0] w_sys_tmp1223;
	wire signed [31:0] w_sys_tmp1226;
	wire signed [31:0] w_sys_tmp1227;
	wire        [31:0] w_sys_tmp1229;
	wire signed [31:0] w_sys_tmp1230;
	wire signed [31:0] w_sys_tmp1231;
	wire signed [31:0] w_sys_tmp1233;
	wire signed [31:0] w_sys_tmp1234;
	wire signed [31:0] w_sys_tmp1235;
	wire signed [31:0] w_sys_tmp1236;
	wire signed [31:0] w_sys_tmp1357;
	wire               w_sys_tmp1358;
	wire               w_sys_tmp1359;
	wire signed [31:0] w_sys_tmp1360;
	wire signed [31:0] w_sys_tmp1363;
	wire signed [31:0] w_sys_tmp1364;
	wire signed [31:0] w_sys_tmp1365;
	wire        [31:0] w_sys_tmp1366;
	wire signed [31:0] w_sys_tmp1367;
	wire signed [31:0] w_sys_tmp1368;
	wire signed [31:0] w_sys_tmp1371;
	wire signed [31:0] w_sys_tmp1372;
	wire        [31:0] w_sys_tmp1374;
	wire signed [31:0] w_sys_tmp1375;
	wire signed [31:0] w_sys_tmp1376;
	wire signed [31:0] w_sys_tmp1378;
	wire signed [31:0] w_sys_tmp1379;
	wire signed [31:0] w_sys_tmp1380;
	wire signed [31:0] w_sys_tmp1381;
	wire               w_sys_tmp1502;
	wire               w_sys_tmp1503;
	wire signed [31:0] w_sys_tmp1504;
	wire signed [31:0] w_sys_tmp1505;
	wire               w_sys_tmp1506;
	wire               w_sys_tmp1507;
	wire signed [31:0] w_sys_tmp1508;
	wire signed [31:0] w_sys_tmp1511;
	wire signed [31:0] w_sys_tmp1512;
	wire signed [31:0] w_sys_tmp1513;
	wire        [31:0] w_sys_tmp1514;
	wire signed [31:0] w_sys_tmp1515;
	wire signed [31:0] w_sys_tmp1516;
	wire signed [31:0] w_sys_tmp1519;
	wire signed [31:0] w_sys_tmp1520;
	wire        [31:0] w_sys_tmp1522;
	wire signed [31:0] w_sys_tmp1523;
	wire signed [31:0] w_sys_tmp1524;
	wire signed [31:0] w_sys_tmp1526;
	wire signed [31:0] w_sys_tmp1527;
	wire signed [31:0] w_sys_tmp1528;
	wire signed [31:0] w_sys_tmp1529;
	wire signed [31:0] w_sys_tmp1650;
	wire               w_sys_tmp1651;
	wire               w_sys_tmp1652;
	wire signed [31:0] w_sys_tmp1653;
	wire signed [31:0] w_sys_tmp1656;
	wire signed [31:0] w_sys_tmp1657;
	wire signed [31:0] w_sys_tmp1658;
	wire        [31:0] w_sys_tmp1659;
	wire signed [31:0] w_sys_tmp1660;
	wire signed [31:0] w_sys_tmp1661;
	wire signed [31:0] w_sys_tmp1664;
	wire signed [31:0] w_sys_tmp1665;
	wire        [31:0] w_sys_tmp1667;
	wire signed [31:0] w_sys_tmp1668;
	wire signed [31:0] w_sys_tmp1669;
	wire signed [31:0] w_sys_tmp1671;
	wire signed [31:0] w_sys_tmp1672;
	wire signed [31:0] w_sys_tmp1673;
	wire signed [31:0] w_sys_tmp1674;
	wire signed [31:0] w_sys_tmp1795;
	wire               w_sys_tmp1796;
	wire               w_sys_tmp1797;
	wire signed [31:0] w_sys_tmp1798;
	wire signed [31:0] w_sys_tmp1801;
	wire signed [31:0] w_sys_tmp1802;
	wire signed [31:0] w_sys_tmp1803;
	wire        [31:0] w_sys_tmp1804;
	wire signed [31:0] w_sys_tmp1805;
	wire signed [31:0] w_sys_tmp1806;
	wire signed [31:0] w_sys_tmp1809;
	wire signed [31:0] w_sys_tmp1810;
	wire        [31:0] w_sys_tmp1812;
	wire signed [31:0] w_sys_tmp1813;
	wire signed [31:0] w_sys_tmp1814;
	wire signed [31:0] w_sys_tmp1816;
	wire signed [31:0] w_sys_tmp1817;
	wire signed [31:0] w_sys_tmp1818;
	wire signed [31:0] w_sys_tmp1819;
	wire signed [31:0] w_sys_tmp1940;
	wire               w_sys_tmp1941;
	wire               w_sys_tmp1942;
	wire signed [31:0] w_sys_tmp1943;
	wire signed [31:0] w_sys_tmp1946;
	wire signed [31:0] w_sys_tmp1947;
	wire signed [31:0] w_sys_tmp1948;
	wire        [31:0] w_sys_tmp1949;
	wire signed [31:0] w_sys_tmp1950;
	wire signed [31:0] w_sys_tmp1951;
	wire signed [31:0] w_sys_tmp1954;
	wire signed [31:0] w_sys_tmp1955;
	wire        [31:0] w_sys_tmp1957;
	wire signed [31:0] w_sys_tmp1958;
	wire signed [31:0] w_sys_tmp1959;
	wire signed [31:0] w_sys_tmp1961;
	wire signed [31:0] w_sys_tmp1962;
	wire signed [31:0] w_sys_tmp1963;
	wire signed [31:0] w_sys_tmp1964;
	wire signed [31:0] w_sys_tmp2085;
	wire               w_sys_tmp2086;
	wire               w_sys_tmp2087;
	wire signed [31:0] w_sys_tmp2088;
	wire signed [31:0] w_sys_tmp2091;
	wire signed [31:0] w_sys_tmp2092;
	wire signed [31:0] w_sys_tmp2093;
	wire        [31:0] w_sys_tmp2094;
	wire signed [31:0] w_sys_tmp2095;
	wire signed [31:0] w_sys_tmp2096;
	wire signed [31:0] w_sys_tmp2099;
	wire signed [31:0] w_sys_tmp2100;
	wire        [31:0] w_sys_tmp2102;
	wire signed [31:0] w_sys_tmp2103;
	wire signed [31:0] w_sys_tmp2104;
	wire signed [31:0] w_sys_tmp2106;
	wire signed [31:0] w_sys_tmp2107;
	wire signed [31:0] w_sys_tmp2108;
	wire signed [31:0] w_sys_tmp2109;
	wire signed [31:0] w_sys_tmp2230;
	wire               w_sys_tmp2231;
	wire               w_sys_tmp2232;
	wire signed [31:0] w_sys_tmp2233;
	wire signed [31:0] w_sys_tmp2236;
	wire signed [31:0] w_sys_tmp2237;
	wire signed [31:0] w_sys_tmp2238;
	wire        [31:0] w_sys_tmp2239;
	wire signed [31:0] w_sys_tmp2240;
	wire signed [31:0] w_sys_tmp2241;
	wire signed [31:0] w_sys_tmp2244;
	wire signed [31:0] w_sys_tmp2245;
	wire        [31:0] w_sys_tmp2247;
	wire signed [31:0] w_sys_tmp2248;
	wire signed [31:0] w_sys_tmp2249;
	wire signed [31:0] w_sys_tmp2251;
	wire signed [31:0] w_sys_tmp2252;
	wire signed [31:0] w_sys_tmp2253;
	wire signed [31:0] w_sys_tmp2254;
	wire signed [31:0] w_sys_tmp2375;
	wire               w_sys_tmp2376;
	wire               w_sys_tmp2377;
	wire signed [31:0] w_sys_tmp2378;
	wire signed [31:0] w_sys_tmp2381;
	wire signed [31:0] w_sys_tmp2382;
	wire signed [31:0] w_sys_tmp2383;
	wire        [31:0] w_sys_tmp2384;
	wire signed [31:0] w_sys_tmp2385;
	wire signed [31:0] w_sys_tmp2386;
	wire signed [31:0] w_sys_tmp2389;
	wire signed [31:0] w_sys_tmp2390;
	wire        [31:0] w_sys_tmp2392;
	wire signed [31:0] w_sys_tmp2393;
	wire signed [31:0] w_sys_tmp2394;
	wire signed [31:0] w_sys_tmp2396;
	wire signed [31:0] w_sys_tmp2397;
	wire signed [31:0] w_sys_tmp2398;
	wire signed [31:0] w_sys_tmp2399;
	wire signed [31:0] w_sys_tmp2520;
	wire               w_sys_tmp2521;
	wire               w_sys_tmp2522;
	wire signed [31:0] w_sys_tmp2523;
	wire signed [31:0] w_sys_tmp2526;
	wire signed [31:0] w_sys_tmp2527;
	wire signed [31:0] w_sys_tmp2528;
	wire        [31:0] w_sys_tmp2529;
	wire signed [31:0] w_sys_tmp2530;
	wire signed [31:0] w_sys_tmp2531;
	wire signed [31:0] w_sys_tmp2534;
	wire signed [31:0] w_sys_tmp2535;
	wire        [31:0] w_sys_tmp2537;
	wire signed [31:0] w_sys_tmp2538;
	wire signed [31:0] w_sys_tmp2539;
	wire signed [31:0] w_sys_tmp2541;
	wire signed [31:0] w_sys_tmp2542;
	wire signed [31:0] w_sys_tmp2543;
	wire signed [31:0] w_sys_tmp2544;
	wire               w_sys_tmp2665;
	wire               w_sys_tmp2666;
	wire signed [31:0] w_sys_tmp2667;
	wire signed [31:0] w_sys_tmp2668;
	wire               w_sys_tmp2669;
	wire               w_sys_tmp2670;
	wire signed [31:0] w_sys_tmp2671;
	wire signed [31:0] w_sys_tmp2674;
	wire signed [31:0] w_sys_tmp2675;
	wire signed [31:0] w_sys_tmp2676;
	wire        [31:0] w_sys_tmp2677;
	wire signed [31:0] w_sys_tmp2678;
	wire signed [31:0] w_sys_tmp2679;
	wire signed [31:0] w_sys_tmp2682;
	wire signed [31:0] w_sys_tmp2683;
	wire        [31:0] w_sys_tmp2685;
	wire signed [31:0] w_sys_tmp2686;
	wire signed [31:0] w_sys_tmp2687;
	wire signed [31:0] w_sys_tmp2689;
	wire signed [31:0] w_sys_tmp2690;
	wire signed [31:0] w_sys_tmp2691;
	wire signed [31:0] w_sys_tmp2692;
	wire signed [31:0] w_sys_tmp2813;
	wire               w_sys_tmp2814;
	wire               w_sys_tmp2815;
	wire signed [31:0] w_sys_tmp2816;
	wire signed [31:0] w_sys_tmp2819;
	wire signed [31:0] w_sys_tmp2820;
	wire signed [31:0] w_sys_tmp2821;
	wire        [31:0] w_sys_tmp2822;
	wire signed [31:0] w_sys_tmp2823;
	wire signed [31:0] w_sys_tmp2824;
	wire signed [31:0] w_sys_tmp2827;
	wire signed [31:0] w_sys_tmp2828;
	wire        [31:0] w_sys_tmp2830;
	wire signed [31:0] w_sys_tmp2831;
	wire signed [31:0] w_sys_tmp2832;
	wire signed [31:0] w_sys_tmp2834;
	wire signed [31:0] w_sys_tmp2835;
	wire signed [31:0] w_sys_tmp2836;
	wire signed [31:0] w_sys_tmp2837;
	wire signed [31:0] w_sys_tmp2958;
	wire               w_sys_tmp2959;
	wire               w_sys_tmp2960;
	wire signed [31:0] w_sys_tmp2961;
	wire signed [31:0] w_sys_tmp2964;
	wire signed [31:0] w_sys_tmp2965;
	wire signed [31:0] w_sys_tmp2966;
	wire        [31:0] w_sys_tmp2967;
	wire signed [31:0] w_sys_tmp2968;
	wire signed [31:0] w_sys_tmp2969;
	wire signed [31:0] w_sys_tmp2972;
	wire signed [31:0] w_sys_tmp2973;
	wire        [31:0] w_sys_tmp2975;
	wire signed [31:0] w_sys_tmp2976;
	wire signed [31:0] w_sys_tmp2977;
	wire signed [31:0] w_sys_tmp2979;
	wire signed [31:0] w_sys_tmp2980;
	wire signed [31:0] w_sys_tmp2981;
	wire signed [31:0] w_sys_tmp2982;
	wire signed [31:0] w_sys_tmp3103;
	wire               w_sys_tmp3104;
	wire               w_sys_tmp3105;
	wire signed [31:0] w_sys_tmp3106;
	wire signed [31:0] w_sys_tmp3109;
	wire signed [31:0] w_sys_tmp3110;
	wire signed [31:0] w_sys_tmp3111;
	wire        [31:0] w_sys_tmp3112;
	wire signed [31:0] w_sys_tmp3113;
	wire signed [31:0] w_sys_tmp3114;
	wire signed [31:0] w_sys_tmp3117;
	wire signed [31:0] w_sys_tmp3118;
	wire        [31:0] w_sys_tmp3120;
	wire signed [31:0] w_sys_tmp3121;
	wire signed [31:0] w_sys_tmp3122;
	wire signed [31:0] w_sys_tmp3124;
	wire signed [31:0] w_sys_tmp3125;
	wire signed [31:0] w_sys_tmp3126;
	wire signed [31:0] w_sys_tmp3127;
	wire signed [31:0] w_sys_tmp3248;
	wire               w_sys_tmp3249;
	wire               w_sys_tmp3250;
	wire signed [31:0] w_sys_tmp3251;
	wire signed [31:0] w_sys_tmp3254;
	wire signed [31:0] w_sys_tmp3255;
	wire signed [31:0] w_sys_tmp3256;
	wire        [31:0] w_sys_tmp3257;
	wire signed [31:0] w_sys_tmp3258;
	wire signed [31:0] w_sys_tmp3259;
	wire signed [31:0] w_sys_tmp3262;
	wire signed [31:0] w_sys_tmp3263;
	wire        [31:0] w_sys_tmp3265;
	wire signed [31:0] w_sys_tmp3266;
	wire signed [31:0] w_sys_tmp3267;
	wire signed [31:0] w_sys_tmp3269;
	wire signed [31:0] w_sys_tmp3270;
	wire signed [31:0] w_sys_tmp3271;
	wire signed [31:0] w_sys_tmp3272;
	wire signed [31:0] w_sys_tmp3393;
	wire               w_sys_tmp3394;
	wire               w_sys_tmp3395;
	wire signed [31:0] w_sys_tmp3396;
	wire signed [31:0] w_sys_tmp3399;
	wire signed [31:0] w_sys_tmp3400;
	wire signed [31:0] w_sys_tmp3401;
	wire        [31:0] w_sys_tmp3402;
	wire signed [31:0] w_sys_tmp3403;
	wire signed [31:0] w_sys_tmp3404;
	wire signed [31:0] w_sys_tmp3407;
	wire signed [31:0] w_sys_tmp3408;
	wire        [31:0] w_sys_tmp3410;
	wire signed [31:0] w_sys_tmp3411;
	wire signed [31:0] w_sys_tmp3412;
	wire signed [31:0] w_sys_tmp3414;
	wire signed [31:0] w_sys_tmp3415;
	wire signed [31:0] w_sys_tmp3416;
	wire signed [31:0] w_sys_tmp3417;
	wire signed [31:0] w_sys_tmp3538;
	wire               w_sys_tmp3539;
	wire               w_sys_tmp3540;
	wire signed [31:0] w_sys_tmp3541;
	wire signed [31:0] w_sys_tmp3544;
	wire signed [31:0] w_sys_tmp3545;
	wire signed [31:0] w_sys_tmp3546;
	wire        [31:0] w_sys_tmp3547;
	wire signed [31:0] w_sys_tmp3548;
	wire signed [31:0] w_sys_tmp3549;
	wire signed [31:0] w_sys_tmp3552;
	wire signed [31:0] w_sys_tmp3553;
	wire        [31:0] w_sys_tmp3555;
	wire signed [31:0] w_sys_tmp3556;
	wire signed [31:0] w_sys_tmp3557;
	wire signed [31:0] w_sys_tmp3559;
	wire signed [31:0] w_sys_tmp3560;
	wire signed [31:0] w_sys_tmp3561;
	wire signed [31:0] w_sys_tmp3562;
	wire signed [31:0] w_sys_tmp3683;
	wire               w_sys_tmp3684;
	wire               w_sys_tmp3685;
	wire signed [31:0] w_sys_tmp3686;
	wire signed [31:0] w_sys_tmp3689;
	wire signed [31:0] w_sys_tmp3690;
	wire signed [31:0] w_sys_tmp3691;
	wire        [31:0] w_sys_tmp3692;
	wire signed [31:0] w_sys_tmp3693;
	wire signed [31:0] w_sys_tmp3694;
	wire signed [31:0] w_sys_tmp3697;
	wire signed [31:0] w_sys_tmp3698;
	wire        [31:0] w_sys_tmp3700;
	wire signed [31:0] w_sys_tmp3701;
	wire signed [31:0] w_sys_tmp3702;
	wire signed [31:0] w_sys_tmp3704;
	wire signed [31:0] w_sys_tmp3705;
	wire signed [31:0] w_sys_tmp3706;
	wire signed [31:0] w_sys_tmp3707;
	wire               w_sys_tmp3828;
	wire               w_sys_tmp3829;
	wire signed [31:0] w_sys_tmp3830;
	wire signed [31:0] w_sys_tmp3831;
	wire               w_sys_tmp3832;
	wire               w_sys_tmp3833;
	wire signed [31:0] w_sys_tmp3834;
	wire signed [31:0] w_sys_tmp3837;
	wire signed [31:0] w_sys_tmp3838;
	wire signed [31:0] w_sys_tmp3839;
	wire        [31:0] w_sys_tmp3840;
	wire signed [31:0] w_sys_tmp3841;
	wire signed [31:0] w_sys_tmp3842;
	wire signed [31:0] w_sys_tmp3845;
	wire signed [31:0] w_sys_tmp3846;
	wire        [31:0] w_sys_tmp3848;
	wire signed [31:0] w_sys_tmp3849;
	wire signed [31:0] w_sys_tmp3850;
	wire signed [31:0] w_sys_tmp3852;
	wire signed [31:0] w_sys_tmp3853;
	wire signed [31:0] w_sys_tmp3854;
	wire signed [31:0] w_sys_tmp3855;
	wire signed [31:0] w_sys_tmp3976;
	wire               w_sys_tmp3977;
	wire               w_sys_tmp3978;
	wire signed [31:0] w_sys_tmp3979;
	wire signed [31:0] w_sys_tmp3982;
	wire signed [31:0] w_sys_tmp3983;
	wire signed [31:0] w_sys_tmp3984;
	wire        [31:0] w_sys_tmp3985;
	wire signed [31:0] w_sys_tmp3986;
	wire signed [31:0] w_sys_tmp3987;
	wire signed [31:0] w_sys_tmp3990;
	wire signed [31:0] w_sys_tmp3991;
	wire        [31:0] w_sys_tmp3993;
	wire signed [31:0] w_sys_tmp3994;
	wire signed [31:0] w_sys_tmp3995;
	wire signed [31:0] w_sys_tmp3997;
	wire signed [31:0] w_sys_tmp3998;
	wire signed [31:0] w_sys_tmp3999;
	wire signed [31:0] w_sys_tmp4000;
	wire signed [31:0] w_sys_tmp4121;
	wire               w_sys_tmp4122;
	wire               w_sys_tmp4123;
	wire signed [31:0] w_sys_tmp4124;
	wire signed [31:0] w_sys_tmp4127;
	wire signed [31:0] w_sys_tmp4128;
	wire signed [31:0] w_sys_tmp4129;
	wire        [31:0] w_sys_tmp4130;
	wire signed [31:0] w_sys_tmp4131;
	wire signed [31:0] w_sys_tmp4132;
	wire signed [31:0] w_sys_tmp4135;
	wire signed [31:0] w_sys_tmp4136;
	wire        [31:0] w_sys_tmp4138;
	wire signed [31:0] w_sys_tmp4139;
	wire signed [31:0] w_sys_tmp4140;
	wire signed [31:0] w_sys_tmp4142;
	wire signed [31:0] w_sys_tmp4143;
	wire signed [31:0] w_sys_tmp4144;
	wire signed [31:0] w_sys_tmp4145;
	wire signed [31:0] w_sys_tmp4266;
	wire               w_sys_tmp4267;
	wire               w_sys_tmp4268;
	wire signed [31:0] w_sys_tmp4269;
	wire signed [31:0] w_sys_tmp4272;
	wire signed [31:0] w_sys_tmp4273;
	wire signed [31:0] w_sys_tmp4274;
	wire        [31:0] w_sys_tmp4275;
	wire signed [31:0] w_sys_tmp4276;
	wire signed [31:0] w_sys_tmp4277;
	wire signed [31:0] w_sys_tmp4280;
	wire signed [31:0] w_sys_tmp4281;
	wire        [31:0] w_sys_tmp4283;
	wire signed [31:0] w_sys_tmp4284;
	wire signed [31:0] w_sys_tmp4285;
	wire signed [31:0] w_sys_tmp4287;
	wire signed [31:0] w_sys_tmp4288;
	wire signed [31:0] w_sys_tmp4289;
	wire signed [31:0] w_sys_tmp4290;
	wire signed [31:0] w_sys_tmp4411;
	wire               w_sys_tmp4412;
	wire               w_sys_tmp4413;
	wire signed [31:0] w_sys_tmp4414;
	wire signed [31:0] w_sys_tmp4417;
	wire signed [31:0] w_sys_tmp4418;
	wire signed [31:0] w_sys_tmp4419;
	wire        [31:0] w_sys_tmp4420;
	wire signed [31:0] w_sys_tmp4421;
	wire signed [31:0] w_sys_tmp4422;
	wire signed [31:0] w_sys_tmp4425;
	wire signed [31:0] w_sys_tmp4426;
	wire        [31:0] w_sys_tmp4428;
	wire signed [31:0] w_sys_tmp4429;
	wire signed [31:0] w_sys_tmp4430;
	wire signed [31:0] w_sys_tmp4432;
	wire signed [31:0] w_sys_tmp4433;
	wire signed [31:0] w_sys_tmp4434;
	wire signed [31:0] w_sys_tmp4435;
	wire signed [31:0] w_sys_tmp4556;
	wire               w_sys_tmp4557;
	wire               w_sys_tmp4558;
	wire signed [31:0] w_sys_tmp4559;
	wire signed [31:0] w_sys_tmp4562;
	wire signed [31:0] w_sys_tmp4563;
	wire signed [31:0] w_sys_tmp4564;
	wire        [31:0] w_sys_tmp4565;
	wire signed [31:0] w_sys_tmp4566;
	wire signed [31:0] w_sys_tmp4567;
	wire signed [31:0] w_sys_tmp4570;
	wire signed [31:0] w_sys_tmp4571;
	wire        [31:0] w_sys_tmp4573;
	wire signed [31:0] w_sys_tmp4574;
	wire signed [31:0] w_sys_tmp4575;
	wire signed [31:0] w_sys_tmp4577;
	wire signed [31:0] w_sys_tmp4578;
	wire signed [31:0] w_sys_tmp4579;
	wire signed [31:0] w_sys_tmp4580;
	wire signed [31:0] w_sys_tmp4701;
	wire               w_sys_tmp4702;
	wire               w_sys_tmp4703;
	wire signed [31:0] w_sys_tmp4704;
	wire signed [31:0] w_sys_tmp4707;
	wire signed [31:0] w_sys_tmp4708;
	wire signed [31:0] w_sys_tmp4709;
	wire        [31:0] w_sys_tmp4710;
	wire signed [31:0] w_sys_tmp4711;
	wire signed [31:0] w_sys_tmp4712;
	wire signed [31:0] w_sys_tmp4715;
	wire signed [31:0] w_sys_tmp4716;
	wire        [31:0] w_sys_tmp4718;
	wire signed [31:0] w_sys_tmp4719;
	wire signed [31:0] w_sys_tmp4720;
	wire signed [31:0] w_sys_tmp4722;
	wire signed [31:0] w_sys_tmp4723;
	wire signed [31:0] w_sys_tmp4724;
	wire signed [31:0] w_sys_tmp4725;
	wire signed [31:0] w_sys_tmp4846;
	wire               w_sys_tmp4847;
	wire               w_sys_tmp4848;
	wire signed [31:0] w_sys_tmp4849;
	wire signed [31:0] w_sys_tmp4852;
	wire signed [31:0] w_sys_tmp4853;
	wire signed [31:0] w_sys_tmp4854;
	wire        [31:0] w_sys_tmp4855;
	wire signed [31:0] w_sys_tmp4856;
	wire signed [31:0] w_sys_tmp4857;
	wire signed [31:0] w_sys_tmp4860;
	wire signed [31:0] w_sys_tmp4861;
	wire        [31:0] w_sys_tmp4863;
	wire signed [31:0] w_sys_tmp4864;
	wire signed [31:0] w_sys_tmp4865;
	wire signed [31:0] w_sys_tmp4867;
	wire signed [31:0] w_sys_tmp4868;
	wire signed [31:0] w_sys_tmp4869;
	wire signed [31:0] w_sys_tmp4870;
	wire               w_sys_tmp4991;
	wire               w_sys_tmp4992;
	wire signed [31:0] w_sys_tmp4993;
	wire signed [31:0] w_sys_tmp4994;
	wire               w_sys_tmp4995;
	wire               w_sys_tmp4996;
	wire signed [31:0] w_sys_tmp4997;
	wire signed [31:0] w_sys_tmp5000;
	wire signed [31:0] w_sys_tmp5001;
	wire        [31:0] w_sys_tmp5002;
	wire signed [31:0] w_sys_tmp5003;
	wire signed [31:0] w_sys_tmp5004;
	wire signed [31:0] w_sys_tmp5006;
	wire signed [31:0] w_sys_tmp5007;
	wire        [31:0] w_sys_tmp5008;
	wire signed [31:0] w_sys_tmp5009;
	wire signed [31:0] w_sys_tmp5010;
	wire signed [31:0] w_sys_tmp5012;
	wire signed [31:0] w_sys_tmp5013;
	wire        [31:0] w_sys_tmp5030;
	wire        [31:0] w_sys_tmp5041;
	wire        [31:0] w_sys_tmp5052;
	wire        [31:0] w_sys_tmp5063;
	wire        [31:0] w_sys_tmp5074;
	wire signed [31:0] w_sys_tmp5077;
	wire signed [31:0] w_sys_tmp5078;
	wire               w_sys_tmp5079;
	wire               w_sys_tmp5080;
	wire signed [31:0] w_sys_tmp5081;
	wire signed [31:0] w_sys_tmp5084;
	wire signed [31:0] w_sys_tmp5085;
	wire        [31:0] w_sys_tmp5086;
	wire signed [31:0] w_sys_tmp5087;
	wire signed [31:0] w_sys_tmp5088;
	wire signed [31:0] w_sys_tmp5090;
	wire signed [31:0] w_sys_tmp5091;
	wire        [31:0] w_sys_tmp5092;
	wire signed [31:0] w_sys_tmp5093;
	wire signed [31:0] w_sys_tmp5094;
	wire signed [31:0] w_sys_tmp5096;
	wire signed [31:0] w_sys_tmp5097;
	wire        [31:0] w_sys_tmp5114;
	wire        [31:0] w_sys_tmp5125;
	wire        [31:0] w_sys_tmp5136;
	wire        [31:0] w_sys_tmp5147;
	wire        [31:0] w_sys_tmp5158;
	wire signed [31:0] w_sys_tmp5161;
	wire signed [31:0] w_sys_tmp5162;
	wire               w_sys_tmp5163;
	wire               w_sys_tmp5164;
	wire signed [31:0] w_sys_tmp5165;
	wire signed [31:0] w_sys_tmp5168;
	wire signed [31:0] w_sys_tmp5169;
	wire        [31:0] w_sys_tmp5170;
	wire signed [31:0] w_sys_tmp5171;
	wire signed [31:0] w_sys_tmp5172;
	wire signed [31:0] w_sys_tmp5174;
	wire signed [31:0] w_sys_tmp5175;
	wire        [31:0] w_sys_tmp5176;
	wire signed [31:0] w_sys_tmp5177;
	wire signed [31:0] w_sys_tmp5178;
	wire signed [31:0] w_sys_tmp5180;
	wire signed [31:0] w_sys_tmp5181;
	wire        [31:0] w_sys_tmp5198;
	wire        [31:0] w_sys_tmp5209;
	wire        [31:0] w_sys_tmp5220;
	wire        [31:0] w_sys_tmp5231;
	wire        [31:0] w_sys_tmp5242;
	wire signed [31:0] w_sys_tmp5245;
	wire signed [31:0] w_sys_tmp5246;
	wire               w_sys_tmp5247;
	wire               w_sys_tmp5248;
	wire signed [31:0] w_sys_tmp5249;
	wire signed [31:0] w_sys_tmp5252;
	wire signed [31:0] w_sys_tmp5253;
	wire        [31:0] w_sys_tmp5254;
	wire signed [31:0] w_sys_tmp5255;
	wire signed [31:0] w_sys_tmp5256;
	wire signed [31:0] w_sys_tmp5258;
	wire signed [31:0] w_sys_tmp5259;
	wire        [31:0] w_sys_tmp5260;
	wire signed [31:0] w_sys_tmp5261;
	wire signed [31:0] w_sys_tmp5262;
	wire signed [31:0] w_sys_tmp5264;
	wire signed [31:0] w_sys_tmp5265;
	wire        [31:0] w_sys_tmp5282;
	wire        [31:0] w_sys_tmp5293;
	wire        [31:0] w_sys_tmp5304;
	wire        [31:0] w_sys_tmp5315;
	wire        [31:0] w_sys_tmp5326;
	wire signed [31:0] w_sys_tmp5329;
	wire               w_sys_tmp5330;
	wire               w_sys_tmp5331;
	wire signed [31:0] w_sys_tmp5332;
	wire signed [31:0] w_sys_tmp5335;
	wire signed [31:0] w_sys_tmp5336;
	wire signed [31:0] w_sys_tmp5337;
	wire signed [31:0] w_sys_tmp5338;
	wire        [31:0] w_sys_tmp5339;
	wire signed [31:0] w_sys_tmp5340;
	wire signed [31:0] w_sys_tmp5341;
	wire signed [31:0] w_sys_tmp5345;
	wire signed [31:0] w_sys_tmp5346;
	wire signed [31:0] w_sys_tmp5348;
	wire        [31:0] w_sys_tmp5349;
	wire signed [31:0] w_sys_tmp5350;
	wire signed [31:0] w_sys_tmp5351;
	wire signed [31:0] w_sys_tmp5355;
	wire signed [31:0] w_sys_tmp5356;
	wire signed [31:0] w_sys_tmp5358;
	wire signed [31:0] w_sys_tmp5359;
	wire signed [31:0] w_sys_tmp5360;
	wire signed [31:0] w_sys_tmp5364;
	wire signed [31:0] w_sys_tmp5365;
	wire signed [31:0] w_sys_tmp5367;
	wire signed [31:0] w_sys_tmp5369;
	wire signed [31:0] w_sys_tmp5370;
	wire signed [31:0] w_sys_tmp5374;
	wire signed [31:0] w_sys_tmp5375;
	wire signed [31:0] w_sys_tmp5377;
	wire signed [31:0] w_sys_tmp5378;
	wire signed [31:0] w_sys_tmp5379;
	wire signed [31:0] w_sys_tmp5383;
	wire signed [31:0] w_sys_tmp5384;
	wire signed [31:0] w_sys_tmp5386;
	wire        [31:0] w_sys_tmp5387;
	wire signed [31:0] w_sys_tmp5388;
	wire signed [31:0] w_sys_tmp5389;
	wire signed [31:0] w_sys_tmp5392;
	wire signed [31:0] w_sys_tmp5393;
	wire signed [31:0] w_sys_tmp5394;
	wire signed [31:0] w_sys_tmp5395;
	wire signed [31:0] w_sys_tmp5396;
	wire signed [31:0] w_sys_tmp5397;
	wire signed [31:0] w_sys_tmp5398;
	wire signed [31:0] w_sys_tmp5399;
	wire signed [31:0] w_sys_tmp5400;
	wire signed [31:0] w_sys_tmp5401;
	wire signed [31:0] w_sys_tmp5402;
	wire signed [31:0] w_sys_tmp5403;
	wire signed [31:0] w_sys_tmp5830;
	wire               w_sys_tmp5831;
	wire               w_sys_tmp5832;
	wire signed [31:0] w_sys_tmp5833;
	wire signed [31:0] w_sys_tmp5836;
	wire signed [31:0] w_sys_tmp5837;
	wire signed [31:0] w_sys_tmp5838;
	wire signed [31:0] w_sys_tmp5839;
	wire        [31:0] w_sys_tmp5840;
	wire signed [31:0] w_sys_tmp5841;
	wire signed [31:0] w_sys_tmp5842;
	wire signed [31:0] w_sys_tmp5846;
	wire signed [31:0] w_sys_tmp5847;
	wire signed [31:0] w_sys_tmp5849;
	wire        [31:0] w_sys_tmp5850;
	wire signed [31:0] w_sys_tmp5851;
	wire signed [31:0] w_sys_tmp5852;
	wire signed [31:0] w_sys_tmp5856;
	wire signed [31:0] w_sys_tmp5857;
	wire signed [31:0] w_sys_tmp5859;
	wire signed [31:0] w_sys_tmp5860;
	wire signed [31:0] w_sys_tmp5861;
	wire signed [31:0] w_sys_tmp5865;
	wire signed [31:0] w_sys_tmp5866;
	wire signed [31:0] w_sys_tmp5868;
	wire signed [31:0] w_sys_tmp5870;
	wire signed [31:0] w_sys_tmp5871;
	wire signed [31:0] w_sys_tmp5875;
	wire signed [31:0] w_sys_tmp5876;
	wire signed [31:0] w_sys_tmp5878;
	wire signed [31:0] w_sys_tmp5879;
	wire signed [31:0] w_sys_tmp5880;
	wire signed [31:0] w_sys_tmp5884;
	wire signed [31:0] w_sys_tmp5885;
	wire signed [31:0] w_sys_tmp5887;
	wire        [31:0] w_sys_tmp5888;
	wire signed [31:0] w_sys_tmp5889;
	wire signed [31:0] w_sys_tmp5890;
	wire signed [31:0] w_sys_tmp5893;
	wire signed [31:0] w_sys_tmp5894;
	wire signed [31:0] w_sys_tmp5895;
	wire signed [31:0] w_sys_tmp5896;
	wire signed [31:0] w_sys_tmp5897;
	wire signed [31:0] w_sys_tmp5898;
	wire signed [31:0] w_sys_tmp5899;
	wire signed [31:0] w_sys_tmp5900;
	wire signed [31:0] w_sys_tmp5901;
	wire signed [31:0] w_sys_tmp5902;
	wire signed [31:0] w_sys_tmp5903;
	wire signed [31:0] w_sys_tmp5904;
	wire signed [31:0] w_sys_tmp6331;
	wire               w_sys_tmp6332;
	wire               w_sys_tmp6333;
	wire signed [31:0] w_sys_tmp6334;
	wire signed [31:0] w_sys_tmp6337;
	wire signed [31:0] w_sys_tmp6338;
	wire signed [31:0] w_sys_tmp6339;
	wire signed [31:0] w_sys_tmp6340;
	wire        [31:0] w_sys_tmp6341;
	wire signed [31:0] w_sys_tmp6342;
	wire signed [31:0] w_sys_tmp6343;
	wire signed [31:0] w_sys_tmp6347;
	wire signed [31:0] w_sys_tmp6348;
	wire signed [31:0] w_sys_tmp6350;
	wire        [31:0] w_sys_tmp6351;
	wire signed [31:0] w_sys_tmp6352;
	wire signed [31:0] w_sys_tmp6353;
	wire signed [31:0] w_sys_tmp6357;
	wire signed [31:0] w_sys_tmp6358;
	wire signed [31:0] w_sys_tmp6360;
	wire signed [31:0] w_sys_tmp6361;
	wire signed [31:0] w_sys_tmp6362;
	wire signed [31:0] w_sys_tmp6366;
	wire signed [31:0] w_sys_tmp6367;
	wire signed [31:0] w_sys_tmp6369;
	wire signed [31:0] w_sys_tmp6371;
	wire signed [31:0] w_sys_tmp6372;
	wire signed [31:0] w_sys_tmp6376;
	wire signed [31:0] w_sys_tmp6377;
	wire signed [31:0] w_sys_tmp6379;
	wire signed [31:0] w_sys_tmp6380;
	wire signed [31:0] w_sys_tmp6381;
	wire signed [31:0] w_sys_tmp6385;
	wire signed [31:0] w_sys_tmp6386;
	wire signed [31:0] w_sys_tmp6388;
	wire        [31:0] w_sys_tmp6389;
	wire signed [31:0] w_sys_tmp6390;
	wire signed [31:0] w_sys_tmp6391;
	wire signed [31:0] w_sys_tmp6394;
	wire signed [31:0] w_sys_tmp6395;
	wire signed [31:0] w_sys_tmp6396;
	wire signed [31:0] w_sys_tmp6397;
	wire signed [31:0] w_sys_tmp6398;
	wire signed [31:0] w_sys_tmp6399;
	wire signed [31:0] w_sys_tmp6400;
	wire signed [31:0] w_sys_tmp6401;
	wire signed [31:0] w_sys_tmp6402;
	wire signed [31:0] w_sys_tmp6403;
	wire signed [31:0] w_sys_tmp6404;
	wire signed [31:0] w_sys_tmp6405;
	wire signed [31:0] w_sys_tmp6832;
	wire               w_sys_tmp6833;
	wire               w_sys_tmp6834;
	wire signed [31:0] w_sys_tmp6835;
	wire signed [31:0] w_sys_tmp6838;
	wire signed [31:0] w_sys_tmp6839;
	wire signed [31:0] w_sys_tmp6840;
	wire signed [31:0] w_sys_tmp6841;
	wire        [31:0] w_sys_tmp6842;
	wire signed [31:0] w_sys_tmp6843;
	wire signed [31:0] w_sys_tmp6844;
	wire signed [31:0] w_sys_tmp6848;
	wire signed [31:0] w_sys_tmp6849;
	wire signed [31:0] w_sys_tmp6851;
	wire        [31:0] w_sys_tmp6852;
	wire signed [31:0] w_sys_tmp6853;
	wire signed [31:0] w_sys_tmp6854;
	wire signed [31:0] w_sys_tmp6858;
	wire signed [31:0] w_sys_tmp6859;
	wire signed [31:0] w_sys_tmp6861;
	wire signed [31:0] w_sys_tmp6862;
	wire signed [31:0] w_sys_tmp6863;
	wire signed [31:0] w_sys_tmp6867;
	wire signed [31:0] w_sys_tmp6868;
	wire signed [31:0] w_sys_tmp6870;
	wire signed [31:0] w_sys_tmp6872;
	wire signed [31:0] w_sys_tmp6873;
	wire signed [31:0] w_sys_tmp6877;
	wire signed [31:0] w_sys_tmp6878;
	wire signed [31:0] w_sys_tmp6880;
	wire signed [31:0] w_sys_tmp6881;
	wire signed [31:0] w_sys_tmp6882;
	wire signed [31:0] w_sys_tmp6886;
	wire signed [31:0] w_sys_tmp6887;
	wire signed [31:0] w_sys_tmp6889;
	wire        [31:0] w_sys_tmp6890;
	wire signed [31:0] w_sys_tmp6891;
	wire signed [31:0] w_sys_tmp6892;
	wire signed [31:0] w_sys_tmp6895;
	wire signed [31:0] w_sys_tmp6896;
	wire signed [31:0] w_sys_tmp6897;
	wire signed [31:0] w_sys_tmp6898;
	wire signed [31:0] w_sys_tmp6899;
	wire signed [31:0] w_sys_tmp6900;
	wire signed [31:0] w_sys_tmp6901;
	wire signed [31:0] w_sys_tmp6902;
	wire signed [31:0] w_sys_tmp6903;
	wire signed [31:0] w_sys_tmp6904;
	wire signed [31:0] w_sys_tmp6905;
	wire signed [31:0] w_sys_tmp6906;
	wire signed [31:0] w_sys_tmp7333;
	wire               w_sys_tmp7334;
	wire               w_sys_tmp7335;
	wire signed [31:0] w_sys_tmp7336;
	wire signed [31:0] w_sys_tmp7339;
	wire signed [31:0] w_sys_tmp7340;
	wire signed [31:0] w_sys_tmp7341;
	wire signed [31:0] w_sys_tmp7342;
	wire        [31:0] w_sys_tmp7343;
	wire signed [31:0] w_sys_tmp7344;
	wire signed [31:0] w_sys_tmp7345;
	wire signed [31:0] w_sys_tmp7349;
	wire signed [31:0] w_sys_tmp7350;
	wire signed [31:0] w_sys_tmp7352;
	wire        [31:0] w_sys_tmp7353;
	wire signed [31:0] w_sys_tmp7354;
	wire signed [31:0] w_sys_tmp7355;
	wire signed [31:0] w_sys_tmp7359;
	wire signed [31:0] w_sys_tmp7360;
	wire signed [31:0] w_sys_tmp7362;
	wire signed [31:0] w_sys_tmp7363;
	wire signed [31:0] w_sys_tmp7364;
	wire signed [31:0] w_sys_tmp7368;
	wire signed [31:0] w_sys_tmp7369;
	wire signed [31:0] w_sys_tmp7371;
	wire signed [31:0] w_sys_tmp7373;
	wire signed [31:0] w_sys_tmp7374;
	wire signed [31:0] w_sys_tmp7378;
	wire signed [31:0] w_sys_tmp7379;
	wire signed [31:0] w_sys_tmp7381;
	wire signed [31:0] w_sys_tmp7382;
	wire signed [31:0] w_sys_tmp7383;
	wire signed [31:0] w_sys_tmp7387;
	wire signed [31:0] w_sys_tmp7388;
	wire signed [31:0] w_sys_tmp7390;
	wire        [31:0] w_sys_tmp7391;
	wire signed [31:0] w_sys_tmp7392;
	wire signed [31:0] w_sys_tmp7393;
	wire signed [31:0] w_sys_tmp7396;
	wire signed [31:0] w_sys_tmp7397;
	wire signed [31:0] w_sys_tmp7398;
	wire signed [31:0] w_sys_tmp7399;
	wire signed [31:0] w_sys_tmp7400;
	wire signed [31:0] w_sys_tmp7401;
	wire signed [31:0] w_sys_tmp7402;
	wire signed [31:0] w_sys_tmp7403;
	wire signed [31:0] w_sys_tmp7404;
	wire signed [31:0] w_sys_tmp7405;
	wire signed [31:0] w_sys_tmp7406;
	wire signed [31:0] w_sys_tmp7407;
	wire signed [31:0] w_sys_tmp7834;
	wire               w_sys_tmp7835;
	wire               w_sys_tmp7836;
	wire signed [31:0] w_sys_tmp7837;
	wire signed [31:0] w_sys_tmp7840;
	wire signed [31:0] w_sys_tmp7841;
	wire signed [31:0] w_sys_tmp7842;
	wire signed [31:0] w_sys_tmp7843;
	wire        [31:0] w_sys_tmp7844;
	wire signed [31:0] w_sys_tmp7845;
	wire signed [31:0] w_sys_tmp7846;
	wire signed [31:0] w_sys_tmp7850;
	wire signed [31:0] w_sys_tmp7851;
	wire signed [31:0] w_sys_tmp7853;
	wire        [31:0] w_sys_tmp7854;
	wire signed [31:0] w_sys_tmp7855;
	wire signed [31:0] w_sys_tmp7856;
	wire signed [31:0] w_sys_tmp7860;
	wire signed [31:0] w_sys_tmp7861;
	wire signed [31:0] w_sys_tmp7863;
	wire signed [31:0] w_sys_tmp7864;
	wire signed [31:0] w_sys_tmp7865;
	wire signed [31:0] w_sys_tmp7869;
	wire signed [31:0] w_sys_tmp7870;
	wire signed [31:0] w_sys_tmp7872;
	wire signed [31:0] w_sys_tmp7874;
	wire signed [31:0] w_sys_tmp7875;
	wire signed [31:0] w_sys_tmp7879;
	wire signed [31:0] w_sys_tmp7880;
	wire signed [31:0] w_sys_tmp7882;
	wire signed [31:0] w_sys_tmp7883;
	wire signed [31:0] w_sys_tmp7884;
	wire signed [31:0] w_sys_tmp7888;
	wire signed [31:0] w_sys_tmp7889;
	wire signed [31:0] w_sys_tmp7891;
	wire        [31:0] w_sys_tmp7892;
	wire signed [31:0] w_sys_tmp7893;
	wire signed [31:0] w_sys_tmp7894;
	wire signed [31:0] w_sys_tmp7897;
	wire signed [31:0] w_sys_tmp7898;
	wire signed [31:0] w_sys_tmp7899;
	wire signed [31:0] w_sys_tmp7900;
	wire signed [31:0] w_sys_tmp7901;
	wire signed [31:0] w_sys_tmp7902;
	wire signed [31:0] w_sys_tmp7903;
	wire signed [31:0] w_sys_tmp7904;
	wire signed [31:0] w_sys_tmp7905;
	wire signed [31:0] w_sys_tmp7906;
	wire signed [31:0] w_sys_tmp7907;
	wire signed [31:0] w_sys_tmp7908;
	wire signed [31:0] w_sys_tmp8335;
	wire               w_sys_tmp8336;
	wire               w_sys_tmp8337;
	wire signed [31:0] w_sys_tmp8338;
	wire signed [31:0] w_sys_tmp8341;
	wire signed [31:0] w_sys_tmp8342;
	wire signed [31:0] w_sys_tmp8343;
	wire signed [31:0] w_sys_tmp8344;
	wire        [31:0] w_sys_tmp8345;
	wire signed [31:0] w_sys_tmp8346;
	wire signed [31:0] w_sys_tmp8347;
	wire signed [31:0] w_sys_tmp8351;
	wire signed [31:0] w_sys_tmp8352;
	wire signed [31:0] w_sys_tmp8354;
	wire        [31:0] w_sys_tmp8355;
	wire signed [31:0] w_sys_tmp8356;
	wire signed [31:0] w_sys_tmp8357;
	wire signed [31:0] w_sys_tmp8361;
	wire signed [31:0] w_sys_tmp8362;
	wire signed [31:0] w_sys_tmp8364;
	wire signed [31:0] w_sys_tmp8365;
	wire signed [31:0] w_sys_tmp8366;
	wire signed [31:0] w_sys_tmp8370;
	wire signed [31:0] w_sys_tmp8371;
	wire signed [31:0] w_sys_tmp8373;
	wire signed [31:0] w_sys_tmp8375;
	wire signed [31:0] w_sys_tmp8376;
	wire signed [31:0] w_sys_tmp8380;
	wire signed [31:0] w_sys_tmp8381;
	wire signed [31:0] w_sys_tmp8383;
	wire signed [31:0] w_sys_tmp8384;
	wire signed [31:0] w_sys_tmp8385;
	wire signed [31:0] w_sys_tmp8389;
	wire signed [31:0] w_sys_tmp8390;
	wire signed [31:0] w_sys_tmp8392;
	wire        [31:0] w_sys_tmp8393;
	wire signed [31:0] w_sys_tmp8394;
	wire signed [31:0] w_sys_tmp8395;
	wire signed [31:0] w_sys_tmp8398;
	wire signed [31:0] w_sys_tmp8399;
	wire signed [31:0] w_sys_tmp8400;
	wire signed [31:0] w_sys_tmp8401;
	wire signed [31:0] w_sys_tmp8402;
	wire signed [31:0] w_sys_tmp8403;
	wire signed [31:0] w_sys_tmp8404;
	wire signed [31:0] w_sys_tmp8405;
	wire signed [31:0] w_sys_tmp8406;
	wire signed [31:0] w_sys_tmp8407;
	wire signed [31:0] w_sys_tmp8408;
	wire signed [31:0] w_sys_tmp8409;
	wire signed [31:0] w_sys_tmp8836;
	wire               w_sys_tmp8837;
	wire               w_sys_tmp8838;
	wire signed [31:0] w_sys_tmp8839;
	wire signed [31:0] w_sys_tmp8842;
	wire signed [31:0] w_sys_tmp8843;
	wire signed [31:0] w_sys_tmp8844;
	wire signed [31:0] w_sys_tmp8845;
	wire        [31:0] w_sys_tmp8846;
	wire signed [31:0] w_sys_tmp8847;
	wire signed [31:0] w_sys_tmp8848;
	wire signed [31:0] w_sys_tmp8852;
	wire signed [31:0] w_sys_tmp8853;
	wire signed [31:0] w_sys_tmp8855;
	wire        [31:0] w_sys_tmp8856;
	wire signed [31:0] w_sys_tmp8857;
	wire signed [31:0] w_sys_tmp8858;
	wire signed [31:0] w_sys_tmp8862;
	wire signed [31:0] w_sys_tmp8863;
	wire signed [31:0] w_sys_tmp8865;
	wire signed [31:0] w_sys_tmp8866;
	wire signed [31:0] w_sys_tmp8867;
	wire signed [31:0] w_sys_tmp8871;
	wire signed [31:0] w_sys_tmp8872;
	wire signed [31:0] w_sys_tmp8874;
	wire signed [31:0] w_sys_tmp8876;
	wire signed [31:0] w_sys_tmp8877;
	wire signed [31:0] w_sys_tmp8881;
	wire signed [31:0] w_sys_tmp8882;
	wire signed [31:0] w_sys_tmp8884;
	wire signed [31:0] w_sys_tmp8885;
	wire signed [31:0] w_sys_tmp8886;
	wire signed [31:0] w_sys_tmp8890;
	wire signed [31:0] w_sys_tmp8891;
	wire signed [31:0] w_sys_tmp8893;
	wire        [31:0] w_sys_tmp8894;
	wire signed [31:0] w_sys_tmp8895;
	wire signed [31:0] w_sys_tmp8896;
	wire signed [31:0] w_sys_tmp8899;
	wire signed [31:0] w_sys_tmp8900;
	wire signed [31:0] w_sys_tmp8901;
	wire signed [31:0] w_sys_tmp8902;
	wire signed [31:0] w_sys_tmp8903;
	wire signed [31:0] w_sys_tmp8904;
	wire signed [31:0] w_sys_tmp8905;
	wire signed [31:0] w_sys_tmp8906;
	wire signed [31:0] w_sys_tmp8907;
	wire signed [31:0] w_sys_tmp8908;
	wire signed [31:0] w_sys_tmp8909;
	wire signed [31:0] w_sys_tmp8910;
	wire signed [31:0] w_sys_tmp9325;
	wire               w_sys_tmp9326;
	wire               w_sys_tmp9327;
	wire signed [31:0] w_sys_tmp9328;
	wire signed [31:0] w_sys_tmp9329;
	wire signed [31:0] w_sys_tmp9330;
	wire               w_sys_tmp9331;
	wire               w_sys_tmp9332;
	wire signed [31:0] w_sys_tmp9333;
	wire signed [31:0] w_sys_tmp9336;
	wire signed [31:0] w_sys_tmp9337;
	wire signed [31:0] w_sys_tmp9338;
	wire        [31:0] w_sys_tmp9339;
	wire signed [31:0] w_sys_tmp9340;
	wire signed [31:0] w_sys_tmp9341;
	wire signed [31:0] w_sys_tmp9343;
	wire signed [31:0] w_sys_tmp9344;
	wire signed [31:0] w_sys_tmp9405;
	wire               w_sys_tmp9406;
	wire               w_sys_tmp9407;
	wire signed [31:0] w_sys_tmp9408;
	wire signed [31:0] w_sys_tmp9410;
	wire signed [31:0] w_sys_tmp9411;
	wire signed [31:0] w_sys_tmp9413;
	wire signed [31:0] w_sys_tmp9414;
	wire signed [31:0] w_sys_tmp9415;
	wire        [31:0] w_sys_tmp9416;
	wire signed [31:0] w_sys_tmp9417;
	wire signed [31:0] w_sys_tmp9418;
	wire signed [31:0] w_sys_tmp9420;
	wire signed [31:0] w_sys_tmp9421;
	wire signed [31:0] w_sys_tmp9422;
	wire signed [31:0] w_sys_tmp9501;
	wire               w_sys_tmp9502;
	wire               w_sys_tmp9503;
	wire signed [31:0] w_sys_tmp9504;
	wire signed [31:0] w_sys_tmp9506;
	wire signed [31:0] w_sys_tmp9507;
	wire signed [31:0] w_sys_tmp9509;
	wire signed [31:0] w_sys_tmp9510;
	wire signed [31:0] w_sys_tmp9511;
	wire        [31:0] w_sys_tmp9512;
	wire signed [31:0] w_sys_tmp9513;
	wire signed [31:0] w_sys_tmp9514;
	wire signed [31:0] w_sys_tmp9516;
	wire signed [31:0] w_sys_tmp9517;
	wire signed [31:0] w_sys_tmp9518;
	wire signed [31:0] w_sys_tmp9597;
	wire               w_sys_tmp9598;
	wire               w_sys_tmp9599;
	wire signed [31:0] w_sys_tmp9600;
	wire signed [31:0] w_sys_tmp9602;
	wire signed [31:0] w_sys_tmp9603;
	wire signed [31:0] w_sys_tmp9605;
	wire signed [31:0] w_sys_tmp9606;
	wire signed [31:0] w_sys_tmp9607;
	wire        [31:0] w_sys_tmp9608;
	wire signed [31:0] w_sys_tmp9609;
	wire signed [31:0] w_sys_tmp9610;
	wire signed [31:0] w_sys_tmp9612;
	wire signed [31:0] w_sys_tmp9613;
	wire signed [31:0] w_sys_tmp9614;
	wire signed [31:0] w_sys_tmp9693;
	wire               w_sys_tmp9694;
	wire               w_sys_tmp9695;
	wire signed [31:0] w_sys_tmp9696;
	wire signed [31:0] w_sys_tmp9698;
	wire signed [31:0] w_sys_tmp9699;
	wire signed [31:0] w_sys_tmp9701;
	wire signed [31:0] w_sys_tmp9702;
	wire signed [31:0] w_sys_tmp9703;
	wire        [31:0] w_sys_tmp9704;
	wire signed [31:0] w_sys_tmp9705;
	wire signed [31:0] w_sys_tmp9706;
	wire signed [31:0] w_sys_tmp9708;
	wire signed [31:0] w_sys_tmp9709;
	wire signed [31:0] w_sys_tmp9710;
	wire signed [31:0] w_sys_tmp9789;
	wire               w_sys_tmp9790;
	wire               w_sys_tmp9791;
	wire signed [31:0] w_sys_tmp9792;
	wire signed [31:0] w_sys_tmp9794;
	wire signed [31:0] w_sys_tmp9795;
	wire signed [31:0] w_sys_tmp9797;
	wire signed [31:0] w_sys_tmp9798;
	wire signed [31:0] w_sys_tmp9799;
	wire        [31:0] w_sys_tmp9800;
	wire signed [31:0] w_sys_tmp9801;
	wire signed [31:0] w_sys_tmp9802;
	wire signed [31:0] w_sys_tmp9804;
	wire signed [31:0] w_sys_tmp9805;
	wire signed [31:0] w_sys_tmp9806;
	wire signed [31:0] w_sys_tmp9885;
	wire               w_sys_tmp9886;
	wire               w_sys_tmp9887;
	wire signed [31:0] w_sys_tmp9888;
	wire signed [31:0] w_sys_tmp9890;
	wire signed [31:0] w_sys_tmp9891;
	wire signed [31:0] w_sys_tmp9893;
	wire signed [31:0] w_sys_tmp9894;
	wire signed [31:0] w_sys_tmp9895;
	wire        [31:0] w_sys_tmp9896;
	wire signed [31:0] w_sys_tmp9897;
	wire signed [31:0] w_sys_tmp9898;
	wire signed [31:0] w_sys_tmp9900;
	wire signed [31:0] w_sys_tmp9901;
	wire signed [31:0] w_sys_tmp9902;
	wire signed [31:0] w_sys_tmp9981;
	wire               w_sys_tmp9982;
	wire               w_sys_tmp9983;
	wire signed [31:0] w_sys_tmp9984;
	wire signed [31:0] w_sys_tmp9986;
	wire signed [31:0] w_sys_tmp9987;
	wire signed [31:0] w_sys_tmp9989;
	wire signed [31:0] w_sys_tmp9990;
	wire signed [31:0] w_sys_tmp9991;
	wire        [31:0] w_sys_tmp9992;
	wire signed [31:0] w_sys_tmp9993;
	wire signed [31:0] w_sys_tmp9994;
	wire signed [31:0] w_sys_tmp9996;
	wire signed [31:0] w_sys_tmp9997;
	wire signed [31:0] w_sys_tmp9998;
	wire signed [31:0] w_sys_tmp10077;
	wire               w_sys_tmp10078;
	wire               w_sys_tmp10079;
	wire signed [31:0] w_sys_tmp10080;
	wire signed [31:0] w_sys_tmp10081;
	wire signed [31:0] w_sys_tmp10082;
	wire               w_sys_tmp10083;
	wire               w_sys_tmp10084;
	wire signed [31:0] w_sys_tmp10085;
	wire signed [31:0] w_sys_tmp10088;
	wire signed [31:0] w_sys_tmp10089;
	wire signed [31:0] w_sys_tmp10090;
	wire        [31:0] w_sys_tmp10091;
	wire signed [31:0] w_sys_tmp10092;
	wire signed [31:0] w_sys_tmp10093;
	wire signed [31:0] w_sys_tmp10095;
	wire signed [31:0] w_sys_tmp10096;
	wire signed [31:0] w_sys_tmp10157;
	wire               w_sys_tmp10158;
	wire               w_sys_tmp10159;
	wire signed [31:0] w_sys_tmp10160;
	wire signed [31:0] w_sys_tmp10162;
	wire signed [31:0] w_sys_tmp10163;
	wire signed [31:0] w_sys_tmp10165;
	wire signed [31:0] w_sys_tmp10166;
	wire signed [31:0] w_sys_tmp10167;
	wire        [31:0] w_sys_tmp10168;
	wire signed [31:0] w_sys_tmp10169;
	wire signed [31:0] w_sys_tmp10170;
	wire signed [31:0] w_sys_tmp10172;
	wire signed [31:0] w_sys_tmp10173;
	wire signed [31:0] w_sys_tmp10174;
	wire signed [31:0] w_sys_tmp10253;
	wire               w_sys_tmp10254;
	wire               w_sys_tmp10255;
	wire signed [31:0] w_sys_tmp10256;
	wire signed [31:0] w_sys_tmp10258;
	wire signed [31:0] w_sys_tmp10259;
	wire signed [31:0] w_sys_tmp10261;
	wire signed [31:0] w_sys_tmp10262;
	wire signed [31:0] w_sys_tmp10263;
	wire        [31:0] w_sys_tmp10264;
	wire signed [31:0] w_sys_tmp10265;
	wire signed [31:0] w_sys_tmp10266;
	wire signed [31:0] w_sys_tmp10268;
	wire signed [31:0] w_sys_tmp10269;
	wire signed [31:0] w_sys_tmp10270;
	wire signed [31:0] w_sys_tmp10349;
	wire               w_sys_tmp10350;
	wire               w_sys_tmp10351;
	wire signed [31:0] w_sys_tmp10352;
	wire signed [31:0] w_sys_tmp10354;
	wire signed [31:0] w_sys_tmp10355;
	wire signed [31:0] w_sys_tmp10357;
	wire signed [31:0] w_sys_tmp10358;
	wire signed [31:0] w_sys_tmp10359;
	wire        [31:0] w_sys_tmp10360;
	wire signed [31:0] w_sys_tmp10361;
	wire signed [31:0] w_sys_tmp10362;
	wire signed [31:0] w_sys_tmp10364;
	wire signed [31:0] w_sys_tmp10365;
	wire signed [31:0] w_sys_tmp10366;
	wire signed [31:0] w_sys_tmp10445;
	wire               w_sys_tmp10446;
	wire               w_sys_tmp10447;
	wire signed [31:0] w_sys_tmp10448;
	wire signed [31:0] w_sys_tmp10450;
	wire signed [31:0] w_sys_tmp10451;
	wire signed [31:0] w_sys_tmp10453;
	wire signed [31:0] w_sys_tmp10454;
	wire signed [31:0] w_sys_tmp10455;
	wire        [31:0] w_sys_tmp10456;
	wire signed [31:0] w_sys_tmp10457;
	wire signed [31:0] w_sys_tmp10458;
	wire signed [31:0] w_sys_tmp10460;
	wire signed [31:0] w_sys_tmp10461;
	wire signed [31:0] w_sys_tmp10462;
	wire signed [31:0] w_sys_tmp10541;
	wire               w_sys_tmp10542;
	wire               w_sys_tmp10543;
	wire signed [31:0] w_sys_tmp10544;
	wire signed [31:0] w_sys_tmp10546;
	wire signed [31:0] w_sys_tmp10547;
	wire signed [31:0] w_sys_tmp10549;
	wire signed [31:0] w_sys_tmp10550;
	wire signed [31:0] w_sys_tmp10551;
	wire        [31:0] w_sys_tmp10552;
	wire signed [31:0] w_sys_tmp10553;
	wire signed [31:0] w_sys_tmp10554;
	wire signed [31:0] w_sys_tmp10556;
	wire signed [31:0] w_sys_tmp10557;
	wire signed [31:0] w_sys_tmp10558;
	wire signed [31:0] w_sys_tmp10637;
	wire               w_sys_tmp10638;
	wire               w_sys_tmp10639;
	wire signed [31:0] w_sys_tmp10640;
	wire signed [31:0] w_sys_tmp10642;
	wire signed [31:0] w_sys_tmp10643;
	wire signed [31:0] w_sys_tmp10645;
	wire signed [31:0] w_sys_tmp10646;
	wire signed [31:0] w_sys_tmp10647;
	wire        [31:0] w_sys_tmp10648;
	wire signed [31:0] w_sys_tmp10649;
	wire signed [31:0] w_sys_tmp10650;
	wire signed [31:0] w_sys_tmp10652;
	wire signed [31:0] w_sys_tmp10653;
	wire signed [31:0] w_sys_tmp10654;
	wire signed [31:0] w_sys_tmp10733;
	wire               w_sys_tmp10734;
	wire               w_sys_tmp10735;
	wire signed [31:0] w_sys_tmp10736;
	wire signed [31:0] w_sys_tmp10738;
	wire signed [31:0] w_sys_tmp10739;
	wire signed [31:0] w_sys_tmp10741;
	wire signed [31:0] w_sys_tmp10742;
	wire signed [31:0] w_sys_tmp10743;
	wire        [31:0] w_sys_tmp10744;
	wire signed [31:0] w_sys_tmp10745;
	wire signed [31:0] w_sys_tmp10746;
	wire signed [31:0] w_sys_tmp10748;
	wire signed [31:0] w_sys_tmp10749;
	wire signed [31:0] w_sys_tmp10750;
	wire signed [31:0] w_sys_tmp10829;
	wire               w_sys_tmp10830;
	wire               w_sys_tmp10831;
	wire signed [31:0] w_sys_tmp10832;
	wire signed [31:0] w_sys_tmp10833;
	wire signed [31:0] w_sys_tmp10834;
	wire               w_sys_tmp10835;
	wire               w_sys_tmp10836;
	wire signed [31:0] w_sys_tmp10837;
	wire signed [31:0] w_sys_tmp10840;
	wire signed [31:0] w_sys_tmp10841;
	wire signed [31:0] w_sys_tmp10842;
	wire        [31:0] w_sys_tmp10843;
	wire signed [31:0] w_sys_tmp10844;
	wire signed [31:0] w_sys_tmp10845;
	wire signed [31:0] w_sys_tmp10847;
	wire signed [31:0] w_sys_tmp10848;
	wire signed [31:0] w_sys_tmp10909;
	wire               w_sys_tmp10910;
	wire               w_sys_tmp10911;
	wire signed [31:0] w_sys_tmp10912;
	wire signed [31:0] w_sys_tmp10914;
	wire signed [31:0] w_sys_tmp10915;
	wire signed [31:0] w_sys_tmp10917;
	wire signed [31:0] w_sys_tmp10918;
	wire signed [31:0] w_sys_tmp10919;
	wire        [31:0] w_sys_tmp10920;
	wire signed [31:0] w_sys_tmp10921;
	wire signed [31:0] w_sys_tmp10922;
	wire signed [31:0] w_sys_tmp10924;
	wire signed [31:0] w_sys_tmp10925;
	wire signed [31:0] w_sys_tmp10926;
	wire signed [31:0] w_sys_tmp11005;
	wire               w_sys_tmp11006;
	wire               w_sys_tmp11007;
	wire signed [31:0] w_sys_tmp11008;
	wire signed [31:0] w_sys_tmp11010;
	wire signed [31:0] w_sys_tmp11011;
	wire signed [31:0] w_sys_tmp11013;
	wire signed [31:0] w_sys_tmp11014;
	wire signed [31:0] w_sys_tmp11015;
	wire        [31:0] w_sys_tmp11016;
	wire signed [31:0] w_sys_tmp11017;
	wire signed [31:0] w_sys_tmp11018;
	wire signed [31:0] w_sys_tmp11020;
	wire signed [31:0] w_sys_tmp11021;
	wire signed [31:0] w_sys_tmp11022;
	wire signed [31:0] w_sys_tmp11101;
	wire               w_sys_tmp11102;
	wire               w_sys_tmp11103;
	wire signed [31:0] w_sys_tmp11104;
	wire signed [31:0] w_sys_tmp11106;
	wire signed [31:0] w_sys_tmp11107;
	wire signed [31:0] w_sys_tmp11109;
	wire signed [31:0] w_sys_tmp11110;
	wire signed [31:0] w_sys_tmp11111;
	wire        [31:0] w_sys_tmp11112;
	wire signed [31:0] w_sys_tmp11113;
	wire signed [31:0] w_sys_tmp11114;
	wire signed [31:0] w_sys_tmp11116;
	wire signed [31:0] w_sys_tmp11117;
	wire signed [31:0] w_sys_tmp11118;
	wire signed [31:0] w_sys_tmp11197;
	wire               w_sys_tmp11198;
	wire               w_sys_tmp11199;
	wire signed [31:0] w_sys_tmp11200;
	wire signed [31:0] w_sys_tmp11202;
	wire signed [31:0] w_sys_tmp11203;
	wire signed [31:0] w_sys_tmp11205;
	wire signed [31:0] w_sys_tmp11206;
	wire signed [31:0] w_sys_tmp11207;
	wire        [31:0] w_sys_tmp11208;
	wire signed [31:0] w_sys_tmp11209;
	wire signed [31:0] w_sys_tmp11210;
	wire signed [31:0] w_sys_tmp11212;
	wire signed [31:0] w_sys_tmp11213;
	wire signed [31:0] w_sys_tmp11214;
	wire signed [31:0] w_sys_tmp11293;
	wire               w_sys_tmp11294;
	wire               w_sys_tmp11295;
	wire signed [31:0] w_sys_tmp11296;
	wire signed [31:0] w_sys_tmp11298;
	wire signed [31:0] w_sys_tmp11299;
	wire signed [31:0] w_sys_tmp11301;
	wire signed [31:0] w_sys_tmp11302;
	wire signed [31:0] w_sys_tmp11303;
	wire        [31:0] w_sys_tmp11304;
	wire signed [31:0] w_sys_tmp11305;
	wire signed [31:0] w_sys_tmp11306;
	wire signed [31:0] w_sys_tmp11308;
	wire signed [31:0] w_sys_tmp11309;
	wire signed [31:0] w_sys_tmp11310;
	wire signed [31:0] w_sys_tmp11389;
	wire               w_sys_tmp11390;
	wire               w_sys_tmp11391;
	wire signed [31:0] w_sys_tmp11392;
	wire signed [31:0] w_sys_tmp11394;
	wire signed [31:0] w_sys_tmp11395;
	wire signed [31:0] w_sys_tmp11397;
	wire signed [31:0] w_sys_tmp11398;
	wire signed [31:0] w_sys_tmp11399;
	wire        [31:0] w_sys_tmp11400;
	wire signed [31:0] w_sys_tmp11401;
	wire signed [31:0] w_sys_tmp11402;
	wire signed [31:0] w_sys_tmp11404;
	wire signed [31:0] w_sys_tmp11405;
	wire signed [31:0] w_sys_tmp11406;
	wire signed [31:0] w_sys_tmp11485;
	wire               w_sys_tmp11486;
	wire               w_sys_tmp11487;
	wire signed [31:0] w_sys_tmp11488;
	wire signed [31:0] w_sys_tmp11490;
	wire signed [31:0] w_sys_tmp11491;
	wire signed [31:0] w_sys_tmp11493;
	wire signed [31:0] w_sys_tmp11494;
	wire signed [31:0] w_sys_tmp11495;
	wire        [31:0] w_sys_tmp11496;
	wire signed [31:0] w_sys_tmp11497;
	wire signed [31:0] w_sys_tmp11498;
	wire signed [31:0] w_sys_tmp11500;
	wire signed [31:0] w_sys_tmp11501;
	wire signed [31:0] w_sys_tmp11502;
	wire signed [31:0] w_sys_tmp11581;
	wire               w_sys_tmp11582;
	wire               w_sys_tmp11583;
	wire signed [31:0] w_sys_tmp11584;
	wire signed [31:0] w_sys_tmp11585;
	wire signed [31:0] w_sys_tmp11586;
	wire               w_sys_tmp11587;
	wire               w_sys_tmp11588;
	wire signed [31:0] w_sys_tmp11589;
	wire signed [31:0] w_sys_tmp11592;
	wire signed [31:0] w_sys_tmp11593;
	wire signed [31:0] w_sys_tmp11594;
	wire        [31:0] w_sys_tmp11595;
	wire signed [31:0] w_sys_tmp11596;
	wire signed [31:0] w_sys_tmp11597;
	wire signed [31:0] w_sys_tmp11599;
	wire signed [31:0] w_sys_tmp11600;
	wire signed [31:0] w_sys_tmp11661;
	wire               w_sys_tmp11662;
	wire               w_sys_tmp11663;
	wire signed [31:0] w_sys_tmp11664;
	wire signed [31:0] w_sys_tmp11666;
	wire signed [31:0] w_sys_tmp11667;
	wire signed [31:0] w_sys_tmp11669;
	wire signed [31:0] w_sys_tmp11670;
	wire signed [31:0] w_sys_tmp11671;
	wire        [31:0] w_sys_tmp11672;
	wire signed [31:0] w_sys_tmp11673;
	wire signed [31:0] w_sys_tmp11674;
	wire signed [31:0] w_sys_tmp11676;
	wire signed [31:0] w_sys_tmp11677;
	wire signed [31:0] w_sys_tmp11678;
	wire signed [31:0] w_sys_tmp11757;
	wire               w_sys_tmp11758;
	wire               w_sys_tmp11759;
	wire signed [31:0] w_sys_tmp11760;
	wire signed [31:0] w_sys_tmp11762;
	wire signed [31:0] w_sys_tmp11763;
	wire signed [31:0] w_sys_tmp11765;
	wire signed [31:0] w_sys_tmp11766;
	wire signed [31:0] w_sys_tmp11767;
	wire        [31:0] w_sys_tmp11768;
	wire signed [31:0] w_sys_tmp11769;
	wire signed [31:0] w_sys_tmp11770;
	wire signed [31:0] w_sys_tmp11772;
	wire signed [31:0] w_sys_tmp11773;
	wire signed [31:0] w_sys_tmp11774;
	wire signed [31:0] w_sys_tmp11853;
	wire               w_sys_tmp11854;
	wire               w_sys_tmp11855;
	wire signed [31:0] w_sys_tmp11856;
	wire signed [31:0] w_sys_tmp11858;
	wire signed [31:0] w_sys_tmp11859;
	wire signed [31:0] w_sys_tmp11861;
	wire signed [31:0] w_sys_tmp11862;
	wire signed [31:0] w_sys_tmp11863;
	wire        [31:0] w_sys_tmp11864;
	wire signed [31:0] w_sys_tmp11865;
	wire signed [31:0] w_sys_tmp11866;
	wire signed [31:0] w_sys_tmp11868;
	wire signed [31:0] w_sys_tmp11869;
	wire signed [31:0] w_sys_tmp11870;
	wire signed [31:0] w_sys_tmp11949;
	wire               w_sys_tmp11950;
	wire               w_sys_tmp11951;
	wire signed [31:0] w_sys_tmp11952;
	wire signed [31:0] w_sys_tmp11954;
	wire signed [31:0] w_sys_tmp11955;
	wire signed [31:0] w_sys_tmp11957;
	wire signed [31:0] w_sys_tmp11958;
	wire signed [31:0] w_sys_tmp11959;
	wire        [31:0] w_sys_tmp11960;
	wire signed [31:0] w_sys_tmp11961;
	wire signed [31:0] w_sys_tmp11962;
	wire signed [31:0] w_sys_tmp11964;
	wire signed [31:0] w_sys_tmp11965;
	wire signed [31:0] w_sys_tmp11966;
	wire signed [31:0] w_sys_tmp12045;
	wire               w_sys_tmp12046;
	wire               w_sys_tmp12047;
	wire signed [31:0] w_sys_tmp12048;
	wire signed [31:0] w_sys_tmp12050;
	wire signed [31:0] w_sys_tmp12051;
	wire signed [31:0] w_sys_tmp12053;
	wire signed [31:0] w_sys_tmp12054;
	wire signed [31:0] w_sys_tmp12055;
	wire        [31:0] w_sys_tmp12056;
	wire signed [31:0] w_sys_tmp12057;
	wire signed [31:0] w_sys_tmp12058;
	wire signed [31:0] w_sys_tmp12060;
	wire signed [31:0] w_sys_tmp12061;
	wire signed [31:0] w_sys_tmp12062;
	wire signed [31:0] w_sys_tmp12141;
	wire               w_sys_tmp12142;
	wire               w_sys_tmp12143;
	wire signed [31:0] w_sys_tmp12144;
	wire signed [31:0] w_sys_tmp12146;
	wire signed [31:0] w_sys_tmp12147;
	wire signed [31:0] w_sys_tmp12149;
	wire signed [31:0] w_sys_tmp12150;
	wire signed [31:0] w_sys_tmp12151;
	wire        [31:0] w_sys_tmp12152;
	wire signed [31:0] w_sys_tmp12153;
	wire signed [31:0] w_sys_tmp12154;
	wire signed [31:0] w_sys_tmp12156;
	wire signed [31:0] w_sys_tmp12157;
	wire signed [31:0] w_sys_tmp12158;
	wire signed [31:0] w_sys_tmp12237;
	wire               w_sys_tmp12238;
	wire               w_sys_tmp12239;
	wire signed [31:0] w_sys_tmp12240;
	wire signed [31:0] w_sys_tmp12242;
	wire signed [31:0] w_sys_tmp12243;
	wire signed [31:0] w_sys_tmp12245;
	wire signed [31:0] w_sys_tmp12246;
	wire signed [31:0] w_sys_tmp12247;
	wire        [31:0] w_sys_tmp12248;
	wire signed [31:0] w_sys_tmp12249;
	wire signed [31:0] w_sys_tmp12250;
	wire signed [31:0] w_sys_tmp12252;
	wire signed [31:0] w_sys_tmp12253;
	wire signed [31:0] w_sys_tmp12254;
	wire        [31:0] w_sys_tmp12333;
	wire signed [31:0] w_sys_tmp12334;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign o_run_return = r_sys_run_return;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 6'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 6'h1);
	assign w_fld_T_0_addr_0 = 15'sh0;
	assign w_fld_T_0_datain_0 = 32'h0;
	assign w_fld_T_0_r_w_0 = 1'h0;
	assign w_fld_T_0_ce_0 = w_sys_ce;
	assign w_fld_T_0_ce_1 = w_sys_ce;
	assign w_fld_TT_1_addr_0 = 15'sh0;
	assign w_fld_TT_1_datain_0 = 32'h0;
	assign w_fld_TT_1_r_w_0 = 1'h0;
	assign w_fld_TT_1_ce_0 = w_sys_ce;
	assign w_fld_TT_1_ce_1 = w_sys_ce;
	assign w_fld_U_2_addr_0 = 15'sh0;
	assign w_fld_U_2_datain_0 = 32'h0;
	assign w_fld_U_2_r_w_0 = 1'h0;
	assign w_fld_U_2_ce_0 = w_sys_ce;
	assign w_fld_U_2_ce_1 = w_sys_ce;
	assign w_sub19_T_addr = ( (|r_sys_processing_methodID) ? r_sub19_T_addr : 12'sh0 ) ;
	assign w_sub19_T_datain = ( (|r_sys_processing_methodID) ? r_sub19_T_datain : 32'h0 ) ;
	assign w_sub19_T_r_w = ( (|r_sys_processing_methodID) ? r_sub19_T_r_w : 1'h0 ) ;
	assign w_sub19_U_addr = ( (|r_sys_processing_methodID) ? r_sub19_U_addr : 12'sh0 ) ;
	assign w_sub19_U_datain = ( (|r_sys_processing_methodID) ? r_sub19_U_datain : 32'h0 ) ;
	assign w_sub19_U_r_w = ( (|r_sys_processing_methodID) ? r_sub19_U_r_w : 1'h0 ) ;
	assign w_sub19_result_addr = ( (|r_sys_processing_methodID) ? r_sub19_result_addr : 12'sh0 ) ;
	assign w_sub19_result_datain = ( (|r_sys_processing_methodID) ? r_sub19_result_datain : 32'h0 ) ;
	assign w_sub19_result_r_w = ( (|r_sys_processing_methodID) ? r_sub19_result_r_w : 1'h0 ) ;
	assign w_sub12_T_addr = ( (|r_sys_processing_methodID) ? r_sub12_T_addr : 12'sh0 ) ;
	assign w_sub12_T_datain = ( (|r_sys_processing_methodID) ? r_sub12_T_datain : 32'h0 ) ;
	assign w_sub12_T_r_w = ( (|r_sys_processing_methodID) ? r_sub12_T_r_w : 1'h0 ) ;
	assign w_sub12_U_addr = ( (|r_sys_processing_methodID) ? r_sub12_U_addr : 12'sh0 ) ;
	assign w_sub12_U_datain = ( (|r_sys_processing_methodID) ? r_sub12_U_datain : 32'h0 ) ;
	assign w_sub12_U_r_w = ( (|r_sys_processing_methodID) ? r_sub12_U_r_w : 1'h0 ) ;
	assign w_sub12_result_addr = ( (|r_sys_processing_methodID) ? r_sub12_result_addr : 12'sh0 ) ;
	assign w_sub12_result_datain = ( (|r_sys_processing_methodID) ? r_sub12_result_datain : 32'h0 ) ;
	assign w_sub12_result_r_w = ( (|r_sys_processing_methodID) ? r_sub12_result_r_w : 1'h0 ) ;
	assign w_sub11_T_addr = ( (|r_sys_processing_methodID) ? r_sub11_T_addr : 12'sh0 ) ;
	assign w_sub11_T_datain = ( (|r_sys_processing_methodID) ? r_sub11_T_datain : 32'h0 ) ;
	assign w_sub11_T_r_w = ( (|r_sys_processing_methodID) ? r_sub11_T_r_w : 1'h0 ) ;
	assign w_sub11_V_addr = ( (|r_sys_processing_methodID) ? r_sub11_V_addr : 12'sh0 ) ;
	assign w_sub11_V_datain = ( (|r_sys_processing_methodID) ? r_sub11_V_datain : 32'h0 ) ;
	assign w_sub11_V_r_w = ( (|r_sys_processing_methodID) ? r_sub11_V_r_w : 1'h0 ) ;
	assign w_sub11_U_addr = ( (|r_sys_processing_methodID) ? r_sub11_U_addr : 12'sh0 ) ;
	assign w_sub11_U_datain = ( (|r_sys_processing_methodID) ? r_sub11_U_datain : 32'h0 ) ;
	assign w_sub11_U_r_w = ( (|r_sys_processing_methodID) ? r_sub11_U_r_w : 1'h0 ) ;
	assign w_sub11_result_addr = ( (|r_sys_processing_methodID) ? r_sub11_result_addr : 12'sh0 ) ;
	assign w_sub11_result_datain = ( (|r_sys_processing_methodID) ? r_sub11_result_datain : 32'h0 ) ;
	assign w_sub11_result_r_w = ( (|r_sys_processing_methodID) ? r_sub11_result_r_w : 1'h0 ) ;
	assign w_sub14_T_addr = ( (|r_sys_processing_methodID) ? r_sub14_T_addr : 12'sh0 ) ;
	assign w_sub14_T_datain = ( (|r_sys_processing_methodID) ? r_sub14_T_datain : 32'h0 ) ;
	assign w_sub14_T_r_w = ( (|r_sys_processing_methodID) ? r_sub14_T_r_w : 1'h0 ) ;
	assign w_sub14_U_addr = ( (|r_sys_processing_methodID) ? r_sub14_U_addr : 12'sh0 ) ;
	assign w_sub14_U_datain = ( (|r_sys_processing_methodID) ? r_sub14_U_datain : 32'h0 ) ;
	assign w_sub14_U_r_w = ( (|r_sys_processing_methodID) ? r_sub14_U_r_w : 1'h0 ) ;
	assign w_sub14_result_addr = ( (|r_sys_processing_methodID) ? r_sub14_result_addr : 12'sh0 ) ;
	assign w_sub14_result_datain = ( (|r_sys_processing_methodID) ? r_sub14_result_datain : 32'h0 ) ;
	assign w_sub14_result_r_w = ( (|r_sys_processing_methodID) ? r_sub14_result_r_w : 1'h0 ) ;
	assign w_sub13_T_addr = ( (|r_sys_processing_methodID) ? r_sub13_T_addr : 12'sh0 ) ;
	assign w_sub13_T_datain = ( (|r_sys_processing_methodID) ? r_sub13_T_datain : 32'h0 ) ;
	assign w_sub13_T_r_w = ( (|r_sys_processing_methodID) ? r_sub13_T_r_w : 1'h0 ) ;
	assign w_sub13_U_addr = ( (|r_sys_processing_methodID) ? r_sub13_U_addr : 12'sh0 ) ;
	assign w_sub13_U_datain = ( (|r_sys_processing_methodID) ? r_sub13_U_datain : 32'h0 ) ;
	assign w_sub13_U_r_w = ( (|r_sys_processing_methodID) ? r_sub13_U_r_w : 1'h0 ) ;
	assign w_sub13_result_addr = ( (|r_sys_processing_methodID) ? r_sub13_result_addr : 12'sh0 ) ;
	assign w_sub13_result_datain = ( (|r_sys_processing_methodID) ? r_sub13_result_datain : 32'h0 ) ;
	assign w_sub13_result_r_w = ( (|r_sys_processing_methodID) ? r_sub13_result_r_w : 1'h0 ) ;
	assign w_sub16_T_addr = ( (|r_sys_processing_methodID) ? r_sub16_T_addr : 12'sh0 ) ;
	assign w_sub16_T_datain = ( (|r_sys_processing_methodID) ? r_sub16_T_datain : 32'h0 ) ;
	assign w_sub16_T_r_w = ( (|r_sys_processing_methodID) ? r_sub16_T_r_w : 1'h0 ) ;
	assign w_sub16_U_addr = ( (|r_sys_processing_methodID) ? r_sub16_U_addr : 12'sh0 ) ;
	assign w_sub16_U_datain = ( (|r_sys_processing_methodID) ? r_sub16_U_datain : 32'h0 ) ;
	assign w_sub16_U_r_w = ( (|r_sys_processing_methodID) ? r_sub16_U_r_w : 1'h0 ) ;
	assign w_sub16_result_addr = ( (|r_sys_processing_methodID) ? r_sub16_result_addr : 12'sh0 ) ;
	assign w_sub16_result_datain = ( (|r_sys_processing_methodID) ? r_sub16_result_datain : 32'h0 ) ;
	assign w_sub16_result_r_w = ( (|r_sys_processing_methodID) ? r_sub16_result_r_w : 1'h0 ) ;
	assign w_sub15_T_addr = ( (|r_sys_processing_methodID) ? r_sub15_T_addr : 12'sh0 ) ;
	assign w_sub15_T_datain = ( (|r_sys_processing_methodID) ? r_sub15_T_datain : 32'h0 ) ;
	assign w_sub15_T_r_w = ( (|r_sys_processing_methodID) ? r_sub15_T_r_w : 1'h0 ) ;
	assign w_sub15_U_addr = ( (|r_sys_processing_methodID) ? r_sub15_U_addr : 12'sh0 ) ;
	assign w_sub15_U_datain = ( (|r_sys_processing_methodID) ? r_sub15_U_datain : 32'h0 ) ;
	assign w_sub15_U_r_w = ( (|r_sys_processing_methodID) ? r_sub15_U_r_w : 1'h0 ) ;
	assign w_sub15_result_addr = ( (|r_sys_processing_methodID) ? r_sub15_result_addr : 12'sh0 ) ;
	assign w_sub15_result_datain = ( (|r_sys_processing_methodID) ? r_sub15_result_datain : 32'h0 ) ;
	assign w_sub15_result_r_w = ( (|r_sys_processing_methodID) ? r_sub15_result_r_w : 1'h0 ) ;
	assign w_sub18_T_addr = ( (|r_sys_processing_methodID) ? r_sub18_T_addr : 12'sh0 ) ;
	assign w_sub18_T_datain = ( (|r_sys_processing_methodID) ? r_sub18_T_datain : 32'h0 ) ;
	assign w_sub18_T_r_w = ( (|r_sys_processing_methodID) ? r_sub18_T_r_w : 1'h0 ) ;
	assign w_sub18_U_addr = ( (|r_sys_processing_methodID) ? r_sub18_U_addr : 12'sh0 ) ;
	assign w_sub18_U_datain = ( (|r_sys_processing_methodID) ? r_sub18_U_datain : 32'h0 ) ;
	assign w_sub18_U_r_w = ( (|r_sys_processing_methodID) ? r_sub18_U_r_w : 1'h0 ) ;
	assign w_sub18_result_addr = ( (|r_sys_processing_methodID) ? r_sub18_result_addr : 12'sh0 ) ;
	assign w_sub18_result_datain = ( (|r_sys_processing_methodID) ? r_sub18_result_datain : 32'h0 ) ;
	assign w_sub18_result_r_w = ( (|r_sys_processing_methodID) ? r_sub18_result_r_w : 1'h0 ) ;
	assign w_sub17_T_addr = ( (|r_sys_processing_methodID) ? r_sub17_T_addr : 12'sh0 ) ;
	assign w_sub17_T_datain = ( (|r_sys_processing_methodID) ? r_sub17_T_datain : 32'h0 ) ;
	assign w_sub17_T_r_w = ( (|r_sys_processing_methodID) ? r_sub17_T_r_w : 1'h0 ) ;
	assign w_sub17_U_addr = ( (|r_sys_processing_methodID) ? r_sub17_U_addr : 12'sh0 ) ;
	assign w_sub17_U_datain = ( (|r_sys_processing_methodID) ? r_sub17_U_datain : 32'h0 ) ;
	assign w_sub17_U_r_w = ( (|r_sys_processing_methodID) ? r_sub17_U_r_w : 1'h0 ) ;
	assign w_sub17_result_addr = ( (|r_sys_processing_methodID) ? r_sub17_result_addr : 12'sh0 ) ;
	assign w_sub17_result_datain = ( (|r_sys_processing_methodID) ? r_sub17_result_datain : 32'h0 ) ;
	assign w_sub17_result_r_w = ( (|r_sys_processing_methodID) ? r_sub17_result_r_w : 1'h0 ) ;
	assign w_sub20_T_addr = ( (|r_sys_processing_methodID) ? r_sub20_T_addr : 12'sh0 ) ;
	assign w_sub20_T_datain = ( (|r_sys_processing_methodID) ? r_sub20_T_datain : 32'h0 ) ;
	assign w_sub20_T_r_w = ( (|r_sys_processing_methodID) ? r_sub20_T_r_w : 1'h0 ) ;
	assign w_sub20_U_addr = ( (|r_sys_processing_methodID) ? r_sub20_U_addr : 12'sh0 ) ;
	assign w_sub20_U_datain = ( (|r_sys_processing_methodID) ? r_sub20_U_datain : 32'h0 ) ;
	assign w_sub20_U_r_w = ( (|r_sys_processing_methodID) ? r_sub20_U_r_w : 1'h0 ) ;
	assign w_sub20_result_addr = ( (|r_sys_processing_methodID) ? r_sub20_result_addr : 12'sh0 ) ;
	assign w_sub20_result_datain = ( (|r_sys_processing_methodID) ? r_sub20_result_datain : 32'h0 ) ;
	assign w_sub20_result_r_w = ( (|r_sys_processing_methodID) ? r_sub20_result_r_w : 1'h0 ) ;
	assign w_sub21_T_addr = ( (|r_sys_processing_methodID) ? r_sub21_T_addr : 12'sh0 ) ;
	assign w_sub21_T_datain = ( (|r_sys_processing_methodID) ? r_sub21_T_datain : 32'h0 ) ;
	assign w_sub21_T_r_w = ( (|r_sys_processing_methodID) ? r_sub21_T_r_w : 1'h0 ) ;
	assign w_sub21_U_addr = ( (|r_sys_processing_methodID) ? r_sub21_U_addr : 12'sh0 ) ;
	assign w_sub21_U_datain = ( (|r_sys_processing_methodID) ? r_sub21_U_datain : 32'h0 ) ;
	assign w_sub21_U_r_w = ( (|r_sys_processing_methodID) ? r_sub21_U_r_w : 1'h0 ) ;
	assign w_sub21_result_addr = ( (|r_sys_processing_methodID) ? r_sub21_result_addr : 12'sh0 ) ;
	assign w_sub21_result_datain = ( (|r_sys_processing_methodID) ? r_sub21_result_datain : 32'h0 ) ;
	assign w_sub21_result_r_w = ( (|r_sys_processing_methodID) ? r_sub21_result_r_w : 1'h0 ) ;
	assign w_sub28_T_addr = ( (|r_sys_processing_methodID) ? r_sub28_T_addr : 12'sh0 ) ;
	assign w_sub28_T_datain = ( (|r_sys_processing_methodID) ? r_sub28_T_datain : 32'h0 ) ;
	assign w_sub28_T_r_w = ( (|r_sys_processing_methodID) ? r_sub28_T_r_w : 1'h0 ) ;
	assign w_sub28_U_addr = ( (|r_sys_processing_methodID) ? r_sub28_U_addr : 12'sh0 ) ;
	assign w_sub28_U_datain = ( (|r_sys_processing_methodID) ? r_sub28_U_datain : 32'h0 ) ;
	assign w_sub28_U_r_w = ( (|r_sys_processing_methodID) ? r_sub28_U_r_w : 1'h0 ) ;
	assign w_sub28_result_addr = ( (|r_sys_processing_methodID) ? r_sub28_result_addr : 12'sh0 ) ;
	assign w_sub28_result_datain = ( (|r_sys_processing_methodID) ? r_sub28_result_datain : 32'h0 ) ;
	assign w_sub28_result_r_w = ( (|r_sys_processing_methodID) ? r_sub28_result_r_w : 1'h0 ) ;
	assign w_sub29_T_addr = ( (|r_sys_processing_methodID) ? r_sub29_T_addr : 12'sh0 ) ;
	assign w_sub29_T_datain = ( (|r_sys_processing_methodID) ? r_sub29_T_datain : 32'h0 ) ;
	assign w_sub29_T_r_w = ( (|r_sys_processing_methodID) ? r_sub29_T_r_w : 1'h0 ) ;
	assign w_sub29_U_addr = ( (|r_sys_processing_methodID) ? r_sub29_U_addr : 12'sh0 ) ;
	assign w_sub29_U_datain = ( (|r_sys_processing_methodID) ? r_sub29_U_datain : 32'h0 ) ;
	assign w_sub29_U_r_w = ( (|r_sys_processing_methodID) ? r_sub29_U_r_w : 1'h0 ) ;
	assign w_sub29_result_addr = ( (|r_sys_processing_methodID) ? r_sub29_result_addr : 12'sh0 ) ;
	assign w_sub29_result_datain = ( (|r_sys_processing_methodID) ? r_sub29_result_datain : 32'h0 ) ;
	assign w_sub29_result_r_w = ( (|r_sys_processing_methodID) ? r_sub29_result_r_w : 1'h0 ) ;
	assign w_sub26_T_addr = ( (|r_sys_processing_methodID) ? r_sub26_T_addr : 12'sh0 ) ;
	assign w_sub26_T_datain = ( (|r_sys_processing_methodID) ? r_sub26_T_datain : 32'h0 ) ;
	assign w_sub26_T_r_w = ( (|r_sys_processing_methodID) ? r_sub26_T_r_w : 1'h0 ) ;
	assign w_sub26_U_addr = ( (|r_sys_processing_methodID) ? r_sub26_U_addr : 12'sh0 ) ;
	assign w_sub26_U_datain = ( (|r_sys_processing_methodID) ? r_sub26_U_datain : 32'h0 ) ;
	assign w_sub26_U_r_w = ( (|r_sys_processing_methodID) ? r_sub26_U_r_w : 1'h0 ) ;
	assign w_sub26_result_addr = ( (|r_sys_processing_methodID) ? r_sub26_result_addr : 12'sh0 ) ;
	assign w_sub26_result_datain = ( (|r_sys_processing_methodID) ? r_sub26_result_datain : 32'h0 ) ;
	assign w_sub26_result_r_w = ( (|r_sys_processing_methodID) ? r_sub26_result_r_w : 1'h0 ) ;
	assign w_sub09_T_addr = ( (|r_sys_processing_methodID) ? r_sub09_T_addr : 12'sh0 ) ;
	assign w_sub09_T_datain = ( (|r_sys_processing_methodID) ? r_sub09_T_datain : 32'h0 ) ;
	assign w_sub09_T_r_w = ( (|r_sys_processing_methodID) ? r_sub09_T_r_w : 1'h0 ) ;
	assign w_sub09_U_addr = ( (|r_sys_processing_methodID) ? r_sub09_U_addr : 12'sh0 ) ;
	assign w_sub09_U_datain = ( (|r_sys_processing_methodID) ? r_sub09_U_datain : 32'h0 ) ;
	assign w_sub09_U_r_w = ( (|r_sys_processing_methodID) ? r_sub09_U_r_w : 1'h0 ) ;
	assign w_sub09_result_addr = ( (|r_sys_processing_methodID) ? r_sub09_result_addr : 12'sh0 ) ;
	assign w_sub09_result_datain = ( (|r_sys_processing_methodID) ? r_sub09_result_datain : 32'h0 ) ;
	assign w_sub09_result_r_w = ( (|r_sys_processing_methodID) ? r_sub09_result_r_w : 1'h0 ) ;
	assign w_sub27_T_addr = ( (|r_sys_processing_methodID) ? r_sub27_T_addr : 12'sh0 ) ;
	assign w_sub27_T_datain = ( (|r_sys_processing_methodID) ? r_sub27_T_datain : 32'h0 ) ;
	assign w_sub27_T_r_w = ( (|r_sys_processing_methodID) ? r_sub27_T_r_w : 1'h0 ) ;
	assign w_sub27_U_addr = ( (|r_sys_processing_methodID) ? r_sub27_U_addr : 12'sh0 ) ;
	assign w_sub27_U_datain = ( (|r_sys_processing_methodID) ? r_sub27_U_datain : 32'h0 ) ;
	assign w_sub27_U_r_w = ( (|r_sys_processing_methodID) ? r_sub27_U_r_w : 1'h0 ) ;
	assign w_sub27_result_addr = ( (|r_sys_processing_methodID) ? r_sub27_result_addr : 12'sh0 ) ;
	assign w_sub27_result_datain = ( (|r_sys_processing_methodID) ? r_sub27_result_datain : 32'h0 ) ;
	assign w_sub27_result_r_w = ( (|r_sys_processing_methodID) ? r_sub27_result_r_w : 1'h0 ) ;
	assign w_sub08_T_addr = ( (|r_sys_processing_methodID) ? r_sub08_T_addr : 12'sh0 ) ;
	assign w_sub08_T_datain = ( (|r_sys_processing_methodID) ? r_sub08_T_datain : 32'h0 ) ;
	assign w_sub08_T_r_w = ( (|r_sys_processing_methodID) ? r_sub08_T_r_w : 1'h0 ) ;
	assign w_sub08_U_addr = ( (|r_sys_processing_methodID) ? r_sub08_U_addr : 12'sh0 ) ;
	assign w_sub08_U_datain = ( (|r_sys_processing_methodID) ? r_sub08_U_datain : 32'h0 ) ;
	assign w_sub08_U_r_w = ( (|r_sys_processing_methodID) ? r_sub08_U_r_w : 1'h0 ) ;
	assign w_sub08_result_addr = ( (|r_sys_processing_methodID) ? r_sub08_result_addr : 12'sh0 ) ;
	assign w_sub08_result_datain = ( (|r_sys_processing_methodID) ? r_sub08_result_datain : 32'h0 ) ;
	assign w_sub08_result_r_w = ( (|r_sys_processing_methodID) ? r_sub08_result_r_w : 1'h0 ) ;
	assign w_sub24_T_addr = ( (|r_sys_processing_methodID) ? r_sub24_T_addr : 12'sh0 ) ;
	assign w_sub24_T_datain = ( (|r_sys_processing_methodID) ? r_sub24_T_datain : 32'h0 ) ;
	assign w_sub24_T_r_w = ( (|r_sys_processing_methodID) ? r_sub24_T_r_w : 1'h0 ) ;
	assign w_sub24_U_addr = ( (|r_sys_processing_methodID) ? r_sub24_U_addr : 12'sh0 ) ;
	assign w_sub24_U_datain = ( (|r_sys_processing_methodID) ? r_sub24_U_datain : 32'h0 ) ;
	assign w_sub24_U_r_w = ( (|r_sys_processing_methodID) ? r_sub24_U_r_w : 1'h0 ) ;
	assign w_sub24_result_addr = ( (|r_sys_processing_methodID) ? r_sub24_result_addr : 12'sh0 ) ;
	assign w_sub24_result_datain = ( (|r_sys_processing_methodID) ? r_sub24_result_datain : 32'h0 ) ;
	assign w_sub24_result_r_w = ( (|r_sys_processing_methodID) ? r_sub24_result_r_w : 1'h0 ) ;
	assign w_sub25_T_addr = ( (|r_sys_processing_methodID) ? r_sub25_T_addr : 12'sh0 ) ;
	assign w_sub25_T_datain = ( (|r_sys_processing_methodID) ? r_sub25_T_datain : 32'h0 ) ;
	assign w_sub25_T_r_w = ( (|r_sys_processing_methodID) ? r_sub25_T_r_w : 1'h0 ) ;
	assign w_sub25_U_addr = ( (|r_sys_processing_methodID) ? r_sub25_U_addr : 12'sh0 ) ;
	assign w_sub25_U_datain = ( (|r_sys_processing_methodID) ? r_sub25_U_datain : 32'h0 ) ;
	assign w_sub25_U_r_w = ( (|r_sys_processing_methodID) ? r_sub25_U_r_w : 1'h0 ) ;
	assign w_sub25_result_addr = ( (|r_sys_processing_methodID) ? r_sub25_result_addr : 12'sh0 ) ;
	assign w_sub25_result_datain = ( (|r_sys_processing_methodID) ? r_sub25_result_datain : 32'h0 ) ;
	assign w_sub25_result_r_w = ( (|r_sys_processing_methodID) ? r_sub25_result_r_w : 1'h0 ) ;
	assign w_sub22_T_addr = ( (|r_sys_processing_methodID) ? r_sub22_T_addr : 12'sh0 ) ;
	assign w_sub22_T_datain = ( (|r_sys_processing_methodID) ? r_sub22_T_datain : 32'h0 ) ;
	assign w_sub22_T_r_w = ( (|r_sys_processing_methodID) ? r_sub22_T_r_w : 1'h0 ) ;
	assign w_sub22_U_addr = ( (|r_sys_processing_methodID) ? r_sub22_U_addr : 12'sh0 ) ;
	assign w_sub22_U_datain = ( (|r_sys_processing_methodID) ? r_sub22_U_datain : 32'h0 ) ;
	assign w_sub22_U_r_w = ( (|r_sys_processing_methodID) ? r_sub22_U_r_w : 1'h0 ) ;
	assign w_sub22_result_addr = ( (|r_sys_processing_methodID) ? r_sub22_result_addr : 12'sh0 ) ;
	assign w_sub22_result_datain = ( (|r_sys_processing_methodID) ? r_sub22_result_datain : 32'h0 ) ;
	assign w_sub22_result_r_w = ( (|r_sys_processing_methodID) ? r_sub22_result_r_w : 1'h0 ) ;
	assign w_sub23_T_addr = ( (|r_sys_processing_methodID) ? r_sub23_T_addr : 12'sh0 ) ;
	assign w_sub23_T_datain = ( (|r_sys_processing_methodID) ? r_sub23_T_datain : 32'h0 ) ;
	assign w_sub23_T_r_w = ( (|r_sys_processing_methodID) ? r_sub23_T_r_w : 1'h0 ) ;
	assign w_sub23_U_addr = ( (|r_sys_processing_methodID) ? r_sub23_U_addr : 12'sh0 ) ;
	assign w_sub23_U_datain = ( (|r_sys_processing_methodID) ? r_sub23_U_datain : 32'h0 ) ;
	assign w_sub23_U_r_w = ( (|r_sys_processing_methodID) ? r_sub23_U_r_w : 1'h0 ) ;
	assign w_sub23_result_addr = ( (|r_sys_processing_methodID) ? r_sub23_result_addr : 12'sh0 ) ;
	assign w_sub23_result_datain = ( (|r_sys_processing_methodID) ? r_sub23_result_datain : 32'h0 ) ;
	assign w_sub23_result_r_w = ( (|r_sys_processing_methodID) ? r_sub23_result_r_w : 1'h0 ) ;
	assign w_sub03_T_addr = ( (|r_sys_processing_methodID) ? r_sub03_T_addr : 12'sh0 ) ;
	assign w_sub03_T_datain = ( (|r_sys_processing_methodID) ? r_sub03_T_datain : 32'h0 ) ;
	assign w_sub03_T_r_w = ( (|r_sys_processing_methodID) ? r_sub03_T_r_w : 1'h0 ) ;
	assign w_sub03_U_addr = ( (|r_sys_processing_methodID) ? r_sub03_U_addr : 12'sh0 ) ;
	assign w_sub03_U_datain = ( (|r_sys_processing_methodID) ? r_sub03_U_datain : 32'h0 ) ;
	assign w_sub03_U_r_w = ( (|r_sys_processing_methodID) ? r_sub03_U_r_w : 1'h0 ) ;
	assign w_sub03_result_addr = ( (|r_sys_processing_methodID) ? r_sub03_result_addr : 12'sh0 ) ;
	assign w_sub03_result_datain = ( (|r_sys_processing_methodID) ? r_sub03_result_datain : 32'h0 ) ;
	assign w_sub03_result_r_w = ( (|r_sys_processing_methodID) ? r_sub03_result_r_w : 1'h0 ) ;
	assign w_sub02_T_addr = ( (|r_sys_processing_methodID) ? r_sub02_T_addr : 12'sh0 ) ;
	assign w_sub02_T_datain = ( (|r_sys_processing_methodID) ? r_sub02_T_datain : 32'h0 ) ;
	assign w_sub02_T_r_w = ( (|r_sys_processing_methodID) ? r_sub02_T_r_w : 1'h0 ) ;
	assign w_sub02_U_addr = ( (|r_sys_processing_methodID) ? r_sub02_U_addr : 12'sh0 ) ;
	assign w_sub02_U_datain = ( (|r_sys_processing_methodID) ? r_sub02_U_datain : 32'h0 ) ;
	assign w_sub02_U_r_w = ( (|r_sys_processing_methodID) ? r_sub02_U_r_w : 1'h0 ) ;
	assign w_sub02_result_addr = ( (|r_sys_processing_methodID) ? r_sub02_result_addr : 12'sh0 ) ;
	assign w_sub02_result_datain = ( (|r_sys_processing_methodID) ? r_sub02_result_datain : 32'h0 ) ;
	assign w_sub02_result_r_w = ( (|r_sys_processing_methodID) ? r_sub02_result_r_w : 1'h0 ) ;
	assign w_sub01_T_addr = ( (|r_sys_processing_methodID) ? r_sub01_T_addr : 12'sh0 ) ;
	assign w_sub01_T_datain = ( (|r_sys_processing_methodID) ? r_sub01_T_datain : 32'h0 ) ;
	assign w_sub01_T_r_w = ( (|r_sys_processing_methodID) ? r_sub01_T_r_w : 1'h0 ) ;
	assign w_sub01_U_addr = ( (|r_sys_processing_methodID) ? r_sub01_U_addr : 12'sh0 ) ;
	assign w_sub01_U_datain = ( (|r_sys_processing_methodID) ? r_sub01_U_datain : 32'h0 ) ;
	assign w_sub01_U_r_w = ( (|r_sys_processing_methodID) ? r_sub01_U_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 12'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub00_T_addr = ( (|r_sys_processing_methodID) ? r_sub00_T_addr : 12'sh0 ) ;
	assign w_sub00_T_datain = ( (|r_sys_processing_methodID) ? r_sub00_T_datain : 32'h0 ) ;
	assign w_sub00_T_r_w = ( (|r_sys_processing_methodID) ? r_sub00_T_r_w : 1'h0 ) ;
	assign w_sub00_U_addr = ( (|r_sys_processing_methodID) ? r_sub00_U_addr : 12'sh0 ) ;
	assign w_sub00_U_datain = ( (|r_sys_processing_methodID) ? r_sub00_U_datain : 32'h0 ) ;
	assign w_sub00_U_r_w = ( (|r_sys_processing_methodID) ? r_sub00_U_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 12'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sub07_T_addr = ( (|r_sys_processing_methodID) ? r_sub07_T_addr : 12'sh0 ) ;
	assign w_sub07_T_datain = ( (|r_sys_processing_methodID) ? r_sub07_T_datain : 32'h0 ) ;
	assign w_sub07_T_r_w = ( (|r_sys_processing_methodID) ? r_sub07_T_r_w : 1'h0 ) ;
	assign w_sub07_U_addr = ( (|r_sys_processing_methodID) ? r_sub07_U_addr : 12'sh0 ) ;
	assign w_sub07_U_datain = ( (|r_sys_processing_methodID) ? r_sub07_U_datain : 32'h0 ) ;
	assign w_sub07_U_r_w = ( (|r_sys_processing_methodID) ? r_sub07_U_r_w : 1'h0 ) ;
	assign w_sub07_result_addr = ( (|r_sys_processing_methodID) ? r_sub07_result_addr : 12'sh0 ) ;
	assign w_sub07_result_datain = ( (|r_sys_processing_methodID) ? r_sub07_result_datain : 32'h0 ) ;
	assign w_sub07_result_r_w = ( (|r_sys_processing_methodID) ? r_sub07_result_r_w : 1'h0 ) ;
	assign w_sub06_T_addr = ( (|r_sys_processing_methodID) ? r_sub06_T_addr : 12'sh0 ) ;
	assign w_sub06_T_datain = ( (|r_sys_processing_methodID) ? r_sub06_T_datain : 32'h0 ) ;
	assign w_sub06_T_r_w = ( (|r_sys_processing_methodID) ? r_sub06_T_r_w : 1'h0 ) ;
	assign w_sub06_U_addr = ( (|r_sys_processing_methodID) ? r_sub06_U_addr : 12'sh0 ) ;
	assign w_sub06_U_datain = ( (|r_sys_processing_methodID) ? r_sub06_U_datain : 32'h0 ) ;
	assign w_sub06_U_r_w = ( (|r_sys_processing_methodID) ? r_sub06_U_r_w : 1'h0 ) ;
	assign w_sub06_result_addr = ( (|r_sys_processing_methodID) ? r_sub06_result_addr : 12'sh0 ) ;
	assign w_sub06_result_datain = ( (|r_sys_processing_methodID) ? r_sub06_result_datain : 32'h0 ) ;
	assign w_sub06_result_r_w = ( (|r_sys_processing_methodID) ? r_sub06_result_r_w : 1'h0 ) ;
	assign w_sub05_T_addr = ( (|r_sys_processing_methodID) ? r_sub05_T_addr : 12'sh0 ) ;
	assign w_sub05_T_datain = ( (|r_sys_processing_methodID) ? r_sub05_T_datain : 32'h0 ) ;
	assign w_sub05_T_r_w = ( (|r_sys_processing_methodID) ? r_sub05_T_r_w : 1'h0 ) ;
	assign w_sub05_U_addr = ( (|r_sys_processing_methodID) ? r_sub05_U_addr : 12'sh0 ) ;
	assign w_sub05_U_datain = ( (|r_sys_processing_methodID) ? r_sub05_U_datain : 32'h0 ) ;
	assign w_sub05_U_r_w = ( (|r_sys_processing_methodID) ? r_sub05_U_r_w : 1'h0 ) ;
	assign w_sub05_result_addr = ( (|r_sys_processing_methodID) ? r_sub05_result_addr : 12'sh0 ) ;
	assign w_sub05_result_datain = ( (|r_sys_processing_methodID) ? r_sub05_result_datain : 32'h0 ) ;
	assign w_sub05_result_r_w = ( (|r_sys_processing_methodID) ? r_sub05_result_r_w : 1'h0 ) ;
	assign w_sub04_T_addr = ( (|r_sys_processing_methodID) ? r_sub04_T_addr : 12'sh0 ) ;
	assign w_sub04_T_datain = ( (|r_sys_processing_methodID) ? r_sub04_T_datain : 32'h0 ) ;
	assign w_sub04_T_r_w = ( (|r_sys_processing_methodID) ? r_sub04_T_r_w : 1'h0 ) ;
	assign w_sub04_U_addr = ( (|r_sys_processing_methodID) ? r_sub04_U_addr : 12'sh0 ) ;
	assign w_sub04_U_datain = ( (|r_sys_processing_methodID) ? r_sub04_U_datain : 32'h0 ) ;
	assign w_sub04_U_r_w = ( (|r_sys_processing_methodID) ? r_sub04_U_r_w : 1'h0 ) ;
	assign w_sub04_result_addr = ( (|r_sys_processing_methodID) ? r_sub04_result_addr : 12'sh0 ) ;
	assign w_sub04_result_datain = ( (|r_sys_processing_methodID) ? r_sub04_result_datain : 32'h0 ) ;
	assign w_sub04_result_r_w = ( (|r_sys_processing_methodID) ? r_sub04_result_r_w : 1'h0 ) ;
	assign w_sub10_T_addr = ( (|r_sys_processing_methodID) ? r_sub10_T_addr : 12'sh0 ) ;
	assign w_sub10_T_datain = ( (|r_sys_processing_methodID) ? r_sub10_T_datain : 32'h0 ) ;
	assign w_sub10_T_r_w = ( (|r_sys_processing_methodID) ? r_sub10_T_r_w : 1'h0 ) ;
	assign w_sub10_U_addr = ( (|r_sys_processing_methodID) ? r_sub10_U_addr : 12'sh0 ) ;
	assign w_sub10_U_datain = ( (|r_sys_processing_methodID) ? r_sub10_U_datain : 32'h0 ) ;
	assign w_sub10_U_r_w = ( (|r_sys_processing_methodID) ? r_sub10_U_r_w : 1'h0 ) ;
	assign w_sub10_result_addr = ( (|r_sys_processing_methodID) ? r_sub10_result_addr : 12'sh0 ) ;
	assign w_sub10_result_datain = ( (|r_sys_processing_methodID) ? r_sub10_result_datain : 32'h0 ) ;
	assign w_sub10_result_r_w = ( (|r_sys_processing_methodID) ? r_sub10_result_r_w : 1'h0 ) ;
	assign w_sub31_T_addr = ( (|r_sys_processing_methodID) ? r_sub31_T_addr : 12'sh0 ) ;
	assign w_sub31_T_datain = ( (|r_sys_processing_methodID) ? r_sub31_T_datain : 32'h0 ) ;
	assign w_sub31_T_r_w = ( (|r_sys_processing_methodID) ? r_sub31_T_r_w : 1'h0 ) ;
	assign w_sub31_U_addr = ( (|r_sys_processing_methodID) ? r_sub31_U_addr : 12'sh0 ) ;
	assign w_sub31_U_datain = ( (|r_sys_processing_methodID) ? r_sub31_U_datain : 32'h0 ) ;
	assign w_sub31_U_r_w = ( (|r_sys_processing_methodID) ? r_sub31_U_r_w : 1'h0 ) ;
	assign w_sub31_result_addr = ( (|r_sys_processing_methodID) ? r_sub31_result_addr : 12'sh0 ) ;
	assign w_sub31_result_datain = ( (|r_sys_processing_methodID) ? r_sub31_result_datain : 32'h0 ) ;
	assign w_sub31_result_r_w = ( (|r_sys_processing_methodID) ? r_sub31_result_r_w : 1'h0 ) ;
	assign w_sub30_T_addr = ( (|r_sys_processing_methodID) ? r_sub30_T_addr : 12'sh0 ) ;
	assign w_sub30_T_datain = ( (|r_sys_processing_methodID) ? r_sub30_T_datain : 32'h0 ) ;
	assign w_sub30_T_r_w = ( (|r_sys_processing_methodID) ? r_sub30_T_r_w : 1'h0 ) ;
	assign w_sub30_U_addr = ( (|r_sys_processing_methodID) ? r_sub30_U_addr : 12'sh0 ) ;
	assign w_sub30_U_datain = ( (|r_sys_processing_methodID) ? r_sub30_U_datain : 32'h0 ) ;
	assign w_sub30_U_r_w = ( (|r_sys_processing_methodID) ? r_sub30_U_r_w : 1'h0 ) ;
	assign w_sub30_result_addr = ( (|r_sys_processing_methodID) ? r_sub30_result_addr : 12'sh0 ) ;
	assign w_sub30_result_datain = ( (|r_sys_processing_methodID) ? r_sub30_result_datain : 32'h0 ) ;
	assign w_sub30_result_r_w = ( (|r_sys_processing_methodID) ? r_sub30_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh00000080;
	assign w_sys_tmp3 = 32'sh00000081;
	assign w_sys_tmp5 = 32'h3a03126f;
	assign w_sys_tmp6 = 32'h3d000000;
	assign w_sys_tmp7 = 32'h3c000000;
	assign w_sys_tmp8 = 32'h3c03126f;
	assign w_sys_tmp9 = 32'h3d03126f;
	assign w_sys_tmp10 = 32'h3f03126f;
	assign w_sys_tmp11 = 32'h4103126f;
	assign w_sys_tmp12 = ( !w_sys_tmp13 );
	assign w_sys_tmp13 = (r_run_my_39 < r_run_k_35);
	assign w_sys_tmp14 = (r_run_k_35 + w_sys_intOne);
	assign w_sys_tmp15 = ( !w_sys_tmp16 );
	assign w_sys_tmp16 = (r_run_mx_38 < r_run_j_36);
	assign w_sys_tmp18 = w_ip_MultFloat_product_0;
	assign w_sys_tmp19 = w_ip_FixedToFloat_floating_0;
	assign w_sys_tmp20 = (r_run_k_35 - w_sys_intOne);
	assign w_sys_tmp22 = (w_sys_tmp23 + r_run_k_35);
	assign w_sys_tmp23 = (r_run_j_36 * w_sys_tmp24);
	assign w_sys_tmp24 = 32'sh00000081;
	assign w_sys_tmp25 = 32'h0;
	assign w_sys_tmp27 = (w_sys_tmp28 + r_run_k_35);
	assign w_sys_tmp28 = (r_run_copy1_j_53 * w_sys_tmp24);
	assign w_sys_tmp32 = (w_sys_tmp33 + r_run_k_35);
	assign w_sys_tmp33 = (r_run_copy0_j_52 * w_sys_tmp24);
	assign w_sys_tmp36 = 32'h42200000;
	assign w_sys_tmp37 = w_sys_tmp18;
	assign w_sys_tmp38 = 32'h3f800000;
	assign w_sys_tmp40 = (r_run_copy0_j_52 + w_sys_intOne);
	assign w_sys_tmp41 = (r_run_copy1_j_53 + w_sys_intOne);
	assign w_sys_tmp42 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp110 = r_sys_tmp4_float;
	assign w_sys_tmp184 = ( !w_sys_tmp185 );
	assign w_sys_tmp185 = (w_sys_tmp186 < r_run_k_35);
	assign w_sys_tmp186 = 32'sh00000081;
	assign w_sys_tmp189 = (w_sys_tmp190 + r_run_k_35);
	assign w_sys_tmp190 = 32'sh00000081;
	assign w_sys_tmp191 = 32'h0;
	assign w_sys_tmp193 = (w_sys_tmp194 + r_run_k_35);
	assign w_sys_tmp194 = (r_run_mx_38 * w_sys_tmp190);
	assign w_sys_tmp196 = w_fld_T_0_dataout_1;
	assign w_sys_tmp197 = (w_sys_tmp198 + r_run_k_35);
	assign w_sys_tmp198 = (w_sys_tmp199 * w_sys_tmp190);
	assign w_sys_tmp199 = (r_run_mx_38 - w_sys_intOne);
	assign w_sys_tmp201 = (r_run_k_35 + w_sys_intOne);
	assign w_sys_tmp202 = ( !w_sys_tmp203 );
	assign w_sys_tmp203 = (w_sys_tmp204 < r_run_j_36);
	assign w_sys_tmp204 = 32'sh00000081;
	assign w_sys_tmp207 = (w_sys_tmp208 + w_sys_intOne);
	assign w_sys_tmp208 = (r_run_j_36 * w_sys_tmp209);
	assign w_sys_tmp209 = 32'sh00000081;
	assign w_sys_tmp210 = 32'h0;
	assign w_sys_tmp212 = (w_sys_tmp213 + r_run_my_39);
	assign w_sys_tmp213 = (r_run_copy0_j_54 * w_sys_tmp209);
	assign w_sys_tmp216 = (r_run_copy0_j_54 + w_sys_intOne);
	assign w_sys_tmp217 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp290 = (r_run_mx_38 / w_sys_tmp291);
	assign w_sys_tmp291 = 32'sh00000004;
	assign w_sys_tmp292 = ( !w_sys_tmp293 );
	assign w_sys_tmp293 = (w_sys_tmp294 < r_run_j_36);
	assign w_sys_tmp294 = (r_run_mx_38 / w_sys_tmp295);
	assign w_sys_tmp295 = 32'sh00000002;
	assign w_sys_tmp298 = (w_sys_tmp299 + w_sys_intOne);
	assign w_sys_tmp299 = (r_run_j_36 * w_sys_tmp300);
	assign w_sys_tmp300 = 32'sh00000081;
	assign w_sys_tmp301 = 32'h3f800000;
	assign w_sys_tmp302 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp339 = ( !w_sys_tmp340 );
	assign w_sys_tmp340 = (w_sys_tmp341 < r_run_k_35);
	assign w_sys_tmp341 = 32'sh00000021;
	assign w_sys_tmp342 = (r_run_k_35 + w_sys_intOne);
	assign w_sys_tmp343 = ( !w_sys_tmp344 );
	assign w_sys_tmp344 = (w_sys_tmp345 < r_run_j_36);
	assign w_sys_tmp345 = 32'sh00000011;
	assign w_sys_tmp348 = (w_sys_tmp349 + r_run_k_35);
	assign w_sys_tmp349 = (r_run_j_36 * w_sys_tmp350);
	assign w_sys_tmp350 = 32'sh00000081;
	assign w_sys_tmp351 = w_fld_U_2_dataout_1;
	assign w_sys_tmp352 = (w_sys_tmp353 + r_run_k_35);
	assign w_sys_tmp353 = (r_run_copy2_j_57 * w_sys_tmp350);
	assign w_sys_tmp356 = (w_sys_tmp357 + r_run_k_35);
	assign w_sys_tmp357 = (r_run_copy1_j_56 * w_sys_tmp350);
	assign w_sys_tmp359 = w_fld_T_0_dataout_1;
	assign w_sys_tmp360 = (w_sys_tmp361 + r_run_k_35);
	assign w_sys_tmp361 = (r_run_copy0_j_55 * w_sys_tmp350);
	assign w_sys_tmp363 = (r_run_copy0_j_55 + w_sys_intOne);
	assign w_sys_tmp364 = (r_run_copy1_j_56 + w_sys_intOne);
	assign w_sys_tmp365 = (r_run_copy2_j_57 + w_sys_intOne);
	assign w_sys_tmp366 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp487 = 32'sh00000010;
	assign w_sys_tmp488 = ( !w_sys_tmp489 );
	assign w_sys_tmp489 = (w_sys_tmp490 < r_run_j_36);
	assign w_sys_tmp490 = 32'sh00000021;
	assign w_sys_tmp493 = (w_sys_tmp494 + r_run_k_35);
	assign w_sys_tmp494 = (r_run_j_36 * w_sys_tmp495);
	assign w_sys_tmp495 = 32'sh00000081;
	assign w_sys_tmp496 = w_fld_U_2_dataout_1;
	assign w_sys_tmp497 = (w_sys_tmp498 + r_run_k_35);
	assign w_sys_tmp498 = (r_run_copy2_j_60 * w_sys_tmp495);
	assign w_sys_tmp501 = (w_sys_tmp502 + r_run_k_35);
	assign w_sys_tmp502 = (r_run_copy1_j_59 * w_sys_tmp495);
	assign w_sys_tmp504 = w_fld_T_0_dataout_1;
	assign w_sys_tmp505 = (w_sys_tmp506 + r_run_k_35);
	assign w_sys_tmp506 = (r_run_copy0_j_58 * w_sys_tmp495);
	assign w_sys_tmp508 = (r_run_copy0_j_58 + w_sys_intOne);
	assign w_sys_tmp509 = (r_run_copy1_j_59 + w_sys_intOne);
	assign w_sys_tmp510 = (r_run_copy2_j_60 + w_sys_intOne);
	assign w_sys_tmp511 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp632 = 32'sh00000020;
	assign w_sys_tmp633 = ( !w_sys_tmp634 );
	assign w_sys_tmp634 = (w_sys_tmp635 < r_run_j_36);
	assign w_sys_tmp635 = 32'sh00000031;
	assign w_sys_tmp638 = (w_sys_tmp639 + r_run_k_35);
	assign w_sys_tmp639 = (r_run_j_36 * w_sys_tmp640);
	assign w_sys_tmp640 = 32'sh00000081;
	assign w_sys_tmp641 = w_fld_U_2_dataout_1;
	assign w_sys_tmp642 = (w_sys_tmp643 + r_run_k_35);
	assign w_sys_tmp643 = (r_run_copy2_j_63 * w_sys_tmp640);
	assign w_sys_tmp646 = (w_sys_tmp647 + r_run_k_35);
	assign w_sys_tmp647 = (r_run_copy1_j_62 * w_sys_tmp640);
	assign w_sys_tmp649 = w_fld_T_0_dataout_1;
	assign w_sys_tmp650 = (w_sys_tmp651 + r_run_k_35);
	assign w_sys_tmp651 = (r_run_copy0_j_61 * w_sys_tmp640);
	assign w_sys_tmp653 = (r_run_copy0_j_61 + w_sys_intOne);
	assign w_sys_tmp654 = (r_run_copy1_j_62 + w_sys_intOne);
	assign w_sys_tmp655 = (r_run_copy2_j_63 + w_sys_intOne);
	assign w_sys_tmp656 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp777 = 32'sh00000030;
	assign w_sys_tmp778 = ( !w_sys_tmp779 );
	assign w_sys_tmp779 = (w_sys_tmp780 < r_run_j_36);
	assign w_sys_tmp780 = 32'sh00000041;
	assign w_sys_tmp783 = (w_sys_tmp784 + r_run_k_35);
	assign w_sys_tmp784 = (r_run_j_36 * w_sys_tmp785);
	assign w_sys_tmp785 = 32'sh00000081;
	assign w_sys_tmp786 = w_fld_U_2_dataout_1;
	assign w_sys_tmp787 = (w_sys_tmp788 + r_run_k_35);
	assign w_sys_tmp788 = (r_run_copy2_j_66 * w_sys_tmp785);
	assign w_sys_tmp791 = (w_sys_tmp792 + r_run_k_35);
	assign w_sys_tmp792 = (r_run_copy1_j_65 * w_sys_tmp785);
	assign w_sys_tmp794 = w_fld_T_0_dataout_1;
	assign w_sys_tmp795 = (w_sys_tmp796 + r_run_k_35);
	assign w_sys_tmp796 = (r_run_copy0_j_64 * w_sys_tmp785);
	assign w_sys_tmp798 = (r_run_copy0_j_64 + w_sys_intOne);
	assign w_sys_tmp799 = (r_run_copy1_j_65 + w_sys_intOne);
	assign w_sys_tmp800 = (r_run_copy2_j_66 + w_sys_intOne);
	assign w_sys_tmp801 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp922 = 32'sh00000040;
	assign w_sys_tmp923 = ( !w_sys_tmp924 );
	assign w_sys_tmp924 = (w_sys_tmp925 < r_run_j_36);
	assign w_sys_tmp925 = 32'sh00000051;
	assign w_sys_tmp928 = (w_sys_tmp929 + r_run_k_35);
	assign w_sys_tmp929 = (r_run_j_36 * w_sys_tmp930);
	assign w_sys_tmp930 = 32'sh00000081;
	assign w_sys_tmp931 = w_fld_U_2_dataout_1;
	assign w_sys_tmp932 = (w_sys_tmp933 + r_run_k_35);
	assign w_sys_tmp933 = (r_run_copy2_j_69 * w_sys_tmp930);
	assign w_sys_tmp936 = (w_sys_tmp937 + r_run_k_35);
	assign w_sys_tmp937 = (r_run_copy1_j_68 * w_sys_tmp930);
	assign w_sys_tmp939 = w_fld_T_0_dataout_1;
	assign w_sys_tmp940 = (w_sys_tmp941 + r_run_k_35);
	assign w_sys_tmp941 = (r_run_copy0_j_67 * w_sys_tmp930);
	assign w_sys_tmp943 = (r_run_copy0_j_67 + w_sys_intOne);
	assign w_sys_tmp944 = (r_run_copy1_j_68 + w_sys_intOne);
	assign w_sys_tmp945 = (r_run_copy2_j_69 + w_sys_intOne);
	assign w_sys_tmp946 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp1067 = 32'sh00000050;
	assign w_sys_tmp1068 = ( !w_sys_tmp1069 );
	assign w_sys_tmp1069 = (w_sys_tmp1070 < r_run_j_36);
	assign w_sys_tmp1070 = 32'sh00000061;
	assign w_sys_tmp1073 = (w_sys_tmp1074 + r_run_k_35);
	assign w_sys_tmp1074 = (r_run_j_36 * w_sys_tmp1075);
	assign w_sys_tmp1075 = 32'sh00000081;
	assign w_sys_tmp1076 = w_fld_U_2_dataout_1;
	assign w_sys_tmp1077 = (w_sys_tmp1078 + r_run_k_35);
	assign w_sys_tmp1078 = (r_run_copy2_j_72 * w_sys_tmp1075);
	assign w_sys_tmp1081 = (w_sys_tmp1082 + r_run_k_35);
	assign w_sys_tmp1082 = (r_run_copy1_j_71 * w_sys_tmp1075);
	assign w_sys_tmp1084 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1085 = (w_sys_tmp1086 + r_run_k_35);
	assign w_sys_tmp1086 = (r_run_copy0_j_70 * w_sys_tmp1075);
	assign w_sys_tmp1088 = (r_run_copy0_j_70 + w_sys_intOne);
	assign w_sys_tmp1089 = (r_run_copy1_j_71 + w_sys_intOne);
	assign w_sys_tmp1090 = (r_run_copy2_j_72 + w_sys_intOne);
	assign w_sys_tmp1091 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp1212 = 32'sh00000060;
	assign w_sys_tmp1213 = ( !w_sys_tmp1214 );
	assign w_sys_tmp1214 = (w_sys_tmp1215 < r_run_j_36);
	assign w_sys_tmp1215 = 32'sh00000071;
	assign w_sys_tmp1218 = (w_sys_tmp1219 + r_run_k_35);
	assign w_sys_tmp1219 = (r_run_j_36 * w_sys_tmp1220);
	assign w_sys_tmp1220 = 32'sh00000081;
	assign w_sys_tmp1221 = w_fld_U_2_dataout_1;
	assign w_sys_tmp1222 = (w_sys_tmp1223 + r_run_k_35);
	assign w_sys_tmp1223 = (r_run_copy2_j_75 * w_sys_tmp1220);
	assign w_sys_tmp1226 = (w_sys_tmp1227 + r_run_k_35);
	assign w_sys_tmp1227 = (r_run_copy1_j_74 * w_sys_tmp1220);
	assign w_sys_tmp1229 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1230 = (w_sys_tmp1231 + r_run_k_35);
	assign w_sys_tmp1231 = (r_run_copy0_j_73 * w_sys_tmp1220);
	assign w_sys_tmp1233 = (r_run_copy0_j_73 + w_sys_intOne);
	assign w_sys_tmp1234 = (r_run_copy1_j_74 + w_sys_intOne);
	assign w_sys_tmp1235 = (r_run_copy2_j_75 + w_sys_intOne);
	assign w_sys_tmp1236 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp1357 = 32'sh00000070;
	assign w_sys_tmp1358 = ( !w_sys_tmp1359 );
	assign w_sys_tmp1359 = (w_sys_tmp1360 < r_run_j_36);
	assign w_sys_tmp1360 = 32'sh00000081;
	assign w_sys_tmp1363 = (w_sys_tmp1364 + r_run_k_35);
	assign w_sys_tmp1364 = (r_run_j_36 * w_sys_tmp1365);
	assign w_sys_tmp1365 = 32'sh00000081;
	assign w_sys_tmp1366 = w_fld_U_2_dataout_1;
	assign w_sys_tmp1367 = (w_sys_tmp1368 + r_run_k_35);
	assign w_sys_tmp1368 = (r_run_copy2_j_78 * w_sys_tmp1365);
	assign w_sys_tmp1371 = (w_sys_tmp1372 + r_run_k_35);
	assign w_sys_tmp1372 = (r_run_copy1_j_77 * w_sys_tmp1365);
	assign w_sys_tmp1374 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1375 = (w_sys_tmp1376 + r_run_k_35);
	assign w_sys_tmp1376 = (r_run_copy0_j_76 * w_sys_tmp1365);
	assign w_sys_tmp1378 = (r_run_copy0_j_76 + w_sys_intOne);
	assign w_sys_tmp1379 = (r_run_copy1_j_77 + w_sys_intOne);
	assign w_sys_tmp1380 = (r_run_copy2_j_78 + w_sys_intOne);
	assign w_sys_tmp1381 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp1502 = ( !w_sys_tmp1503 );
	assign w_sys_tmp1503 = (w_sys_tmp1504 < r_run_k_35);
	assign w_sys_tmp1504 = 32'sh00000021;
	assign w_sys_tmp1505 = (r_run_k_35 + w_sys_intOne);
	assign w_sys_tmp1506 = ( !w_sys_tmp1507 );
	assign w_sys_tmp1507 = (w_sys_tmp1508 < r_run_j_36);
	assign w_sys_tmp1508 = 32'sh00000011;
	assign w_sys_tmp1511 = (w_sys_tmp1512 + r_run_k_35);
	assign w_sys_tmp1512 = (r_run_j_36 * w_sys_tmp1513);
	assign w_sys_tmp1513 = 32'sh00000081;
	assign w_sys_tmp1514 = w_fld_U_2_dataout_1;
	assign w_sys_tmp1515 = (w_sys_tmp1516 + r_run_k_35);
	assign w_sys_tmp1516 = (r_run_copy2_j_81 * w_sys_tmp1513);
	assign w_sys_tmp1519 = (w_sys_tmp1520 + r_run_k_35);
	assign w_sys_tmp1520 = (r_run_copy1_j_80 * w_sys_tmp1513);
	assign w_sys_tmp1522 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1523 = (w_sys_tmp1524 + r_run_k_35);
	assign w_sys_tmp1524 = (r_run_copy0_j_79 * w_sys_tmp1513);
	assign w_sys_tmp1526 = (r_run_copy0_j_79 + w_sys_intOne);
	assign w_sys_tmp1527 = (r_run_copy1_j_80 + w_sys_intOne);
	assign w_sys_tmp1528 = (r_run_copy2_j_81 + w_sys_intOne);
	assign w_sys_tmp1529 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp1650 = 32'sh00000010;
	assign w_sys_tmp1651 = ( !w_sys_tmp1652 );
	assign w_sys_tmp1652 = (w_sys_tmp1653 < r_run_j_36);
	assign w_sys_tmp1653 = 32'sh00000021;
	assign w_sys_tmp1656 = (w_sys_tmp1657 + r_run_k_35);
	assign w_sys_tmp1657 = (r_run_j_36 * w_sys_tmp1658);
	assign w_sys_tmp1658 = 32'sh00000081;
	assign w_sys_tmp1659 = w_fld_U_2_dataout_1;
	assign w_sys_tmp1660 = (w_sys_tmp1661 + r_run_k_35);
	assign w_sys_tmp1661 = (r_run_copy2_j_84 * w_sys_tmp1658);
	assign w_sys_tmp1664 = (w_sys_tmp1665 + r_run_k_35);
	assign w_sys_tmp1665 = (r_run_copy1_j_83 * w_sys_tmp1658);
	assign w_sys_tmp1667 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1668 = (w_sys_tmp1669 + r_run_k_35);
	assign w_sys_tmp1669 = (r_run_copy0_j_82 * w_sys_tmp1658);
	assign w_sys_tmp1671 = (r_run_copy0_j_82 + w_sys_intOne);
	assign w_sys_tmp1672 = (r_run_copy1_j_83 + w_sys_intOne);
	assign w_sys_tmp1673 = (r_run_copy2_j_84 + w_sys_intOne);
	assign w_sys_tmp1674 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp1795 = 32'sh00000020;
	assign w_sys_tmp1796 = ( !w_sys_tmp1797 );
	assign w_sys_tmp1797 = (w_sys_tmp1798 < r_run_j_36);
	assign w_sys_tmp1798 = 32'sh00000031;
	assign w_sys_tmp1801 = (w_sys_tmp1802 + r_run_k_35);
	assign w_sys_tmp1802 = (r_run_j_36 * w_sys_tmp1803);
	assign w_sys_tmp1803 = 32'sh00000081;
	assign w_sys_tmp1804 = w_fld_U_2_dataout_1;
	assign w_sys_tmp1805 = (w_sys_tmp1806 + r_run_k_35);
	assign w_sys_tmp1806 = (r_run_copy2_j_87 * w_sys_tmp1803);
	assign w_sys_tmp1809 = (w_sys_tmp1810 + r_run_k_35);
	assign w_sys_tmp1810 = (r_run_copy1_j_86 * w_sys_tmp1803);
	assign w_sys_tmp1812 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1813 = (w_sys_tmp1814 + r_run_k_35);
	assign w_sys_tmp1814 = (r_run_copy0_j_85 * w_sys_tmp1803);
	assign w_sys_tmp1816 = (r_run_copy0_j_85 + w_sys_intOne);
	assign w_sys_tmp1817 = (r_run_copy1_j_86 + w_sys_intOne);
	assign w_sys_tmp1818 = (r_run_copy2_j_87 + w_sys_intOne);
	assign w_sys_tmp1819 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp1940 = 32'sh00000030;
	assign w_sys_tmp1941 = ( !w_sys_tmp1942 );
	assign w_sys_tmp1942 = (w_sys_tmp1943 < r_run_j_36);
	assign w_sys_tmp1943 = 32'sh00000041;
	assign w_sys_tmp1946 = (w_sys_tmp1947 + r_run_k_35);
	assign w_sys_tmp1947 = (r_run_j_36 * w_sys_tmp1948);
	assign w_sys_tmp1948 = 32'sh00000081;
	assign w_sys_tmp1949 = w_fld_U_2_dataout_1;
	assign w_sys_tmp1950 = (w_sys_tmp1951 + r_run_k_35);
	assign w_sys_tmp1951 = (r_run_copy2_j_90 * w_sys_tmp1948);
	assign w_sys_tmp1954 = (w_sys_tmp1955 + r_run_k_35);
	assign w_sys_tmp1955 = (r_run_copy1_j_89 * w_sys_tmp1948);
	assign w_sys_tmp1957 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1958 = (w_sys_tmp1959 + r_run_k_35);
	assign w_sys_tmp1959 = (r_run_copy0_j_88 * w_sys_tmp1948);
	assign w_sys_tmp1961 = (r_run_copy0_j_88 + w_sys_intOne);
	assign w_sys_tmp1962 = (r_run_copy1_j_89 + w_sys_intOne);
	assign w_sys_tmp1963 = (r_run_copy2_j_90 + w_sys_intOne);
	assign w_sys_tmp1964 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp2085 = 32'sh00000040;
	assign w_sys_tmp2086 = ( !w_sys_tmp2087 );
	assign w_sys_tmp2087 = (w_sys_tmp2088 < r_run_j_36);
	assign w_sys_tmp2088 = 32'sh00000051;
	assign w_sys_tmp2091 = (w_sys_tmp2092 + r_run_k_35);
	assign w_sys_tmp2092 = (r_run_j_36 * w_sys_tmp2093);
	assign w_sys_tmp2093 = 32'sh00000081;
	assign w_sys_tmp2094 = w_fld_U_2_dataout_1;
	assign w_sys_tmp2095 = (w_sys_tmp2096 + r_run_k_35);
	assign w_sys_tmp2096 = (r_run_copy2_j_93 * w_sys_tmp2093);
	assign w_sys_tmp2099 = (w_sys_tmp2100 + r_run_k_35);
	assign w_sys_tmp2100 = (r_run_copy1_j_92 * w_sys_tmp2093);
	assign w_sys_tmp2102 = w_fld_T_0_dataout_1;
	assign w_sys_tmp2103 = (w_sys_tmp2104 + r_run_k_35);
	assign w_sys_tmp2104 = (r_run_copy0_j_91 * w_sys_tmp2093);
	assign w_sys_tmp2106 = (r_run_copy0_j_91 + w_sys_intOne);
	assign w_sys_tmp2107 = (r_run_copy1_j_92 + w_sys_intOne);
	assign w_sys_tmp2108 = (r_run_copy2_j_93 + w_sys_intOne);
	assign w_sys_tmp2109 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp2230 = 32'sh00000050;
	assign w_sys_tmp2231 = ( !w_sys_tmp2232 );
	assign w_sys_tmp2232 = (w_sys_tmp2233 < r_run_j_36);
	assign w_sys_tmp2233 = 32'sh00000061;
	assign w_sys_tmp2236 = (w_sys_tmp2237 + r_run_k_35);
	assign w_sys_tmp2237 = (r_run_j_36 * w_sys_tmp2238);
	assign w_sys_tmp2238 = 32'sh00000081;
	assign w_sys_tmp2239 = w_fld_U_2_dataout_1;
	assign w_sys_tmp2240 = (w_sys_tmp2241 + r_run_k_35);
	assign w_sys_tmp2241 = (r_run_copy2_j_96 * w_sys_tmp2238);
	assign w_sys_tmp2244 = (w_sys_tmp2245 + r_run_k_35);
	assign w_sys_tmp2245 = (r_run_copy1_j_95 * w_sys_tmp2238);
	assign w_sys_tmp2247 = w_fld_T_0_dataout_1;
	assign w_sys_tmp2248 = (w_sys_tmp2249 + r_run_k_35);
	assign w_sys_tmp2249 = (r_run_copy0_j_94 * w_sys_tmp2238);
	assign w_sys_tmp2251 = (r_run_copy0_j_94 + w_sys_intOne);
	assign w_sys_tmp2252 = (r_run_copy1_j_95 + w_sys_intOne);
	assign w_sys_tmp2253 = (r_run_copy2_j_96 + w_sys_intOne);
	assign w_sys_tmp2254 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp2375 = 32'sh00000060;
	assign w_sys_tmp2376 = ( !w_sys_tmp2377 );
	assign w_sys_tmp2377 = (w_sys_tmp2378 < r_run_j_36);
	assign w_sys_tmp2378 = 32'sh00000071;
	assign w_sys_tmp2381 = (w_sys_tmp2382 + r_run_k_35);
	assign w_sys_tmp2382 = (r_run_j_36 * w_sys_tmp2383);
	assign w_sys_tmp2383 = 32'sh00000081;
	assign w_sys_tmp2384 = w_fld_U_2_dataout_1;
	assign w_sys_tmp2385 = (w_sys_tmp2386 + r_run_k_35);
	assign w_sys_tmp2386 = (r_run_copy2_j_99 * w_sys_tmp2383);
	assign w_sys_tmp2389 = (w_sys_tmp2390 + r_run_k_35);
	assign w_sys_tmp2390 = (r_run_copy1_j_98 * w_sys_tmp2383);
	assign w_sys_tmp2392 = w_fld_T_0_dataout_1;
	assign w_sys_tmp2393 = (w_sys_tmp2394 + r_run_k_35);
	assign w_sys_tmp2394 = (r_run_copy0_j_97 * w_sys_tmp2383);
	assign w_sys_tmp2396 = (r_run_copy0_j_97 + w_sys_intOne);
	assign w_sys_tmp2397 = (r_run_copy1_j_98 + w_sys_intOne);
	assign w_sys_tmp2398 = (r_run_copy2_j_99 + w_sys_intOne);
	assign w_sys_tmp2399 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp2520 = 32'sh00000070;
	assign w_sys_tmp2521 = ( !w_sys_tmp2522 );
	assign w_sys_tmp2522 = (w_sys_tmp2523 < r_run_j_36);
	assign w_sys_tmp2523 = 32'sh00000081;
	assign w_sys_tmp2526 = (w_sys_tmp2527 + r_run_k_35);
	assign w_sys_tmp2527 = (r_run_j_36 * w_sys_tmp2528);
	assign w_sys_tmp2528 = 32'sh00000081;
	assign w_sys_tmp2529 = w_fld_U_2_dataout_1;
	assign w_sys_tmp2530 = (w_sys_tmp2531 + r_run_k_35);
	assign w_sys_tmp2531 = (r_run_copy2_j_102 * w_sys_tmp2528);
	assign w_sys_tmp2534 = (w_sys_tmp2535 + r_run_k_35);
	assign w_sys_tmp2535 = (r_run_copy1_j_101 * w_sys_tmp2528);
	assign w_sys_tmp2537 = w_fld_T_0_dataout_1;
	assign w_sys_tmp2538 = (w_sys_tmp2539 + r_run_k_35);
	assign w_sys_tmp2539 = (r_run_copy0_j_100 * w_sys_tmp2528);
	assign w_sys_tmp2541 = (r_run_copy0_j_100 + w_sys_intOne);
	assign w_sys_tmp2542 = (r_run_copy1_j_101 + w_sys_intOne);
	assign w_sys_tmp2543 = (r_run_copy2_j_102 + w_sys_intOne);
	assign w_sys_tmp2544 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp2665 = ( !w_sys_tmp2666 );
	assign w_sys_tmp2666 = (w_sys_tmp2667 < r_run_k_35);
	assign w_sys_tmp2667 = 32'sh00000021;
	assign w_sys_tmp2668 = (r_run_k_35 + w_sys_intOne);
	assign w_sys_tmp2669 = ( !w_sys_tmp2670 );
	assign w_sys_tmp2670 = (w_sys_tmp2671 < r_run_j_36);
	assign w_sys_tmp2671 = 32'sh00000011;
	assign w_sys_tmp2674 = (w_sys_tmp2675 + r_run_k_35);
	assign w_sys_tmp2675 = (r_run_j_36 * w_sys_tmp2676);
	assign w_sys_tmp2676 = 32'sh00000081;
	assign w_sys_tmp2677 = w_fld_U_2_dataout_1;
	assign w_sys_tmp2678 = (w_sys_tmp2679 + r_run_k_35);
	assign w_sys_tmp2679 = (r_run_copy2_j_105 * w_sys_tmp2676);
	assign w_sys_tmp2682 = (w_sys_tmp2683 + r_run_k_35);
	assign w_sys_tmp2683 = (r_run_copy1_j_104 * w_sys_tmp2676);
	assign w_sys_tmp2685 = w_fld_T_0_dataout_1;
	assign w_sys_tmp2686 = (w_sys_tmp2687 + r_run_k_35);
	assign w_sys_tmp2687 = (r_run_copy0_j_103 * w_sys_tmp2676);
	assign w_sys_tmp2689 = (r_run_copy0_j_103 + w_sys_intOne);
	assign w_sys_tmp2690 = (r_run_copy1_j_104 + w_sys_intOne);
	assign w_sys_tmp2691 = (r_run_copy2_j_105 + w_sys_intOne);
	assign w_sys_tmp2692 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp2813 = 32'sh00000010;
	assign w_sys_tmp2814 = ( !w_sys_tmp2815 );
	assign w_sys_tmp2815 = (w_sys_tmp2816 < r_run_j_36);
	assign w_sys_tmp2816 = 32'sh00000021;
	assign w_sys_tmp2819 = (w_sys_tmp2820 + r_run_k_35);
	assign w_sys_tmp2820 = (r_run_j_36 * w_sys_tmp2821);
	assign w_sys_tmp2821 = 32'sh00000081;
	assign w_sys_tmp2822 = w_fld_U_2_dataout_1;
	assign w_sys_tmp2823 = (w_sys_tmp2824 + r_run_k_35);
	assign w_sys_tmp2824 = (r_run_copy2_j_108 * w_sys_tmp2821);
	assign w_sys_tmp2827 = (w_sys_tmp2828 + r_run_k_35);
	assign w_sys_tmp2828 = (r_run_copy1_j_107 * w_sys_tmp2821);
	assign w_sys_tmp2830 = w_fld_T_0_dataout_1;
	assign w_sys_tmp2831 = (w_sys_tmp2832 + r_run_k_35);
	assign w_sys_tmp2832 = (r_run_copy0_j_106 * w_sys_tmp2821);
	assign w_sys_tmp2834 = (r_run_copy0_j_106 + w_sys_intOne);
	assign w_sys_tmp2835 = (r_run_copy1_j_107 + w_sys_intOne);
	assign w_sys_tmp2836 = (r_run_copy2_j_108 + w_sys_intOne);
	assign w_sys_tmp2837 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp2958 = 32'sh00000020;
	assign w_sys_tmp2959 = ( !w_sys_tmp2960 );
	assign w_sys_tmp2960 = (w_sys_tmp2961 < r_run_j_36);
	assign w_sys_tmp2961 = 32'sh00000031;
	assign w_sys_tmp2964 = (w_sys_tmp2965 + r_run_k_35);
	assign w_sys_tmp2965 = (r_run_j_36 * w_sys_tmp2966);
	assign w_sys_tmp2966 = 32'sh00000081;
	assign w_sys_tmp2967 = w_fld_U_2_dataout_1;
	assign w_sys_tmp2968 = (w_sys_tmp2969 + r_run_k_35);
	assign w_sys_tmp2969 = (r_run_copy2_j_111 * w_sys_tmp2966);
	assign w_sys_tmp2972 = (w_sys_tmp2973 + r_run_k_35);
	assign w_sys_tmp2973 = (r_run_copy1_j_110 * w_sys_tmp2966);
	assign w_sys_tmp2975 = w_fld_T_0_dataout_1;
	assign w_sys_tmp2976 = (w_sys_tmp2977 + r_run_k_35);
	assign w_sys_tmp2977 = (r_run_copy0_j_109 * w_sys_tmp2966);
	assign w_sys_tmp2979 = (r_run_copy0_j_109 + w_sys_intOne);
	assign w_sys_tmp2980 = (r_run_copy1_j_110 + w_sys_intOne);
	assign w_sys_tmp2981 = (r_run_copy2_j_111 + w_sys_intOne);
	assign w_sys_tmp2982 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp3103 = 32'sh00000030;
	assign w_sys_tmp3104 = ( !w_sys_tmp3105 );
	assign w_sys_tmp3105 = (w_sys_tmp3106 < r_run_j_36);
	assign w_sys_tmp3106 = 32'sh00000041;
	assign w_sys_tmp3109 = (w_sys_tmp3110 + r_run_k_35);
	assign w_sys_tmp3110 = (r_run_j_36 * w_sys_tmp3111);
	assign w_sys_tmp3111 = 32'sh00000081;
	assign w_sys_tmp3112 = w_fld_U_2_dataout_1;
	assign w_sys_tmp3113 = (w_sys_tmp3114 + r_run_k_35);
	assign w_sys_tmp3114 = (r_run_copy2_j_114 * w_sys_tmp3111);
	assign w_sys_tmp3117 = (w_sys_tmp3118 + r_run_k_35);
	assign w_sys_tmp3118 = (r_run_copy1_j_113 * w_sys_tmp3111);
	assign w_sys_tmp3120 = w_fld_T_0_dataout_1;
	assign w_sys_tmp3121 = (w_sys_tmp3122 + r_run_k_35);
	assign w_sys_tmp3122 = (r_run_copy0_j_112 * w_sys_tmp3111);
	assign w_sys_tmp3124 = (r_run_copy0_j_112 + w_sys_intOne);
	assign w_sys_tmp3125 = (r_run_copy1_j_113 + w_sys_intOne);
	assign w_sys_tmp3126 = (r_run_copy2_j_114 + w_sys_intOne);
	assign w_sys_tmp3127 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp3248 = 32'sh00000040;
	assign w_sys_tmp3249 = ( !w_sys_tmp3250 );
	assign w_sys_tmp3250 = (w_sys_tmp3251 < r_run_j_36);
	assign w_sys_tmp3251 = 32'sh00000051;
	assign w_sys_tmp3254 = (w_sys_tmp3255 + r_run_k_35);
	assign w_sys_tmp3255 = (r_run_j_36 * w_sys_tmp3256);
	assign w_sys_tmp3256 = 32'sh00000081;
	assign w_sys_tmp3257 = w_fld_U_2_dataout_1;
	assign w_sys_tmp3258 = (w_sys_tmp3259 + r_run_k_35);
	assign w_sys_tmp3259 = (r_run_copy2_j_117 * w_sys_tmp3256);
	assign w_sys_tmp3262 = (w_sys_tmp3263 + r_run_k_35);
	assign w_sys_tmp3263 = (r_run_copy1_j_116 * w_sys_tmp3256);
	assign w_sys_tmp3265 = w_fld_T_0_dataout_1;
	assign w_sys_tmp3266 = (w_sys_tmp3267 + r_run_k_35);
	assign w_sys_tmp3267 = (r_run_copy0_j_115 * w_sys_tmp3256);
	assign w_sys_tmp3269 = (r_run_copy0_j_115 + w_sys_intOne);
	assign w_sys_tmp3270 = (r_run_copy1_j_116 + w_sys_intOne);
	assign w_sys_tmp3271 = (r_run_copy2_j_117 + w_sys_intOne);
	assign w_sys_tmp3272 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp3393 = 32'sh00000050;
	assign w_sys_tmp3394 = ( !w_sys_tmp3395 );
	assign w_sys_tmp3395 = (w_sys_tmp3396 < r_run_j_36);
	assign w_sys_tmp3396 = 32'sh00000061;
	assign w_sys_tmp3399 = (w_sys_tmp3400 + r_run_k_35);
	assign w_sys_tmp3400 = (r_run_j_36 * w_sys_tmp3401);
	assign w_sys_tmp3401 = 32'sh00000081;
	assign w_sys_tmp3402 = w_fld_U_2_dataout_1;
	assign w_sys_tmp3403 = (w_sys_tmp3404 + r_run_k_35);
	assign w_sys_tmp3404 = (r_run_copy2_j_120 * w_sys_tmp3401);
	assign w_sys_tmp3407 = (w_sys_tmp3408 + r_run_k_35);
	assign w_sys_tmp3408 = (r_run_copy1_j_119 * w_sys_tmp3401);
	assign w_sys_tmp3410 = w_fld_T_0_dataout_1;
	assign w_sys_tmp3411 = (w_sys_tmp3412 + r_run_k_35);
	assign w_sys_tmp3412 = (r_run_copy0_j_118 * w_sys_tmp3401);
	assign w_sys_tmp3414 = (r_run_copy0_j_118 + w_sys_intOne);
	assign w_sys_tmp3415 = (r_run_copy1_j_119 + w_sys_intOne);
	assign w_sys_tmp3416 = (r_run_copy2_j_120 + w_sys_intOne);
	assign w_sys_tmp3417 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp3538 = 32'sh00000060;
	assign w_sys_tmp3539 = ( !w_sys_tmp3540 );
	assign w_sys_tmp3540 = (w_sys_tmp3541 < r_run_j_36);
	assign w_sys_tmp3541 = 32'sh00000071;
	assign w_sys_tmp3544 = (w_sys_tmp3545 + r_run_k_35);
	assign w_sys_tmp3545 = (r_run_j_36 * w_sys_tmp3546);
	assign w_sys_tmp3546 = 32'sh00000081;
	assign w_sys_tmp3547 = w_fld_U_2_dataout_1;
	assign w_sys_tmp3548 = (w_sys_tmp3549 + r_run_k_35);
	assign w_sys_tmp3549 = (r_run_copy2_j_123 * w_sys_tmp3546);
	assign w_sys_tmp3552 = (w_sys_tmp3553 + r_run_k_35);
	assign w_sys_tmp3553 = (r_run_copy1_j_122 * w_sys_tmp3546);
	assign w_sys_tmp3555 = w_fld_T_0_dataout_1;
	assign w_sys_tmp3556 = (w_sys_tmp3557 + r_run_k_35);
	assign w_sys_tmp3557 = (r_run_copy0_j_121 * w_sys_tmp3546);
	assign w_sys_tmp3559 = (r_run_copy0_j_121 + w_sys_intOne);
	assign w_sys_tmp3560 = (r_run_copy1_j_122 + w_sys_intOne);
	assign w_sys_tmp3561 = (r_run_copy2_j_123 + w_sys_intOne);
	assign w_sys_tmp3562 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp3683 = 32'sh00000070;
	assign w_sys_tmp3684 = ( !w_sys_tmp3685 );
	assign w_sys_tmp3685 = (w_sys_tmp3686 < r_run_j_36);
	assign w_sys_tmp3686 = 32'sh00000081;
	assign w_sys_tmp3689 = (w_sys_tmp3690 + r_run_k_35);
	assign w_sys_tmp3690 = (r_run_j_36 * w_sys_tmp3691);
	assign w_sys_tmp3691 = 32'sh00000081;
	assign w_sys_tmp3692 = w_fld_U_2_dataout_1;
	assign w_sys_tmp3693 = (w_sys_tmp3694 + r_run_k_35);
	assign w_sys_tmp3694 = (r_run_copy2_j_126 * w_sys_tmp3691);
	assign w_sys_tmp3697 = (w_sys_tmp3698 + r_run_k_35);
	assign w_sys_tmp3698 = (r_run_copy1_j_125 * w_sys_tmp3691);
	assign w_sys_tmp3700 = w_fld_T_0_dataout_1;
	assign w_sys_tmp3701 = (w_sys_tmp3702 + r_run_k_35);
	assign w_sys_tmp3702 = (r_run_copy0_j_124 * w_sys_tmp3691);
	assign w_sys_tmp3704 = (r_run_copy0_j_124 + w_sys_intOne);
	assign w_sys_tmp3705 = (r_run_copy1_j_125 + w_sys_intOne);
	assign w_sys_tmp3706 = (r_run_copy2_j_126 + w_sys_intOne);
	assign w_sys_tmp3707 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp3828 = ( !w_sys_tmp3829 );
	assign w_sys_tmp3829 = (w_sys_tmp3830 < r_run_k_35);
	assign w_sys_tmp3830 = 32'sh00000021;
	assign w_sys_tmp3831 = (r_run_k_35 + w_sys_intOne);
	assign w_sys_tmp3832 = ( !w_sys_tmp3833 );
	assign w_sys_tmp3833 = (w_sys_tmp3834 < r_run_j_36);
	assign w_sys_tmp3834 = 32'sh00000011;
	assign w_sys_tmp3837 = (w_sys_tmp3838 + r_run_k_35);
	assign w_sys_tmp3838 = (r_run_j_36 * w_sys_tmp3839);
	assign w_sys_tmp3839 = 32'sh00000081;
	assign w_sys_tmp3840 = w_fld_U_2_dataout_1;
	assign w_sys_tmp3841 = (w_sys_tmp3842 + r_run_k_35);
	assign w_sys_tmp3842 = (r_run_copy2_j_129 * w_sys_tmp3839);
	assign w_sys_tmp3845 = (w_sys_tmp3846 + r_run_k_35);
	assign w_sys_tmp3846 = (r_run_copy1_j_128 * w_sys_tmp3839);
	assign w_sys_tmp3848 = w_fld_T_0_dataout_1;
	assign w_sys_tmp3849 = (w_sys_tmp3850 + r_run_k_35);
	assign w_sys_tmp3850 = (r_run_copy0_j_127 * w_sys_tmp3839);
	assign w_sys_tmp3852 = (r_run_copy0_j_127 + w_sys_intOne);
	assign w_sys_tmp3853 = (r_run_copy1_j_128 + w_sys_intOne);
	assign w_sys_tmp3854 = (r_run_copy2_j_129 + w_sys_intOne);
	assign w_sys_tmp3855 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp3976 = 32'sh00000010;
	assign w_sys_tmp3977 = ( !w_sys_tmp3978 );
	assign w_sys_tmp3978 = (w_sys_tmp3979 < r_run_j_36);
	assign w_sys_tmp3979 = 32'sh00000021;
	assign w_sys_tmp3982 = (w_sys_tmp3983 + r_run_k_35);
	assign w_sys_tmp3983 = (r_run_j_36 * w_sys_tmp3984);
	assign w_sys_tmp3984 = 32'sh00000081;
	assign w_sys_tmp3985 = w_fld_U_2_dataout_1;
	assign w_sys_tmp3986 = (w_sys_tmp3987 + r_run_k_35);
	assign w_sys_tmp3987 = (r_run_copy2_j_132 * w_sys_tmp3984);
	assign w_sys_tmp3990 = (w_sys_tmp3991 + r_run_k_35);
	assign w_sys_tmp3991 = (r_run_copy1_j_131 * w_sys_tmp3984);
	assign w_sys_tmp3993 = w_fld_T_0_dataout_1;
	assign w_sys_tmp3994 = (w_sys_tmp3995 + r_run_k_35);
	assign w_sys_tmp3995 = (r_run_copy0_j_130 * w_sys_tmp3984);
	assign w_sys_tmp3997 = (r_run_copy0_j_130 + w_sys_intOne);
	assign w_sys_tmp3998 = (r_run_copy1_j_131 + w_sys_intOne);
	assign w_sys_tmp3999 = (r_run_copy2_j_132 + w_sys_intOne);
	assign w_sys_tmp4000 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp4121 = 32'sh00000020;
	assign w_sys_tmp4122 = ( !w_sys_tmp4123 );
	assign w_sys_tmp4123 = (w_sys_tmp4124 < r_run_j_36);
	assign w_sys_tmp4124 = 32'sh00000031;
	assign w_sys_tmp4127 = (w_sys_tmp4128 + r_run_k_35);
	assign w_sys_tmp4128 = (r_run_j_36 * w_sys_tmp4129);
	assign w_sys_tmp4129 = 32'sh00000081;
	assign w_sys_tmp4130 = w_fld_U_2_dataout_1;
	assign w_sys_tmp4131 = (w_sys_tmp4132 + r_run_k_35);
	assign w_sys_tmp4132 = (r_run_copy2_j_135 * w_sys_tmp4129);
	assign w_sys_tmp4135 = (w_sys_tmp4136 + r_run_k_35);
	assign w_sys_tmp4136 = (r_run_copy1_j_134 * w_sys_tmp4129);
	assign w_sys_tmp4138 = w_fld_T_0_dataout_1;
	assign w_sys_tmp4139 = (w_sys_tmp4140 + r_run_k_35);
	assign w_sys_tmp4140 = (r_run_copy0_j_133 * w_sys_tmp4129);
	assign w_sys_tmp4142 = (r_run_copy0_j_133 + w_sys_intOne);
	assign w_sys_tmp4143 = (r_run_copy1_j_134 + w_sys_intOne);
	assign w_sys_tmp4144 = (r_run_copy2_j_135 + w_sys_intOne);
	assign w_sys_tmp4145 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp4266 = 32'sh00000030;
	assign w_sys_tmp4267 = ( !w_sys_tmp4268 );
	assign w_sys_tmp4268 = (w_sys_tmp4269 < r_run_j_36);
	assign w_sys_tmp4269 = 32'sh00000041;
	assign w_sys_tmp4272 = (w_sys_tmp4273 + r_run_k_35);
	assign w_sys_tmp4273 = (r_run_j_36 * w_sys_tmp4274);
	assign w_sys_tmp4274 = 32'sh00000081;
	assign w_sys_tmp4275 = w_fld_U_2_dataout_1;
	assign w_sys_tmp4276 = (w_sys_tmp4277 + r_run_k_35);
	assign w_sys_tmp4277 = (r_run_copy2_j_138 * w_sys_tmp4274);
	assign w_sys_tmp4280 = (w_sys_tmp4281 + r_run_k_35);
	assign w_sys_tmp4281 = (r_run_copy1_j_137 * w_sys_tmp4274);
	assign w_sys_tmp4283 = w_fld_T_0_dataout_1;
	assign w_sys_tmp4284 = (w_sys_tmp4285 + r_run_k_35);
	assign w_sys_tmp4285 = (r_run_copy0_j_136 * w_sys_tmp4274);
	assign w_sys_tmp4287 = (r_run_copy0_j_136 + w_sys_intOne);
	assign w_sys_tmp4288 = (r_run_copy1_j_137 + w_sys_intOne);
	assign w_sys_tmp4289 = (r_run_copy2_j_138 + w_sys_intOne);
	assign w_sys_tmp4290 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp4411 = 32'sh00000040;
	assign w_sys_tmp4412 = ( !w_sys_tmp4413 );
	assign w_sys_tmp4413 = (w_sys_tmp4414 < r_run_j_36);
	assign w_sys_tmp4414 = 32'sh00000051;
	assign w_sys_tmp4417 = (w_sys_tmp4418 + r_run_k_35);
	assign w_sys_tmp4418 = (r_run_j_36 * w_sys_tmp4419);
	assign w_sys_tmp4419 = 32'sh00000081;
	assign w_sys_tmp4420 = w_fld_U_2_dataout_1;
	assign w_sys_tmp4421 = (w_sys_tmp4422 + r_run_k_35);
	assign w_sys_tmp4422 = (r_run_copy2_j_141 * w_sys_tmp4419);
	assign w_sys_tmp4425 = (w_sys_tmp4426 + r_run_k_35);
	assign w_sys_tmp4426 = (r_run_copy1_j_140 * w_sys_tmp4419);
	assign w_sys_tmp4428 = w_fld_T_0_dataout_1;
	assign w_sys_tmp4429 = (w_sys_tmp4430 + r_run_k_35);
	assign w_sys_tmp4430 = (r_run_copy0_j_139 * w_sys_tmp4419);
	assign w_sys_tmp4432 = (r_run_copy0_j_139 + w_sys_intOne);
	assign w_sys_tmp4433 = (r_run_copy1_j_140 + w_sys_intOne);
	assign w_sys_tmp4434 = (r_run_copy2_j_141 + w_sys_intOne);
	assign w_sys_tmp4435 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp4556 = 32'sh00000050;
	assign w_sys_tmp4557 = ( !w_sys_tmp4558 );
	assign w_sys_tmp4558 = (w_sys_tmp4559 < r_run_j_36);
	assign w_sys_tmp4559 = 32'sh00000061;
	assign w_sys_tmp4562 = (w_sys_tmp4563 + r_run_k_35);
	assign w_sys_tmp4563 = (r_run_j_36 * w_sys_tmp4564);
	assign w_sys_tmp4564 = 32'sh00000081;
	assign w_sys_tmp4565 = w_fld_U_2_dataout_1;
	assign w_sys_tmp4566 = (w_sys_tmp4567 + r_run_k_35);
	assign w_sys_tmp4567 = (r_run_copy2_j_144 * w_sys_tmp4564);
	assign w_sys_tmp4570 = (w_sys_tmp4571 + r_run_k_35);
	assign w_sys_tmp4571 = (r_run_copy1_j_143 * w_sys_tmp4564);
	assign w_sys_tmp4573 = w_fld_T_0_dataout_1;
	assign w_sys_tmp4574 = (w_sys_tmp4575 + r_run_k_35);
	assign w_sys_tmp4575 = (r_run_copy0_j_142 * w_sys_tmp4564);
	assign w_sys_tmp4577 = (r_run_copy0_j_142 + w_sys_intOne);
	assign w_sys_tmp4578 = (r_run_copy1_j_143 + w_sys_intOne);
	assign w_sys_tmp4579 = (r_run_copy2_j_144 + w_sys_intOne);
	assign w_sys_tmp4580 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp4701 = 32'sh00000060;
	assign w_sys_tmp4702 = ( !w_sys_tmp4703 );
	assign w_sys_tmp4703 = (w_sys_tmp4704 < r_run_j_36);
	assign w_sys_tmp4704 = 32'sh00000071;
	assign w_sys_tmp4707 = (w_sys_tmp4708 + r_run_k_35);
	assign w_sys_tmp4708 = (r_run_j_36 * w_sys_tmp4709);
	assign w_sys_tmp4709 = 32'sh00000081;
	assign w_sys_tmp4710 = w_fld_U_2_dataout_1;
	assign w_sys_tmp4711 = (w_sys_tmp4712 + r_run_k_35);
	assign w_sys_tmp4712 = (r_run_copy2_j_147 * w_sys_tmp4709);
	assign w_sys_tmp4715 = (w_sys_tmp4716 + r_run_k_35);
	assign w_sys_tmp4716 = (r_run_copy1_j_146 * w_sys_tmp4709);
	assign w_sys_tmp4718 = w_fld_T_0_dataout_1;
	assign w_sys_tmp4719 = (w_sys_tmp4720 + r_run_k_35);
	assign w_sys_tmp4720 = (r_run_copy0_j_145 * w_sys_tmp4709);
	assign w_sys_tmp4722 = (r_run_copy0_j_145 + w_sys_intOne);
	assign w_sys_tmp4723 = (r_run_copy1_j_146 + w_sys_intOne);
	assign w_sys_tmp4724 = (r_run_copy2_j_147 + w_sys_intOne);
	assign w_sys_tmp4725 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp4846 = 32'sh00000070;
	assign w_sys_tmp4847 = ( !w_sys_tmp4848 );
	assign w_sys_tmp4848 = (w_sys_tmp4849 < r_run_j_36);
	assign w_sys_tmp4849 = 32'sh00000081;
	assign w_sys_tmp4852 = (w_sys_tmp4853 + r_run_k_35);
	assign w_sys_tmp4853 = (r_run_j_36 * w_sys_tmp4854);
	assign w_sys_tmp4854 = 32'sh00000081;
	assign w_sys_tmp4855 = w_fld_U_2_dataout_1;
	assign w_sys_tmp4856 = (w_sys_tmp4857 + r_run_k_35);
	assign w_sys_tmp4857 = (r_run_copy2_j_150 * w_sys_tmp4854);
	assign w_sys_tmp4860 = (w_sys_tmp4861 + r_run_k_35);
	assign w_sys_tmp4861 = (r_run_copy1_j_149 * w_sys_tmp4854);
	assign w_sys_tmp4863 = w_fld_T_0_dataout_1;
	assign w_sys_tmp4864 = (w_sys_tmp4865 + r_run_k_35);
	assign w_sys_tmp4865 = (r_run_copy0_j_148 * w_sys_tmp4854);
	assign w_sys_tmp4867 = (r_run_copy0_j_148 + w_sys_intOne);
	assign w_sys_tmp4868 = (r_run_copy1_j_149 + w_sys_intOne);
	assign w_sys_tmp4869 = (r_run_copy2_j_150 + w_sys_intOne);
	assign w_sys_tmp4870 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp4991 = ( !w_sys_tmp4992 );
	assign w_sys_tmp4992 = (r_run_nlast_50 < r_run_n_37);
	assign w_sys_tmp4993 = (r_run_n_37 + w_sys_intOne);
	assign w_sys_tmp4994 = 32'sh00000002;
	assign w_sys_tmp4995 = ( !w_sys_tmp4996 );
	assign w_sys_tmp4996 = (w_sys_tmp4997 < r_run_k_35);
	assign w_sys_tmp4997 = 32'sh00000020;
	assign w_sys_tmp5000 = (w_sys_tmp5001 + r_run_k_35);
	assign w_sys_tmp5001 = 32'sh00000891;
	assign w_sys_tmp5002 = w_sub01_result_dataout;
	assign w_sys_tmp5003 = (w_sys_tmp5004 + r_run_k_35);
	assign w_sys_tmp5004 = 32'sh00000102;
	assign w_sys_tmp5006 = (w_sys_tmp5007 + r_run_k_35);
	assign w_sys_tmp5007 = 32'sh00000081;
	assign w_sys_tmp5008 = w_sub00_result_dataout;
	assign w_sys_tmp5009 = (w_sys_tmp5010 + r_run_k_35);
	assign w_sys_tmp5010 = 32'sh00000810;
	assign w_sys_tmp5012 = (w_sys_tmp5013 + r_run_k_35);
	assign w_sys_tmp5013 = 32'sh00000912;
	assign w_sys_tmp5030 = w_sub02_result_dataout;
	assign w_sys_tmp5041 = w_sub03_result_dataout;
	assign w_sys_tmp5052 = w_sub04_result_dataout;
	assign w_sys_tmp5063 = w_sub05_result_dataout;
	assign w_sys_tmp5074 = w_sub06_result_dataout;
	assign w_sys_tmp5077 = (r_run_k_35 + w_sys_intOne);
	assign w_sys_tmp5078 = 32'sh00000020;
	assign w_sys_tmp5079 = ( !w_sys_tmp5080 );
	assign w_sys_tmp5080 = (w_sys_tmp5081 < r_run_k_35);
	assign w_sys_tmp5081 = 32'sh00000041;
	assign w_sys_tmp5084 = (w_sys_tmp5085 + r_run_k_35);
	assign w_sys_tmp5085 = 32'sh00000891;
	assign w_sys_tmp5086 = w_sub09_result_dataout;
	assign w_sys_tmp5087 = (w_sys_tmp5088 + r_run_k_35);
	assign w_sys_tmp5088 = 32'sh00000102;
	assign w_sys_tmp5090 = (w_sys_tmp5091 + r_run_k_35);
	assign w_sys_tmp5091 = 32'sh00000081;
	assign w_sys_tmp5092 = w_sub08_result_dataout;
	assign w_sys_tmp5093 = (w_sys_tmp5094 + r_run_k_35);
	assign w_sys_tmp5094 = 32'sh00000810;
	assign w_sys_tmp5096 = (w_sys_tmp5097 + r_run_k_35);
	assign w_sys_tmp5097 = 32'sh00000912;
	assign w_sys_tmp5114 = w_sub10_result_dataout;
	assign w_sys_tmp5125 = w_sub11_result_dataout;
	assign w_sys_tmp5136 = w_sub12_result_dataout;
	assign w_sys_tmp5147 = w_sub13_result_dataout;
	assign w_sys_tmp5158 = w_sub14_result_dataout;
	assign w_sys_tmp5161 = (r_run_k_35 + w_sys_intOne);
	assign w_sys_tmp5162 = 32'sh00000040;
	assign w_sys_tmp5163 = ( !w_sys_tmp5164 );
	assign w_sys_tmp5164 = (w_sys_tmp5165 < r_run_k_35);
	assign w_sys_tmp5165 = 32'sh00000061;
	assign w_sys_tmp5168 = (w_sys_tmp5169 + r_run_k_35);
	assign w_sys_tmp5169 = 32'sh00000891;
	assign w_sys_tmp5170 = w_sub17_result_dataout;
	assign w_sys_tmp5171 = (w_sys_tmp5172 + r_run_k_35);
	assign w_sys_tmp5172 = 32'sh00000102;
	assign w_sys_tmp5174 = (w_sys_tmp5175 + r_run_k_35);
	assign w_sys_tmp5175 = 32'sh00000081;
	assign w_sys_tmp5176 = w_sub16_result_dataout;
	assign w_sys_tmp5177 = (w_sys_tmp5178 + r_run_k_35);
	assign w_sys_tmp5178 = 32'sh00000810;
	assign w_sys_tmp5180 = (w_sys_tmp5181 + r_run_k_35);
	assign w_sys_tmp5181 = 32'sh00000912;
	assign w_sys_tmp5198 = w_sub18_result_dataout;
	assign w_sys_tmp5209 = w_sub19_result_dataout;
	assign w_sys_tmp5220 = w_sub20_result_dataout;
	assign w_sys_tmp5231 = w_sub21_result_dataout;
	assign w_sys_tmp5242 = w_sub22_result_dataout;
	assign w_sys_tmp5245 = (r_run_k_35 + w_sys_intOne);
	assign w_sys_tmp5246 = 32'sh00000060;
	assign w_sys_tmp5247 = ( !w_sys_tmp5248 );
	assign w_sys_tmp5248 = (w_sys_tmp5249 < r_run_k_35);
	assign w_sys_tmp5249 = 32'sh00000081;
	assign w_sys_tmp5252 = (w_sys_tmp5253 + r_run_k_35);
	assign w_sys_tmp5253 = 32'sh00000891;
	assign w_sys_tmp5254 = w_sub25_result_dataout;
	assign w_sys_tmp5255 = (w_sys_tmp5256 + r_run_k_35);
	assign w_sys_tmp5256 = 32'sh00000102;
	assign w_sys_tmp5258 = (w_sys_tmp5259 + r_run_k_35);
	assign w_sys_tmp5259 = 32'sh00000081;
	assign w_sys_tmp5260 = w_sub24_result_dataout;
	assign w_sys_tmp5261 = (w_sys_tmp5262 + r_run_k_35);
	assign w_sys_tmp5262 = 32'sh00000810;
	assign w_sys_tmp5264 = (w_sys_tmp5265 + r_run_k_35);
	assign w_sys_tmp5265 = 32'sh00000912;
	assign w_sys_tmp5282 = w_sub26_result_dataout;
	assign w_sys_tmp5293 = w_sub27_result_dataout;
	assign w_sys_tmp5304 = w_sub28_result_dataout;
	assign w_sys_tmp5315 = w_sub29_result_dataout;
	assign w_sys_tmp5326 = w_sub30_result_dataout;
	assign w_sys_tmp5329 = (r_run_k_35 + w_sys_intOne);
	assign w_sys_tmp5330 = ( !w_sys_tmp5331 );
	assign w_sys_tmp5331 = (w_sys_tmp5332 < r_run_j_36);
	assign w_sys_tmp5332 = 32'sh00000011;
	assign w_sys_tmp5335 = (w_sys_tmp5336 + w_sys_tmp5338);
	assign w_sys_tmp5336 = (r_run_j_36 * w_sys_tmp5337);
	assign w_sys_tmp5337 = 32'sh00000081;
	assign w_sys_tmp5338 = 32'sh00000021;
	assign w_sys_tmp5339 = w_sub08_result_dataout;
	assign w_sys_tmp5340 = (w_sys_tmp5341 + w_sys_tmp5338);
	assign w_sys_tmp5341 = (r_run_copy10_j_161 * w_sys_tmp5337);
	assign w_sys_tmp5345 = (w_sys_tmp5346 + w_sys_tmp5348);
	assign w_sys_tmp5346 = (r_run_copy9_j_160 * w_sys_tmp5337);
	assign w_sys_tmp5348 = 32'sh00000020;
	assign w_sys_tmp5349 = w_sub00_result_dataout;
	assign w_sys_tmp5350 = (w_sys_tmp5351 + w_sys_tmp5348);
	assign w_sys_tmp5351 = (r_run_copy8_j_159 * w_sys_tmp5337);
	assign w_sys_tmp5355 = (w_sys_tmp5356 + w_sys_tmp5358);
	assign w_sys_tmp5356 = (r_run_copy7_j_158 * w_sys_tmp5337);
	assign w_sys_tmp5358 = 32'sh00000041;
	assign w_sys_tmp5359 = (w_sys_tmp5360 + w_sys_tmp5358);
	assign w_sys_tmp5360 = (r_run_copy6_j_157 * w_sys_tmp5337);
	assign w_sys_tmp5364 = (w_sys_tmp5365 + w_sys_tmp5367);
	assign w_sys_tmp5365 = (r_run_copy5_j_156 * w_sys_tmp5337);
	assign w_sys_tmp5367 = 32'sh00000040;
	assign w_sys_tmp5369 = (w_sys_tmp5370 + w_sys_tmp5367);
	assign w_sys_tmp5370 = (r_run_copy4_j_155 * w_sys_tmp5337);
	assign w_sys_tmp5374 = (w_sys_tmp5375 + w_sys_tmp5377);
	assign w_sys_tmp5375 = (r_run_copy3_j_154 * w_sys_tmp5337);
	assign w_sys_tmp5377 = 32'sh00000061;
	assign w_sys_tmp5378 = (w_sys_tmp5379 + w_sys_tmp5377);
	assign w_sys_tmp5379 = (r_run_copy2_j_153 * w_sys_tmp5337);
	assign w_sys_tmp5383 = (w_sys_tmp5384 + w_sys_tmp5386);
	assign w_sys_tmp5384 = (r_run_copy1_j_152 * w_sys_tmp5337);
	assign w_sys_tmp5386 = 32'sh00000060;
	assign w_sys_tmp5387 = w_sub16_result_dataout;
	assign w_sys_tmp5388 = (w_sys_tmp5389 + w_sys_tmp5386);
	assign w_sys_tmp5389 = (r_run_copy0_j_151 * w_sys_tmp5337);
	assign w_sys_tmp5392 = (r_run_copy0_j_151 + w_sys_intOne);
	assign w_sys_tmp5393 = (r_run_copy1_j_152 + w_sys_intOne);
	assign w_sys_tmp5394 = (r_run_copy2_j_153 + w_sys_intOne);
	assign w_sys_tmp5395 = (r_run_copy3_j_154 + w_sys_intOne);
	assign w_sys_tmp5396 = (r_run_copy4_j_155 + w_sys_intOne);
	assign w_sys_tmp5397 = (r_run_copy5_j_156 + w_sys_intOne);
	assign w_sys_tmp5398 = (r_run_copy6_j_157 + w_sys_intOne);
	assign w_sys_tmp5399 = (r_run_copy7_j_158 + w_sys_intOne);
	assign w_sys_tmp5400 = (r_run_copy8_j_159 + w_sys_intOne);
	assign w_sys_tmp5401 = (r_run_copy9_j_160 + w_sys_intOne);
	assign w_sys_tmp5402 = (r_run_copy10_j_161 + w_sys_intOne);
	assign w_sys_tmp5403 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp5830 = 32'sh00000010;
	assign w_sys_tmp5831 = ( !w_sys_tmp5832 );
	assign w_sys_tmp5832 = (w_sys_tmp5833 < r_run_j_36);
	assign w_sys_tmp5833 = 32'sh00000021;
	assign w_sys_tmp5836 = (w_sys_tmp5837 + w_sys_tmp5839);
	assign w_sys_tmp5837 = (r_run_j_36 * w_sys_tmp5838);
	assign w_sys_tmp5838 = 32'sh00000081;
	assign w_sys_tmp5839 = 32'sh00000021;
	assign w_sys_tmp5840 = w_sub09_result_dataout;
	assign w_sys_tmp5841 = (w_sys_tmp5842 + w_sys_tmp5839);
	assign w_sys_tmp5842 = (r_run_copy10_j_172 * w_sys_tmp5838);
	assign w_sys_tmp5846 = (w_sys_tmp5847 + w_sys_tmp5849);
	assign w_sys_tmp5847 = (r_run_copy9_j_171 * w_sys_tmp5838);
	assign w_sys_tmp5849 = 32'sh00000020;
	assign w_sys_tmp5850 = w_sub01_result_dataout;
	assign w_sys_tmp5851 = (w_sys_tmp5852 + w_sys_tmp5849);
	assign w_sys_tmp5852 = (r_run_copy8_j_170 * w_sys_tmp5838);
	assign w_sys_tmp5856 = (w_sys_tmp5857 + w_sys_tmp5859);
	assign w_sys_tmp5857 = (r_run_copy7_j_169 * w_sys_tmp5838);
	assign w_sys_tmp5859 = 32'sh00000041;
	assign w_sys_tmp5860 = (w_sys_tmp5861 + w_sys_tmp5859);
	assign w_sys_tmp5861 = (r_run_copy6_j_168 * w_sys_tmp5838);
	assign w_sys_tmp5865 = (w_sys_tmp5866 + w_sys_tmp5868);
	assign w_sys_tmp5866 = (r_run_copy5_j_167 * w_sys_tmp5838);
	assign w_sys_tmp5868 = 32'sh00000040;
	assign w_sys_tmp5870 = (w_sys_tmp5871 + w_sys_tmp5868);
	assign w_sys_tmp5871 = (r_run_copy4_j_166 * w_sys_tmp5838);
	assign w_sys_tmp5875 = (w_sys_tmp5876 + w_sys_tmp5878);
	assign w_sys_tmp5876 = (r_run_copy3_j_165 * w_sys_tmp5838);
	assign w_sys_tmp5878 = 32'sh00000061;
	assign w_sys_tmp5879 = (w_sys_tmp5880 + w_sys_tmp5878);
	assign w_sys_tmp5880 = (r_run_copy2_j_164 * w_sys_tmp5838);
	assign w_sys_tmp5884 = (w_sys_tmp5885 + w_sys_tmp5887);
	assign w_sys_tmp5885 = (r_run_copy1_j_163 * w_sys_tmp5838);
	assign w_sys_tmp5887 = 32'sh00000060;
	assign w_sys_tmp5888 = w_sub17_result_dataout;
	assign w_sys_tmp5889 = (w_sys_tmp5890 + w_sys_tmp5887);
	assign w_sys_tmp5890 = (r_run_copy0_j_162 * w_sys_tmp5838);
	assign w_sys_tmp5893 = (r_run_copy0_j_162 + w_sys_intOne);
	assign w_sys_tmp5894 = (r_run_copy1_j_163 + w_sys_intOne);
	assign w_sys_tmp5895 = (r_run_copy2_j_164 + w_sys_intOne);
	assign w_sys_tmp5896 = (r_run_copy3_j_165 + w_sys_intOne);
	assign w_sys_tmp5897 = (r_run_copy4_j_166 + w_sys_intOne);
	assign w_sys_tmp5898 = (r_run_copy5_j_167 + w_sys_intOne);
	assign w_sys_tmp5899 = (r_run_copy6_j_168 + w_sys_intOne);
	assign w_sys_tmp5900 = (r_run_copy7_j_169 + w_sys_intOne);
	assign w_sys_tmp5901 = (r_run_copy8_j_170 + w_sys_intOne);
	assign w_sys_tmp5902 = (r_run_copy9_j_171 + w_sys_intOne);
	assign w_sys_tmp5903 = (r_run_copy10_j_172 + w_sys_intOne);
	assign w_sys_tmp5904 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp6331 = 32'sh00000020;
	assign w_sys_tmp6332 = ( !w_sys_tmp6333 );
	assign w_sys_tmp6333 = (w_sys_tmp6334 < r_run_j_36);
	assign w_sys_tmp6334 = 32'sh00000031;
	assign w_sys_tmp6337 = (w_sys_tmp6338 + w_sys_tmp6340);
	assign w_sys_tmp6338 = (r_run_j_36 * w_sys_tmp6339);
	assign w_sys_tmp6339 = 32'sh00000081;
	assign w_sys_tmp6340 = 32'sh00000021;
	assign w_sys_tmp6341 = w_sub10_result_dataout;
	assign w_sys_tmp6342 = (w_sys_tmp6343 + w_sys_tmp6340);
	assign w_sys_tmp6343 = (r_run_copy10_j_183 * w_sys_tmp6339);
	assign w_sys_tmp6347 = (w_sys_tmp6348 + w_sys_tmp6350);
	assign w_sys_tmp6348 = (r_run_copy9_j_182 * w_sys_tmp6339);
	assign w_sys_tmp6350 = 32'sh00000020;
	assign w_sys_tmp6351 = w_sub02_result_dataout;
	assign w_sys_tmp6352 = (w_sys_tmp6353 + w_sys_tmp6350);
	assign w_sys_tmp6353 = (r_run_copy8_j_181 * w_sys_tmp6339);
	assign w_sys_tmp6357 = (w_sys_tmp6358 + w_sys_tmp6360);
	assign w_sys_tmp6358 = (r_run_copy7_j_180 * w_sys_tmp6339);
	assign w_sys_tmp6360 = 32'sh00000041;
	assign w_sys_tmp6361 = (w_sys_tmp6362 + w_sys_tmp6360);
	assign w_sys_tmp6362 = (r_run_copy6_j_179 * w_sys_tmp6339);
	assign w_sys_tmp6366 = (w_sys_tmp6367 + w_sys_tmp6369);
	assign w_sys_tmp6367 = (r_run_copy5_j_178 * w_sys_tmp6339);
	assign w_sys_tmp6369 = 32'sh00000040;
	assign w_sys_tmp6371 = (w_sys_tmp6372 + w_sys_tmp6369);
	assign w_sys_tmp6372 = (r_run_copy4_j_177 * w_sys_tmp6339);
	assign w_sys_tmp6376 = (w_sys_tmp6377 + w_sys_tmp6379);
	assign w_sys_tmp6377 = (r_run_copy3_j_176 * w_sys_tmp6339);
	assign w_sys_tmp6379 = 32'sh00000061;
	assign w_sys_tmp6380 = (w_sys_tmp6381 + w_sys_tmp6379);
	assign w_sys_tmp6381 = (r_run_copy2_j_175 * w_sys_tmp6339);
	assign w_sys_tmp6385 = (w_sys_tmp6386 + w_sys_tmp6388);
	assign w_sys_tmp6386 = (r_run_copy1_j_174 * w_sys_tmp6339);
	assign w_sys_tmp6388 = 32'sh00000060;
	assign w_sys_tmp6389 = w_sub18_result_dataout;
	assign w_sys_tmp6390 = (w_sys_tmp6391 + w_sys_tmp6388);
	assign w_sys_tmp6391 = (r_run_copy0_j_173 * w_sys_tmp6339);
	assign w_sys_tmp6394 = (r_run_copy0_j_173 + w_sys_intOne);
	assign w_sys_tmp6395 = (r_run_copy1_j_174 + w_sys_intOne);
	assign w_sys_tmp6396 = (r_run_copy2_j_175 + w_sys_intOne);
	assign w_sys_tmp6397 = (r_run_copy3_j_176 + w_sys_intOne);
	assign w_sys_tmp6398 = (r_run_copy4_j_177 + w_sys_intOne);
	assign w_sys_tmp6399 = (r_run_copy5_j_178 + w_sys_intOne);
	assign w_sys_tmp6400 = (r_run_copy6_j_179 + w_sys_intOne);
	assign w_sys_tmp6401 = (r_run_copy7_j_180 + w_sys_intOne);
	assign w_sys_tmp6402 = (r_run_copy8_j_181 + w_sys_intOne);
	assign w_sys_tmp6403 = (r_run_copy9_j_182 + w_sys_intOne);
	assign w_sys_tmp6404 = (r_run_copy10_j_183 + w_sys_intOne);
	assign w_sys_tmp6405 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp6832 = 32'sh00000030;
	assign w_sys_tmp6833 = ( !w_sys_tmp6834 );
	assign w_sys_tmp6834 = (w_sys_tmp6835 < r_run_j_36);
	assign w_sys_tmp6835 = 32'sh00000041;
	assign w_sys_tmp6838 = (w_sys_tmp6839 + w_sys_tmp6841);
	assign w_sys_tmp6839 = (r_run_j_36 * w_sys_tmp6840);
	assign w_sys_tmp6840 = 32'sh00000081;
	assign w_sys_tmp6841 = 32'sh00000021;
	assign w_sys_tmp6842 = w_sub11_result_dataout;
	assign w_sys_tmp6843 = (w_sys_tmp6844 + w_sys_tmp6841);
	assign w_sys_tmp6844 = (r_run_copy10_j_194 * w_sys_tmp6840);
	assign w_sys_tmp6848 = (w_sys_tmp6849 + w_sys_tmp6851);
	assign w_sys_tmp6849 = (r_run_copy9_j_193 * w_sys_tmp6840);
	assign w_sys_tmp6851 = 32'sh00000020;
	assign w_sys_tmp6852 = w_sub03_result_dataout;
	assign w_sys_tmp6853 = (w_sys_tmp6854 + w_sys_tmp6851);
	assign w_sys_tmp6854 = (r_run_copy8_j_192 * w_sys_tmp6840);
	assign w_sys_tmp6858 = (w_sys_tmp6859 + w_sys_tmp6861);
	assign w_sys_tmp6859 = (r_run_copy7_j_191 * w_sys_tmp6840);
	assign w_sys_tmp6861 = 32'sh00000041;
	assign w_sys_tmp6862 = (w_sys_tmp6863 + w_sys_tmp6861);
	assign w_sys_tmp6863 = (r_run_copy6_j_190 * w_sys_tmp6840);
	assign w_sys_tmp6867 = (w_sys_tmp6868 + w_sys_tmp6870);
	assign w_sys_tmp6868 = (r_run_copy5_j_189 * w_sys_tmp6840);
	assign w_sys_tmp6870 = 32'sh00000040;
	assign w_sys_tmp6872 = (w_sys_tmp6873 + w_sys_tmp6870);
	assign w_sys_tmp6873 = (r_run_copy4_j_188 * w_sys_tmp6840);
	assign w_sys_tmp6877 = (w_sys_tmp6878 + w_sys_tmp6880);
	assign w_sys_tmp6878 = (r_run_copy3_j_187 * w_sys_tmp6840);
	assign w_sys_tmp6880 = 32'sh00000061;
	assign w_sys_tmp6881 = (w_sys_tmp6882 + w_sys_tmp6880);
	assign w_sys_tmp6882 = (r_run_copy2_j_186 * w_sys_tmp6840);
	assign w_sys_tmp6886 = (w_sys_tmp6887 + w_sys_tmp6889);
	assign w_sys_tmp6887 = (r_run_copy1_j_185 * w_sys_tmp6840);
	assign w_sys_tmp6889 = 32'sh00000060;
	assign w_sys_tmp6890 = w_sub19_result_dataout;
	assign w_sys_tmp6891 = (w_sys_tmp6892 + w_sys_tmp6889);
	assign w_sys_tmp6892 = (r_run_copy0_j_184 * w_sys_tmp6840);
	assign w_sys_tmp6895 = (r_run_copy0_j_184 + w_sys_intOne);
	assign w_sys_tmp6896 = (r_run_copy1_j_185 + w_sys_intOne);
	assign w_sys_tmp6897 = (r_run_copy2_j_186 + w_sys_intOne);
	assign w_sys_tmp6898 = (r_run_copy3_j_187 + w_sys_intOne);
	assign w_sys_tmp6899 = (r_run_copy4_j_188 + w_sys_intOne);
	assign w_sys_tmp6900 = (r_run_copy5_j_189 + w_sys_intOne);
	assign w_sys_tmp6901 = (r_run_copy6_j_190 + w_sys_intOne);
	assign w_sys_tmp6902 = (r_run_copy7_j_191 + w_sys_intOne);
	assign w_sys_tmp6903 = (r_run_copy8_j_192 + w_sys_intOne);
	assign w_sys_tmp6904 = (r_run_copy9_j_193 + w_sys_intOne);
	assign w_sys_tmp6905 = (r_run_copy10_j_194 + w_sys_intOne);
	assign w_sys_tmp6906 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp7333 = 32'sh00000040;
	assign w_sys_tmp7334 = ( !w_sys_tmp7335 );
	assign w_sys_tmp7335 = (w_sys_tmp7336 < r_run_j_36);
	assign w_sys_tmp7336 = 32'sh00000051;
	assign w_sys_tmp7339 = (w_sys_tmp7340 + w_sys_tmp7342);
	assign w_sys_tmp7340 = (r_run_j_36 * w_sys_tmp7341);
	assign w_sys_tmp7341 = 32'sh00000081;
	assign w_sys_tmp7342 = 32'sh00000021;
	assign w_sys_tmp7343 = w_sub12_result_dataout;
	assign w_sys_tmp7344 = (w_sys_tmp7345 + w_sys_tmp7342);
	assign w_sys_tmp7345 = (r_run_copy10_j_205 * w_sys_tmp7341);
	assign w_sys_tmp7349 = (w_sys_tmp7350 + w_sys_tmp7352);
	assign w_sys_tmp7350 = (r_run_copy9_j_204 * w_sys_tmp7341);
	assign w_sys_tmp7352 = 32'sh00000020;
	assign w_sys_tmp7353 = w_sub04_result_dataout;
	assign w_sys_tmp7354 = (w_sys_tmp7355 + w_sys_tmp7352);
	assign w_sys_tmp7355 = (r_run_copy8_j_203 * w_sys_tmp7341);
	assign w_sys_tmp7359 = (w_sys_tmp7360 + w_sys_tmp7362);
	assign w_sys_tmp7360 = (r_run_copy7_j_202 * w_sys_tmp7341);
	assign w_sys_tmp7362 = 32'sh00000041;
	assign w_sys_tmp7363 = (w_sys_tmp7364 + w_sys_tmp7362);
	assign w_sys_tmp7364 = (r_run_copy6_j_201 * w_sys_tmp7341);
	assign w_sys_tmp7368 = (w_sys_tmp7369 + w_sys_tmp7371);
	assign w_sys_tmp7369 = (r_run_copy5_j_200 * w_sys_tmp7341);
	assign w_sys_tmp7371 = 32'sh00000040;
	assign w_sys_tmp7373 = (w_sys_tmp7374 + w_sys_tmp7371);
	assign w_sys_tmp7374 = (r_run_copy4_j_199 * w_sys_tmp7341);
	assign w_sys_tmp7378 = (w_sys_tmp7379 + w_sys_tmp7381);
	assign w_sys_tmp7379 = (r_run_copy3_j_198 * w_sys_tmp7341);
	assign w_sys_tmp7381 = 32'sh00000061;
	assign w_sys_tmp7382 = (w_sys_tmp7383 + w_sys_tmp7381);
	assign w_sys_tmp7383 = (r_run_copy2_j_197 * w_sys_tmp7341);
	assign w_sys_tmp7387 = (w_sys_tmp7388 + w_sys_tmp7390);
	assign w_sys_tmp7388 = (r_run_copy1_j_196 * w_sys_tmp7341);
	assign w_sys_tmp7390 = 32'sh00000060;
	assign w_sys_tmp7391 = w_sub20_result_dataout;
	assign w_sys_tmp7392 = (w_sys_tmp7393 + w_sys_tmp7390);
	assign w_sys_tmp7393 = (r_run_copy0_j_195 * w_sys_tmp7341);
	assign w_sys_tmp7396 = (r_run_copy0_j_195 + w_sys_intOne);
	assign w_sys_tmp7397 = (r_run_copy1_j_196 + w_sys_intOne);
	assign w_sys_tmp7398 = (r_run_copy2_j_197 + w_sys_intOne);
	assign w_sys_tmp7399 = (r_run_copy3_j_198 + w_sys_intOne);
	assign w_sys_tmp7400 = (r_run_copy4_j_199 + w_sys_intOne);
	assign w_sys_tmp7401 = (r_run_copy5_j_200 + w_sys_intOne);
	assign w_sys_tmp7402 = (r_run_copy6_j_201 + w_sys_intOne);
	assign w_sys_tmp7403 = (r_run_copy7_j_202 + w_sys_intOne);
	assign w_sys_tmp7404 = (r_run_copy8_j_203 + w_sys_intOne);
	assign w_sys_tmp7405 = (r_run_copy9_j_204 + w_sys_intOne);
	assign w_sys_tmp7406 = (r_run_copy10_j_205 + w_sys_intOne);
	assign w_sys_tmp7407 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp7834 = 32'sh00000050;
	assign w_sys_tmp7835 = ( !w_sys_tmp7836 );
	assign w_sys_tmp7836 = (w_sys_tmp7837 < r_run_j_36);
	assign w_sys_tmp7837 = 32'sh00000061;
	assign w_sys_tmp7840 = (w_sys_tmp7841 + w_sys_tmp7843);
	assign w_sys_tmp7841 = (r_run_j_36 * w_sys_tmp7842);
	assign w_sys_tmp7842 = 32'sh00000081;
	assign w_sys_tmp7843 = 32'sh00000021;
	assign w_sys_tmp7844 = w_sub13_result_dataout;
	assign w_sys_tmp7845 = (w_sys_tmp7846 + w_sys_tmp7843);
	assign w_sys_tmp7846 = (r_run_copy10_j_216 * w_sys_tmp7842);
	assign w_sys_tmp7850 = (w_sys_tmp7851 + w_sys_tmp7853);
	assign w_sys_tmp7851 = (r_run_copy9_j_215 * w_sys_tmp7842);
	assign w_sys_tmp7853 = 32'sh00000020;
	assign w_sys_tmp7854 = w_sub05_result_dataout;
	assign w_sys_tmp7855 = (w_sys_tmp7856 + w_sys_tmp7853);
	assign w_sys_tmp7856 = (r_run_copy8_j_214 * w_sys_tmp7842);
	assign w_sys_tmp7860 = (w_sys_tmp7861 + w_sys_tmp7863);
	assign w_sys_tmp7861 = (r_run_copy7_j_213 * w_sys_tmp7842);
	assign w_sys_tmp7863 = 32'sh00000041;
	assign w_sys_tmp7864 = (w_sys_tmp7865 + w_sys_tmp7863);
	assign w_sys_tmp7865 = (r_run_copy6_j_212 * w_sys_tmp7842);
	assign w_sys_tmp7869 = (w_sys_tmp7870 + w_sys_tmp7872);
	assign w_sys_tmp7870 = (r_run_copy5_j_211 * w_sys_tmp7842);
	assign w_sys_tmp7872 = 32'sh00000040;
	assign w_sys_tmp7874 = (w_sys_tmp7875 + w_sys_tmp7872);
	assign w_sys_tmp7875 = (r_run_copy4_j_210 * w_sys_tmp7842);
	assign w_sys_tmp7879 = (w_sys_tmp7880 + w_sys_tmp7882);
	assign w_sys_tmp7880 = (r_run_copy3_j_209 * w_sys_tmp7842);
	assign w_sys_tmp7882 = 32'sh00000061;
	assign w_sys_tmp7883 = (w_sys_tmp7884 + w_sys_tmp7882);
	assign w_sys_tmp7884 = (r_run_copy2_j_208 * w_sys_tmp7842);
	assign w_sys_tmp7888 = (w_sys_tmp7889 + w_sys_tmp7891);
	assign w_sys_tmp7889 = (r_run_copy1_j_207 * w_sys_tmp7842);
	assign w_sys_tmp7891 = 32'sh00000060;
	assign w_sys_tmp7892 = w_sub21_result_dataout;
	assign w_sys_tmp7893 = (w_sys_tmp7894 + w_sys_tmp7891);
	assign w_sys_tmp7894 = (r_run_copy0_j_206 * w_sys_tmp7842);
	assign w_sys_tmp7897 = (r_run_copy0_j_206 + w_sys_intOne);
	assign w_sys_tmp7898 = (r_run_copy1_j_207 + w_sys_intOne);
	assign w_sys_tmp7899 = (r_run_copy2_j_208 + w_sys_intOne);
	assign w_sys_tmp7900 = (r_run_copy3_j_209 + w_sys_intOne);
	assign w_sys_tmp7901 = (r_run_copy4_j_210 + w_sys_intOne);
	assign w_sys_tmp7902 = (r_run_copy5_j_211 + w_sys_intOne);
	assign w_sys_tmp7903 = (r_run_copy6_j_212 + w_sys_intOne);
	assign w_sys_tmp7904 = (r_run_copy7_j_213 + w_sys_intOne);
	assign w_sys_tmp7905 = (r_run_copy8_j_214 + w_sys_intOne);
	assign w_sys_tmp7906 = (r_run_copy9_j_215 + w_sys_intOne);
	assign w_sys_tmp7907 = (r_run_copy10_j_216 + w_sys_intOne);
	assign w_sys_tmp7908 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp8335 = 32'sh00000060;
	assign w_sys_tmp8336 = ( !w_sys_tmp8337 );
	assign w_sys_tmp8337 = (w_sys_tmp8338 < r_run_j_36);
	assign w_sys_tmp8338 = 32'sh00000071;
	assign w_sys_tmp8341 = (w_sys_tmp8342 + w_sys_tmp8344);
	assign w_sys_tmp8342 = (r_run_j_36 * w_sys_tmp8343);
	assign w_sys_tmp8343 = 32'sh00000081;
	assign w_sys_tmp8344 = 32'sh00000021;
	assign w_sys_tmp8345 = w_sub14_result_dataout;
	assign w_sys_tmp8346 = (w_sys_tmp8347 + w_sys_tmp8344);
	assign w_sys_tmp8347 = (r_run_copy10_j_227 * w_sys_tmp8343);
	assign w_sys_tmp8351 = (w_sys_tmp8352 + w_sys_tmp8354);
	assign w_sys_tmp8352 = (r_run_copy9_j_226 * w_sys_tmp8343);
	assign w_sys_tmp8354 = 32'sh00000020;
	assign w_sys_tmp8355 = w_sub06_result_dataout;
	assign w_sys_tmp8356 = (w_sys_tmp8357 + w_sys_tmp8354);
	assign w_sys_tmp8357 = (r_run_copy8_j_225 * w_sys_tmp8343);
	assign w_sys_tmp8361 = (w_sys_tmp8362 + w_sys_tmp8364);
	assign w_sys_tmp8362 = (r_run_copy7_j_224 * w_sys_tmp8343);
	assign w_sys_tmp8364 = 32'sh00000041;
	assign w_sys_tmp8365 = (w_sys_tmp8366 + w_sys_tmp8364);
	assign w_sys_tmp8366 = (r_run_copy6_j_223 * w_sys_tmp8343);
	assign w_sys_tmp8370 = (w_sys_tmp8371 + w_sys_tmp8373);
	assign w_sys_tmp8371 = (r_run_copy5_j_222 * w_sys_tmp8343);
	assign w_sys_tmp8373 = 32'sh00000040;
	assign w_sys_tmp8375 = (w_sys_tmp8376 + w_sys_tmp8373);
	assign w_sys_tmp8376 = (r_run_copy4_j_221 * w_sys_tmp8343);
	assign w_sys_tmp8380 = (w_sys_tmp8381 + w_sys_tmp8383);
	assign w_sys_tmp8381 = (r_run_copy3_j_220 * w_sys_tmp8343);
	assign w_sys_tmp8383 = 32'sh00000061;
	assign w_sys_tmp8384 = (w_sys_tmp8385 + w_sys_tmp8383);
	assign w_sys_tmp8385 = (r_run_copy2_j_219 * w_sys_tmp8343);
	assign w_sys_tmp8389 = (w_sys_tmp8390 + w_sys_tmp8392);
	assign w_sys_tmp8390 = (r_run_copy1_j_218 * w_sys_tmp8343);
	assign w_sys_tmp8392 = 32'sh00000060;
	assign w_sys_tmp8393 = w_sub22_result_dataout;
	assign w_sys_tmp8394 = (w_sys_tmp8395 + w_sys_tmp8392);
	assign w_sys_tmp8395 = (r_run_copy0_j_217 * w_sys_tmp8343);
	assign w_sys_tmp8398 = (r_run_copy0_j_217 + w_sys_intOne);
	assign w_sys_tmp8399 = (r_run_copy1_j_218 + w_sys_intOne);
	assign w_sys_tmp8400 = (r_run_copy2_j_219 + w_sys_intOne);
	assign w_sys_tmp8401 = (r_run_copy3_j_220 + w_sys_intOne);
	assign w_sys_tmp8402 = (r_run_copy4_j_221 + w_sys_intOne);
	assign w_sys_tmp8403 = (r_run_copy5_j_222 + w_sys_intOne);
	assign w_sys_tmp8404 = (r_run_copy6_j_223 + w_sys_intOne);
	assign w_sys_tmp8405 = (r_run_copy7_j_224 + w_sys_intOne);
	assign w_sys_tmp8406 = (r_run_copy8_j_225 + w_sys_intOne);
	assign w_sys_tmp8407 = (r_run_copy9_j_226 + w_sys_intOne);
	assign w_sys_tmp8408 = (r_run_copy10_j_227 + w_sys_intOne);
	assign w_sys_tmp8409 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp8836 = 32'sh00000070;
	assign w_sys_tmp8837 = ( !w_sys_tmp8838 );
	assign w_sys_tmp8838 = (w_sys_tmp8839 < r_run_j_36);
	assign w_sys_tmp8839 = 32'sh00000081;
	assign w_sys_tmp8842 = (w_sys_tmp8843 + w_sys_tmp8845);
	assign w_sys_tmp8843 = (r_run_j_36 * w_sys_tmp8844);
	assign w_sys_tmp8844 = 32'sh00000081;
	assign w_sys_tmp8845 = 32'sh00000021;
	assign w_sys_tmp8846 = w_sub15_result_dataout;
	assign w_sys_tmp8847 = (w_sys_tmp8848 + w_sys_tmp8845);
	assign w_sys_tmp8848 = (r_run_copy10_j_238 * w_sys_tmp8844);
	assign w_sys_tmp8852 = (w_sys_tmp8853 + w_sys_tmp8855);
	assign w_sys_tmp8853 = (r_run_copy9_j_237 * w_sys_tmp8844);
	assign w_sys_tmp8855 = 32'sh00000020;
	assign w_sys_tmp8856 = w_sub07_result_dataout;
	assign w_sys_tmp8857 = (w_sys_tmp8858 + w_sys_tmp8855);
	assign w_sys_tmp8858 = (r_run_copy8_j_236 * w_sys_tmp8844);
	assign w_sys_tmp8862 = (w_sys_tmp8863 + w_sys_tmp8865);
	assign w_sys_tmp8863 = (r_run_copy7_j_235 * w_sys_tmp8844);
	assign w_sys_tmp8865 = 32'sh00000041;
	assign w_sys_tmp8866 = (w_sys_tmp8867 + w_sys_tmp8865);
	assign w_sys_tmp8867 = (r_run_copy6_j_234 * w_sys_tmp8844);
	assign w_sys_tmp8871 = (w_sys_tmp8872 + w_sys_tmp8874);
	assign w_sys_tmp8872 = (r_run_copy5_j_233 * w_sys_tmp8844);
	assign w_sys_tmp8874 = 32'sh00000040;
	assign w_sys_tmp8876 = (w_sys_tmp8877 + w_sys_tmp8874);
	assign w_sys_tmp8877 = (r_run_copy4_j_232 * w_sys_tmp8844);
	assign w_sys_tmp8881 = (w_sys_tmp8882 + w_sys_tmp8884);
	assign w_sys_tmp8882 = (r_run_copy3_j_231 * w_sys_tmp8844);
	assign w_sys_tmp8884 = 32'sh00000061;
	assign w_sys_tmp8885 = (w_sys_tmp8886 + w_sys_tmp8884);
	assign w_sys_tmp8886 = (r_run_copy2_j_230 * w_sys_tmp8844);
	assign w_sys_tmp8890 = (w_sys_tmp8891 + w_sys_tmp8893);
	assign w_sys_tmp8891 = (r_run_copy1_j_229 * w_sys_tmp8844);
	assign w_sys_tmp8893 = 32'sh00000060;
	assign w_sys_tmp8894 = w_sub16_result_dataout;
	assign w_sys_tmp8895 = (w_sys_tmp8896 + w_sys_tmp8893);
	assign w_sys_tmp8896 = (r_run_copy0_j_228 * w_sys_tmp8844);
	assign w_sys_tmp8899 = (r_run_copy0_j_228 + w_sys_intOne);
	assign w_sys_tmp8900 = (r_run_copy1_j_229 + w_sys_intOne);
	assign w_sys_tmp8901 = (r_run_copy2_j_230 + w_sys_intOne);
	assign w_sys_tmp8902 = (r_run_copy3_j_231 + w_sys_intOne);
	assign w_sys_tmp8903 = (r_run_copy4_j_232 + w_sys_intOne);
	assign w_sys_tmp8904 = (r_run_copy5_j_233 + w_sys_intOne);
	assign w_sys_tmp8905 = (r_run_copy6_j_234 + w_sys_intOne);
	assign w_sys_tmp8906 = (r_run_copy7_j_235 + w_sys_intOne);
	assign w_sys_tmp8907 = (r_run_copy8_j_236 + w_sys_intOne);
	assign w_sys_tmp8908 = (r_run_copy9_j_237 + w_sys_intOne);
	assign w_sys_tmp8909 = (r_run_copy10_j_238 + w_sys_intOne);
	assign w_sys_tmp8910 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp9325 = 32'sh00000002;
	assign w_sys_tmp9326 = ( !w_sys_tmp9327 );
	assign w_sys_tmp9327 = (w_sys_tmp9328 < r_run_k_35);
	assign w_sys_tmp9328 = 32'sh00000020;
	assign w_sys_tmp9329 = (r_run_k_35 + w_sys_intOne);
	assign w_sys_tmp9330 = 32'sh00000002;
	assign w_sys_tmp9331 = ( !w_sys_tmp9332 );
	assign w_sys_tmp9332 = (w_sys_tmp9333 < r_run_j_36);
	assign w_sys_tmp9333 = 32'sh00000010;
	assign w_sys_tmp9336 = (w_sys_tmp9337 + r_run_k_35);
	assign w_sys_tmp9337 = (r_run_j_36 * w_sys_tmp9338);
	assign w_sys_tmp9338 = 32'sh00000081;
	assign w_sys_tmp9339 = w_sub00_result_dataout;
	assign w_sys_tmp9340 = (w_sys_tmp9341 + r_run_k_35);
	assign w_sys_tmp9341 = (r_run_copy0_j_239 * w_sys_tmp9338);
	assign w_sys_tmp9343 = (r_run_copy0_j_239 + w_sys_intOne);
	assign w_sys_tmp9344 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp9405 = 32'sh00000011;
	assign w_sys_tmp9406 = ( !w_sys_tmp9407 );
	assign w_sys_tmp9407 = (w_sys_tmp9408 < r_run_j_36);
	assign w_sys_tmp9408 = 32'sh00000020;
	assign w_sys_tmp9410 = (r_run_j_36 - w_sys_tmp9411);
	assign w_sys_tmp9411 = 32'sh0000000f;
	assign w_sys_tmp9413 = (w_sys_tmp9414 + r_run_k_35);
	assign w_sys_tmp9414 = (r_run_copy1_j_241 * w_sys_tmp9415);
	assign w_sys_tmp9415 = 32'sh00000081;
	assign w_sys_tmp9416 = w_sub01_result_dataout;
	assign w_sys_tmp9417 = (w_sys_tmp9418 + r_run_k_35);
	assign w_sys_tmp9418 = (r_run_copy0_j_240 * w_sys_tmp9415);
	assign w_sys_tmp9420 = (r_run_copy0_j_240 + w_sys_intOne);
	assign w_sys_tmp9421 = (r_run_copy1_j_241 + w_sys_intOne);
	assign w_sys_tmp9422 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp9501 = 32'sh00000021;
	assign w_sys_tmp9502 = ( !w_sys_tmp9503 );
	assign w_sys_tmp9503 = (w_sys_tmp9504 < r_run_j_36);
	assign w_sys_tmp9504 = 32'sh00000030;
	assign w_sys_tmp9506 = (r_run_j_36 - w_sys_tmp9507);
	assign w_sys_tmp9507 = 32'sh0000001f;
	assign w_sys_tmp9509 = (w_sys_tmp9510 + r_run_k_35);
	assign w_sys_tmp9510 = (r_run_copy1_j_243 * w_sys_tmp9511);
	assign w_sys_tmp9511 = 32'sh00000081;
	assign w_sys_tmp9512 = w_sub02_result_dataout;
	assign w_sys_tmp9513 = (w_sys_tmp9514 + r_run_k_35);
	assign w_sys_tmp9514 = (r_run_copy0_j_242 * w_sys_tmp9511);
	assign w_sys_tmp9516 = (r_run_copy0_j_242 + w_sys_intOne);
	assign w_sys_tmp9517 = (r_run_copy1_j_243 + w_sys_intOne);
	assign w_sys_tmp9518 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp9597 = 32'sh00000031;
	assign w_sys_tmp9598 = ( !w_sys_tmp9599 );
	assign w_sys_tmp9599 = (w_sys_tmp9600 < r_run_j_36);
	assign w_sys_tmp9600 = 32'sh00000040;
	assign w_sys_tmp9602 = (r_run_j_36 - w_sys_tmp9603);
	assign w_sys_tmp9603 = 32'sh0000002f;
	assign w_sys_tmp9605 = (w_sys_tmp9606 + r_run_k_35);
	assign w_sys_tmp9606 = (r_run_copy1_j_245 * w_sys_tmp9607);
	assign w_sys_tmp9607 = 32'sh00000081;
	assign w_sys_tmp9608 = w_sub03_result_dataout;
	assign w_sys_tmp9609 = (w_sys_tmp9610 + r_run_k_35);
	assign w_sys_tmp9610 = (r_run_copy0_j_244 * w_sys_tmp9607);
	assign w_sys_tmp9612 = (r_run_copy0_j_244 + w_sys_intOne);
	assign w_sys_tmp9613 = (r_run_copy1_j_245 + w_sys_intOne);
	assign w_sys_tmp9614 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp9693 = 32'sh00000041;
	assign w_sys_tmp9694 = ( !w_sys_tmp9695 );
	assign w_sys_tmp9695 = (w_sys_tmp9696 < r_run_j_36);
	assign w_sys_tmp9696 = 32'sh00000050;
	assign w_sys_tmp9698 = (r_run_j_36 - w_sys_tmp9699);
	assign w_sys_tmp9699 = 32'sh0000003f;
	assign w_sys_tmp9701 = (w_sys_tmp9702 + r_run_k_35);
	assign w_sys_tmp9702 = (r_run_copy1_j_247 * w_sys_tmp9703);
	assign w_sys_tmp9703 = 32'sh00000081;
	assign w_sys_tmp9704 = w_sub04_result_dataout;
	assign w_sys_tmp9705 = (w_sys_tmp9706 + r_run_k_35);
	assign w_sys_tmp9706 = (r_run_copy0_j_246 * w_sys_tmp9703);
	assign w_sys_tmp9708 = (r_run_copy0_j_246 + w_sys_intOne);
	assign w_sys_tmp9709 = (r_run_copy1_j_247 + w_sys_intOne);
	assign w_sys_tmp9710 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp9789 = 32'sh00000051;
	assign w_sys_tmp9790 = ( !w_sys_tmp9791 );
	assign w_sys_tmp9791 = (w_sys_tmp9792 < r_run_j_36);
	assign w_sys_tmp9792 = 32'sh00000060;
	assign w_sys_tmp9794 = (r_run_j_36 - w_sys_tmp9795);
	assign w_sys_tmp9795 = 32'sh0000004f;
	assign w_sys_tmp9797 = (w_sys_tmp9798 + r_run_k_35);
	assign w_sys_tmp9798 = (r_run_copy1_j_249 * w_sys_tmp9799);
	assign w_sys_tmp9799 = 32'sh00000081;
	assign w_sys_tmp9800 = w_sub05_result_dataout;
	assign w_sys_tmp9801 = (w_sys_tmp9802 + r_run_k_35);
	assign w_sys_tmp9802 = (r_run_copy0_j_248 * w_sys_tmp9799);
	assign w_sys_tmp9804 = (r_run_copy0_j_248 + w_sys_intOne);
	assign w_sys_tmp9805 = (r_run_copy1_j_249 + w_sys_intOne);
	assign w_sys_tmp9806 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp9885 = 32'sh00000061;
	assign w_sys_tmp9886 = ( !w_sys_tmp9887 );
	assign w_sys_tmp9887 = (w_sys_tmp9888 < r_run_j_36);
	assign w_sys_tmp9888 = 32'sh00000070;
	assign w_sys_tmp9890 = (r_run_j_36 - w_sys_tmp9891);
	assign w_sys_tmp9891 = 32'sh0000005f;
	assign w_sys_tmp9893 = (w_sys_tmp9894 + r_run_k_35);
	assign w_sys_tmp9894 = (r_run_copy1_j_251 * w_sys_tmp9895);
	assign w_sys_tmp9895 = 32'sh00000081;
	assign w_sys_tmp9896 = w_sub06_result_dataout;
	assign w_sys_tmp9897 = (w_sys_tmp9898 + r_run_k_35);
	assign w_sys_tmp9898 = (r_run_copy0_j_250 * w_sys_tmp9895);
	assign w_sys_tmp9900 = (r_run_copy0_j_250 + w_sys_intOne);
	assign w_sys_tmp9901 = (r_run_copy1_j_251 + w_sys_intOne);
	assign w_sys_tmp9902 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp9981 = 32'sh00000071;
	assign w_sys_tmp9982 = ( !w_sys_tmp9983 );
	assign w_sys_tmp9983 = (w_sys_tmp9984 < r_run_j_36);
	assign w_sys_tmp9984 = 32'sh00000080;
	assign w_sys_tmp9986 = (r_run_j_36 - w_sys_tmp9987);
	assign w_sys_tmp9987 = 32'sh0000006f;
	assign w_sys_tmp9989 = (w_sys_tmp9990 + r_run_k_35);
	assign w_sys_tmp9990 = (r_run_copy1_j_253 * w_sys_tmp9991);
	assign w_sys_tmp9991 = 32'sh00000081;
	assign w_sys_tmp9992 = w_sub07_result_dataout;
	assign w_sys_tmp9993 = (w_sys_tmp9994 + r_run_k_35);
	assign w_sys_tmp9994 = (r_run_copy0_j_252 * w_sys_tmp9991);
	assign w_sys_tmp9996 = (r_run_copy0_j_252 + w_sys_intOne);
	assign w_sys_tmp9997 = (r_run_copy1_j_253 + w_sys_intOne);
	assign w_sys_tmp9998 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp10077 = 32'sh00000021;
	assign w_sys_tmp10078 = ( !w_sys_tmp10079 );
	assign w_sys_tmp10079 = (w_sys_tmp10080 < r_run_k_35);
	assign w_sys_tmp10080 = 32'sh00000040;
	assign w_sys_tmp10081 = (r_run_k_35 + w_sys_intOne);
	assign w_sys_tmp10082 = 32'sh00000002;
	assign w_sys_tmp10083 = ( !w_sys_tmp10084 );
	assign w_sys_tmp10084 = (w_sys_tmp10085 < r_run_j_36);
	assign w_sys_tmp10085 = 32'sh00000010;
	assign w_sys_tmp10088 = (w_sys_tmp10089 + r_run_k_35);
	assign w_sys_tmp10089 = (r_run_j_36 * w_sys_tmp10090);
	assign w_sys_tmp10090 = 32'sh00000081;
	assign w_sys_tmp10091 = w_sub08_result_dataout;
	assign w_sys_tmp10092 = (w_sys_tmp10093 + r_run_k_35);
	assign w_sys_tmp10093 = (r_run_copy0_j_254 * w_sys_tmp10090);
	assign w_sys_tmp10095 = (r_run_copy0_j_254 + w_sys_intOne);
	assign w_sys_tmp10096 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp10157 = 32'sh00000011;
	assign w_sys_tmp10158 = ( !w_sys_tmp10159 );
	assign w_sys_tmp10159 = (w_sys_tmp10160 < r_run_j_36);
	assign w_sys_tmp10160 = 32'sh00000020;
	assign w_sys_tmp10162 = (r_run_j_36 - w_sys_tmp10163);
	assign w_sys_tmp10163 = 32'sh0000000f;
	assign w_sys_tmp10165 = (w_sys_tmp10166 + r_run_k_35);
	assign w_sys_tmp10166 = (r_run_copy1_j_256 * w_sys_tmp10167);
	assign w_sys_tmp10167 = 32'sh00000081;
	assign w_sys_tmp10168 = w_sub09_result_dataout;
	assign w_sys_tmp10169 = (w_sys_tmp10170 + r_run_k_35);
	assign w_sys_tmp10170 = (r_run_copy0_j_255 * w_sys_tmp10167);
	assign w_sys_tmp10172 = (r_run_copy0_j_255 + w_sys_intOne);
	assign w_sys_tmp10173 = (r_run_copy1_j_256 + w_sys_intOne);
	assign w_sys_tmp10174 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp10253 = 32'sh00000021;
	assign w_sys_tmp10254 = ( !w_sys_tmp10255 );
	assign w_sys_tmp10255 = (w_sys_tmp10256 < r_run_j_36);
	assign w_sys_tmp10256 = 32'sh00000030;
	assign w_sys_tmp10258 = (r_run_j_36 - w_sys_tmp10259);
	assign w_sys_tmp10259 = 32'sh0000001f;
	assign w_sys_tmp10261 = (w_sys_tmp10262 + r_run_k_35);
	assign w_sys_tmp10262 = (r_run_copy1_j_258 * w_sys_tmp10263);
	assign w_sys_tmp10263 = 32'sh00000081;
	assign w_sys_tmp10264 = w_sub10_result_dataout;
	assign w_sys_tmp10265 = (w_sys_tmp10266 + r_run_k_35);
	assign w_sys_tmp10266 = (r_run_copy0_j_257 * w_sys_tmp10263);
	assign w_sys_tmp10268 = (r_run_copy0_j_257 + w_sys_intOne);
	assign w_sys_tmp10269 = (r_run_copy1_j_258 + w_sys_intOne);
	assign w_sys_tmp10270 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp10349 = 32'sh00000031;
	assign w_sys_tmp10350 = ( !w_sys_tmp10351 );
	assign w_sys_tmp10351 = (w_sys_tmp10352 < r_run_j_36);
	assign w_sys_tmp10352 = 32'sh00000040;
	assign w_sys_tmp10354 = (r_run_j_36 - w_sys_tmp10355);
	assign w_sys_tmp10355 = 32'sh0000002f;
	assign w_sys_tmp10357 = (w_sys_tmp10358 + r_run_k_35);
	assign w_sys_tmp10358 = (r_run_copy1_j_260 * w_sys_tmp10359);
	assign w_sys_tmp10359 = 32'sh00000081;
	assign w_sys_tmp10360 = w_sub11_result_dataout;
	assign w_sys_tmp10361 = (w_sys_tmp10362 + r_run_k_35);
	assign w_sys_tmp10362 = (r_run_copy0_j_259 * w_sys_tmp10359);
	assign w_sys_tmp10364 = (r_run_copy0_j_259 + w_sys_intOne);
	assign w_sys_tmp10365 = (r_run_copy1_j_260 + w_sys_intOne);
	assign w_sys_tmp10366 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp10445 = 32'sh00000041;
	assign w_sys_tmp10446 = ( !w_sys_tmp10447 );
	assign w_sys_tmp10447 = (w_sys_tmp10448 < r_run_j_36);
	assign w_sys_tmp10448 = 32'sh00000050;
	assign w_sys_tmp10450 = (r_run_j_36 - w_sys_tmp10451);
	assign w_sys_tmp10451 = 32'sh0000003f;
	assign w_sys_tmp10453 = (w_sys_tmp10454 + r_run_k_35);
	assign w_sys_tmp10454 = (r_run_copy1_j_262 * w_sys_tmp10455);
	assign w_sys_tmp10455 = 32'sh00000081;
	assign w_sys_tmp10456 = w_sub12_result_dataout;
	assign w_sys_tmp10457 = (w_sys_tmp10458 + r_run_k_35);
	assign w_sys_tmp10458 = (r_run_copy0_j_261 * w_sys_tmp10455);
	assign w_sys_tmp10460 = (r_run_copy0_j_261 + w_sys_intOne);
	assign w_sys_tmp10461 = (r_run_copy1_j_262 + w_sys_intOne);
	assign w_sys_tmp10462 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp10541 = 32'sh00000051;
	assign w_sys_tmp10542 = ( !w_sys_tmp10543 );
	assign w_sys_tmp10543 = (w_sys_tmp10544 < r_run_j_36);
	assign w_sys_tmp10544 = 32'sh00000060;
	assign w_sys_tmp10546 = (r_run_j_36 - w_sys_tmp10547);
	assign w_sys_tmp10547 = 32'sh0000004f;
	assign w_sys_tmp10549 = (w_sys_tmp10550 + r_run_k_35);
	assign w_sys_tmp10550 = (r_run_copy1_j_264 * w_sys_tmp10551);
	assign w_sys_tmp10551 = 32'sh00000081;
	assign w_sys_tmp10552 = w_sub13_result_dataout;
	assign w_sys_tmp10553 = (w_sys_tmp10554 + r_run_k_35);
	assign w_sys_tmp10554 = (r_run_copy0_j_263 * w_sys_tmp10551);
	assign w_sys_tmp10556 = (r_run_copy0_j_263 + w_sys_intOne);
	assign w_sys_tmp10557 = (r_run_copy1_j_264 + w_sys_intOne);
	assign w_sys_tmp10558 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp10637 = 32'sh00000061;
	assign w_sys_tmp10638 = ( !w_sys_tmp10639 );
	assign w_sys_tmp10639 = (w_sys_tmp10640 < r_run_j_36);
	assign w_sys_tmp10640 = 32'sh00000070;
	assign w_sys_tmp10642 = (r_run_j_36 - w_sys_tmp10643);
	assign w_sys_tmp10643 = 32'sh0000005f;
	assign w_sys_tmp10645 = (w_sys_tmp10646 + r_run_k_35);
	assign w_sys_tmp10646 = (r_run_copy1_j_266 * w_sys_tmp10647);
	assign w_sys_tmp10647 = 32'sh00000081;
	assign w_sys_tmp10648 = w_sub14_result_dataout;
	assign w_sys_tmp10649 = (w_sys_tmp10650 + r_run_k_35);
	assign w_sys_tmp10650 = (r_run_copy0_j_265 * w_sys_tmp10647);
	assign w_sys_tmp10652 = (r_run_copy0_j_265 + w_sys_intOne);
	assign w_sys_tmp10653 = (r_run_copy1_j_266 + w_sys_intOne);
	assign w_sys_tmp10654 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp10733 = 32'sh00000071;
	assign w_sys_tmp10734 = ( !w_sys_tmp10735 );
	assign w_sys_tmp10735 = (w_sys_tmp10736 < r_run_j_36);
	assign w_sys_tmp10736 = 32'sh00000080;
	assign w_sys_tmp10738 = (r_run_j_36 - w_sys_tmp10739);
	assign w_sys_tmp10739 = 32'sh0000006f;
	assign w_sys_tmp10741 = (w_sys_tmp10742 + r_run_k_35);
	assign w_sys_tmp10742 = (r_run_copy1_j_268 * w_sys_tmp10743);
	assign w_sys_tmp10743 = 32'sh00000081;
	assign w_sys_tmp10744 = w_sub15_result_dataout;
	assign w_sys_tmp10745 = (w_sys_tmp10746 + r_run_k_35);
	assign w_sys_tmp10746 = (r_run_copy0_j_267 * w_sys_tmp10743);
	assign w_sys_tmp10748 = (r_run_copy0_j_267 + w_sys_intOne);
	assign w_sys_tmp10749 = (r_run_copy1_j_268 + w_sys_intOne);
	assign w_sys_tmp10750 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp10829 = 32'sh00000041;
	assign w_sys_tmp10830 = ( !w_sys_tmp10831 );
	assign w_sys_tmp10831 = (w_sys_tmp10832 < r_run_k_35);
	assign w_sys_tmp10832 = 32'sh00000060;
	assign w_sys_tmp10833 = (r_run_k_35 + w_sys_intOne);
	assign w_sys_tmp10834 = 32'sh00000002;
	assign w_sys_tmp10835 = ( !w_sys_tmp10836 );
	assign w_sys_tmp10836 = (w_sys_tmp10837 < r_run_j_36);
	assign w_sys_tmp10837 = 32'sh00000010;
	assign w_sys_tmp10840 = (w_sys_tmp10841 + r_run_k_35);
	assign w_sys_tmp10841 = (r_run_j_36 * w_sys_tmp10842);
	assign w_sys_tmp10842 = 32'sh00000081;
	assign w_sys_tmp10843 = w_sub16_result_dataout;
	assign w_sys_tmp10844 = (w_sys_tmp10845 + r_run_k_35);
	assign w_sys_tmp10845 = (r_run_copy0_j_269 * w_sys_tmp10842);
	assign w_sys_tmp10847 = (r_run_copy0_j_269 + w_sys_intOne);
	assign w_sys_tmp10848 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp10909 = 32'sh00000011;
	assign w_sys_tmp10910 = ( !w_sys_tmp10911 );
	assign w_sys_tmp10911 = (w_sys_tmp10912 < r_run_j_36);
	assign w_sys_tmp10912 = 32'sh00000020;
	assign w_sys_tmp10914 = (r_run_j_36 - w_sys_tmp10915);
	assign w_sys_tmp10915 = 32'sh0000000f;
	assign w_sys_tmp10917 = (w_sys_tmp10918 + r_run_k_35);
	assign w_sys_tmp10918 = (r_run_copy1_j_271 * w_sys_tmp10919);
	assign w_sys_tmp10919 = 32'sh00000081;
	assign w_sys_tmp10920 = w_sub17_result_dataout;
	assign w_sys_tmp10921 = (w_sys_tmp10922 + r_run_k_35);
	assign w_sys_tmp10922 = (r_run_copy0_j_270 * w_sys_tmp10919);
	assign w_sys_tmp10924 = (r_run_copy0_j_270 + w_sys_intOne);
	assign w_sys_tmp10925 = (r_run_copy1_j_271 + w_sys_intOne);
	assign w_sys_tmp10926 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp11005 = 32'sh00000021;
	assign w_sys_tmp11006 = ( !w_sys_tmp11007 );
	assign w_sys_tmp11007 = (w_sys_tmp11008 < r_run_j_36);
	assign w_sys_tmp11008 = 32'sh00000030;
	assign w_sys_tmp11010 = (r_run_j_36 - w_sys_tmp11011);
	assign w_sys_tmp11011 = 32'sh0000001f;
	assign w_sys_tmp11013 = (w_sys_tmp11014 + r_run_k_35);
	assign w_sys_tmp11014 = (r_run_copy1_j_273 * w_sys_tmp11015);
	assign w_sys_tmp11015 = 32'sh00000081;
	assign w_sys_tmp11016 = w_sub18_result_dataout;
	assign w_sys_tmp11017 = (w_sys_tmp11018 + r_run_k_35);
	assign w_sys_tmp11018 = (r_run_copy0_j_272 * w_sys_tmp11015);
	assign w_sys_tmp11020 = (r_run_copy0_j_272 + w_sys_intOne);
	assign w_sys_tmp11021 = (r_run_copy1_j_273 + w_sys_intOne);
	assign w_sys_tmp11022 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp11101 = 32'sh00000031;
	assign w_sys_tmp11102 = ( !w_sys_tmp11103 );
	assign w_sys_tmp11103 = (w_sys_tmp11104 < r_run_j_36);
	assign w_sys_tmp11104 = 32'sh00000040;
	assign w_sys_tmp11106 = (r_run_j_36 - w_sys_tmp11107);
	assign w_sys_tmp11107 = 32'sh0000002f;
	assign w_sys_tmp11109 = (w_sys_tmp11110 + r_run_k_35);
	assign w_sys_tmp11110 = (r_run_copy1_j_275 * w_sys_tmp11111);
	assign w_sys_tmp11111 = 32'sh00000081;
	assign w_sys_tmp11112 = w_sub19_result_dataout;
	assign w_sys_tmp11113 = (w_sys_tmp11114 + r_run_k_35);
	assign w_sys_tmp11114 = (r_run_copy0_j_274 * w_sys_tmp11111);
	assign w_sys_tmp11116 = (r_run_copy0_j_274 + w_sys_intOne);
	assign w_sys_tmp11117 = (r_run_copy1_j_275 + w_sys_intOne);
	assign w_sys_tmp11118 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp11197 = 32'sh00000041;
	assign w_sys_tmp11198 = ( !w_sys_tmp11199 );
	assign w_sys_tmp11199 = (w_sys_tmp11200 < r_run_j_36);
	assign w_sys_tmp11200 = 32'sh00000050;
	assign w_sys_tmp11202 = (r_run_j_36 - w_sys_tmp11203);
	assign w_sys_tmp11203 = 32'sh0000003f;
	assign w_sys_tmp11205 = (w_sys_tmp11206 + r_run_k_35);
	assign w_sys_tmp11206 = (r_run_copy1_j_277 * w_sys_tmp11207);
	assign w_sys_tmp11207 = 32'sh00000081;
	assign w_sys_tmp11208 = w_sub20_result_dataout;
	assign w_sys_tmp11209 = (w_sys_tmp11210 + r_run_k_35);
	assign w_sys_tmp11210 = (r_run_copy0_j_276 * w_sys_tmp11207);
	assign w_sys_tmp11212 = (r_run_copy0_j_276 + w_sys_intOne);
	assign w_sys_tmp11213 = (r_run_copy1_j_277 + w_sys_intOne);
	assign w_sys_tmp11214 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp11293 = 32'sh00000051;
	assign w_sys_tmp11294 = ( !w_sys_tmp11295 );
	assign w_sys_tmp11295 = (w_sys_tmp11296 < r_run_j_36);
	assign w_sys_tmp11296 = 32'sh00000060;
	assign w_sys_tmp11298 = (r_run_j_36 - w_sys_tmp11299);
	assign w_sys_tmp11299 = 32'sh0000004f;
	assign w_sys_tmp11301 = (w_sys_tmp11302 + r_run_k_35);
	assign w_sys_tmp11302 = (r_run_copy1_j_279 * w_sys_tmp11303);
	assign w_sys_tmp11303 = 32'sh00000081;
	assign w_sys_tmp11304 = w_sub21_result_dataout;
	assign w_sys_tmp11305 = (w_sys_tmp11306 + r_run_k_35);
	assign w_sys_tmp11306 = (r_run_copy0_j_278 * w_sys_tmp11303);
	assign w_sys_tmp11308 = (r_run_copy0_j_278 + w_sys_intOne);
	assign w_sys_tmp11309 = (r_run_copy1_j_279 + w_sys_intOne);
	assign w_sys_tmp11310 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp11389 = 32'sh00000061;
	assign w_sys_tmp11390 = ( !w_sys_tmp11391 );
	assign w_sys_tmp11391 = (w_sys_tmp11392 < r_run_j_36);
	assign w_sys_tmp11392 = 32'sh00000070;
	assign w_sys_tmp11394 = (r_run_j_36 - w_sys_tmp11395);
	assign w_sys_tmp11395 = 32'sh0000005f;
	assign w_sys_tmp11397 = (w_sys_tmp11398 + r_run_k_35);
	assign w_sys_tmp11398 = (r_run_copy1_j_281 * w_sys_tmp11399);
	assign w_sys_tmp11399 = 32'sh00000081;
	assign w_sys_tmp11400 = w_sub22_result_dataout;
	assign w_sys_tmp11401 = (w_sys_tmp11402 + r_run_k_35);
	assign w_sys_tmp11402 = (r_run_copy0_j_280 * w_sys_tmp11399);
	assign w_sys_tmp11404 = (r_run_copy0_j_280 + w_sys_intOne);
	assign w_sys_tmp11405 = (r_run_copy1_j_281 + w_sys_intOne);
	assign w_sys_tmp11406 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp11485 = 32'sh00000071;
	assign w_sys_tmp11486 = ( !w_sys_tmp11487 );
	assign w_sys_tmp11487 = (w_sys_tmp11488 < r_run_j_36);
	assign w_sys_tmp11488 = 32'sh00000080;
	assign w_sys_tmp11490 = (r_run_j_36 - w_sys_tmp11491);
	assign w_sys_tmp11491 = 32'sh0000006f;
	assign w_sys_tmp11493 = (w_sys_tmp11494 + r_run_k_35);
	assign w_sys_tmp11494 = (r_run_copy1_j_283 * w_sys_tmp11495);
	assign w_sys_tmp11495 = 32'sh00000081;
	assign w_sys_tmp11496 = w_sub23_result_dataout;
	assign w_sys_tmp11497 = (w_sys_tmp11498 + r_run_k_35);
	assign w_sys_tmp11498 = (r_run_copy0_j_282 * w_sys_tmp11495);
	assign w_sys_tmp11500 = (r_run_copy0_j_282 + w_sys_intOne);
	assign w_sys_tmp11501 = (r_run_copy1_j_283 + w_sys_intOne);
	assign w_sys_tmp11502 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp11581 = 32'sh00000061;
	assign w_sys_tmp11582 = ( !w_sys_tmp11583 );
	assign w_sys_tmp11583 = (w_sys_tmp11584 < r_run_k_35);
	assign w_sys_tmp11584 = 32'sh00000080;
	assign w_sys_tmp11585 = (r_run_k_35 + w_sys_intOne);
	assign w_sys_tmp11586 = 32'sh00000002;
	assign w_sys_tmp11587 = ( !w_sys_tmp11588 );
	assign w_sys_tmp11588 = (w_sys_tmp11589 < r_run_j_36);
	assign w_sys_tmp11589 = 32'sh00000010;
	assign w_sys_tmp11592 = (w_sys_tmp11593 + r_run_k_35);
	assign w_sys_tmp11593 = (r_run_j_36 * w_sys_tmp11594);
	assign w_sys_tmp11594 = 32'sh00000081;
	assign w_sys_tmp11595 = w_sub24_result_dataout;
	assign w_sys_tmp11596 = (w_sys_tmp11597 + r_run_k_35);
	assign w_sys_tmp11597 = (r_run_copy0_j_284 * w_sys_tmp11594);
	assign w_sys_tmp11599 = (r_run_copy0_j_284 + w_sys_intOne);
	assign w_sys_tmp11600 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp11661 = 32'sh00000011;
	assign w_sys_tmp11662 = ( !w_sys_tmp11663 );
	assign w_sys_tmp11663 = (w_sys_tmp11664 < r_run_j_36);
	assign w_sys_tmp11664 = 32'sh00000020;
	assign w_sys_tmp11666 = (r_run_j_36 - w_sys_tmp11667);
	assign w_sys_tmp11667 = 32'sh0000000f;
	assign w_sys_tmp11669 = (w_sys_tmp11670 + r_run_k_35);
	assign w_sys_tmp11670 = (r_run_copy1_j_286 * w_sys_tmp11671);
	assign w_sys_tmp11671 = 32'sh00000081;
	assign w_sys_tmp11672 = w_sub25_result_dataout;
	assign w_sys_tmp11673 = (w_sys_tmp11674 + r_run_k_35);
	assign w_sys_tmp11674 = (r_run_copy0_j_285 * w_sys_tmp11671);
	assign w_sys_tmp11676 = (r_run_copy0_j_285 + w_sys_intOne);
	assign w_sys_tmp11677 = (r_run_copy1_j_286 + w_sys_intOne);
	assign w_sys_tmp11678 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp11757 = 32'sh00000021;
	assign w_sys_tmp11758 = ( !w_sys_tmp11759 );
	assign w_sys_tmp11759 = (w_sys_tmp11760 < r_run_j_36);
	assign w_sys_tmp11760 = 32'sh00000030;
	assign w_sys_tmp11762 = (r_run_j_36 - w_sys_tmp11763);
	assign w_sys_tmp11763 = 32'sh0000001f;
	assign w_sys_tmp11765 = (w_sys_tmp11766 + r_run_k_35);
	assign w_sys_tmp11766 = (r_run_copy1_j_288 * w_sys_tmp11767);
	assign w_sys_tmp11767 = 32'sh00000081;
	assign w_sys_tmp11768 = w_sub26_result_dataout;
	assign w_sys_tmp11769 = (w_sys_tmp11770 + r_run_k_35);
	assign w_sys_tmp11770 = (r_run_copy0_j_287 * w_sys_tmp11767);
	assign w_sys_tmp11772 = (r_run_copy0_j_287 + w_sys_intOne);
	assign w_sys_tmp11773 = (r_run_copy1_j_288 + w_sys_intOne);
	assign w_sys_tmp11774 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp11853 = 32'sh00000031;
	assign w_sys_tmp11854 = ( !w_sys_tmp11855 );
	assign w_sys_tmp11855 = (w_sys_tmp11856 < r_run_j_36);
	assign w_sys_tmp11856 = 32'sh00000040;
	assign w_sys_tmp11858 = (r_run_j_36 - w_sys_tmp11859);
	assign w_sys_tmp11859 = 32'sh0000002f;
	assign w_sys_tmp11861 = (w_sys_tmp11862 + r_run_k_35);
	assign w_sys_tmp11862 = (r_run_copy1_j_290 * w_sys_tmp11863);
	assign w_sys_tmp11863 = 32'sh00000081;
	assign w_sys_tmp11864 = w_sub27_result_dataout;
	assign w_sys_tmp11865 = (w_sys_tmp11866 + r_run_k_35);
	assign w_sys_tmp11866 = (r_run_copy0_j_289 * w_sys_tmp11863);
	assign w_sys_tmp11868 = (r_run_copy0_j_289 + w_sys_intOne);
	assign w_sys_tmp11869 = (r_run_copy1_j_290 + w_sys_intOne);
	assign w_sys_tmp11870 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp11949 = 32'sh00000041;
	assign w_sys_tmp11950 = ( !w_sys_tmp11951 );
	assign w_sys_tmp11951 = (w_sys_tmp11952 < r_run_j_36);
	assign w_sys_tmp11952 = 32'sh00000050;
	assign w_sys_tmp11954 = (r_run_j_36 - w_sys_tmp11955);
	assign w_sys_tmp11955 = 32'sh0000003f;
	assign w_sys_tmp11957 = (w_sys_tmp11958 + r_run_k_35);
	assign w_sys_tmp11958 = (r_run_copy1_j_292 * w_sys_tmp11959);
	assign w_sys_tmp11959 = 32'sh00000081;
	assign w_sys_tmp11960 = w_sub28_result_dataout;
	assign w_sys_tmp11961 = (w_sys_tmp11962 + r_run_k_35);
	assign w_sys_tmp11962 = (r_run_copy0_j_291 * w_sys_tmp11959);
	assign w_sys_tmp11964 = (r_run_copy0_j_291 + w_sys_intOne);
	assign w_sys_tmp11965 = (r_run_copy1_j_292 + w_sys_intOne);
	assign w_sys_tmp11966 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp12045 = 32'sh00000051;
	assign w_sys_tmp12046 = ( !w_sys_tmp12047 );
	assign w_sys_tmp12047 = (w_sys_tmp12048 < r_run_j_36);
	assign w_sys_tmp12048 = 32'sh00000060;
	assign w_sys_tmp12050 = (r_run_j_36 - w_sys_tmp12051);
	assign w_sys_tmp12051 = 32'sh0000004f;
	assign w_sys_tmp12053 = (w_sys_tmp12054 + r_run_k_35);
	assign w_sys_tmp12054 = (r_run_copy1_j_294 * w_sys_tmp12055);
	assign w_sys_tmp12055 = 32'sh00000081;
	assign w_sys_tmp12056 = w_sub29_result_dataout;
	assign w_sys_tmp12057 = (w_sys_tmp12058 + r_run_k_35);
	assign w_sys_tmp12058 = (r_run_copy0_j_293 * w_sys_tmp12055);
	assign w_sys_tmp12060 = (r_run_copy0_j_293 + w_sys_intOne);
	assign w_sys_tmp12061 = (r_run_copy1_j_294 + w_sys_intOne);
	assign w_sys_tmp12062 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp12141 = 32'sh00000061;
	assign w_sys_tmp12142 = ( !w_sys_tmp12143 );
	assign w_sys_tmp12143 = (w_sys_tmp12144 < r_run_j_36);
	assign w_sys_tmp12144 = 32'sh00000070;
	assign w_sys_tmp12146 = (r_run_j_36 - w_sys_tmp12147);
	assign w_sys_tmp12147 = 32'sh0000005f;
	assign w_sys_tmp12149 = (w_sys_tmp12150 + r_run_k_35);
	assign w_sys_tmp12150 = (r_run_copy1_j_296 * w_sys_tmp12151);
	assign w_sys_tmp12151 = 32'sh00000081;
	assign w_sys_tmp12152 = w_sub30_result_dataout;
	assign w_sys_tmp12153 = (w_sys_tmp12154 + r_run_k_35);
	assign w_sys_tmp12154 = (r_run_copy0_j_295 * w_sys_tmp12151);
	assign w_sys_tmp12156 = (r_run_copy0_j_295 + w_sys_intOne);
	assign w_sys_tmp12157 = (r_run_copy1_j_296 + w_sys_intOne);
	assign w_sys_tmp12158 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp12237 = 32'sh00000071;
	assign w_sys_tmp12238 = ( !w_sys_tmp12239 );
	assign w_sys_tmp12239 = (w_sys_tmp12240 < r_run_j_36);
	assign w_sys_tmp12240 = 32'sh00000080;
	assign w_sys_tmp12242 = (r_run_j_36 - w_sys_tmp12243);
	assign w_sys_tmp12243 = 32'sh0000006f;
	assign w_sys_tmp12245 = (w_sys_tmp12246 + r_run_k_35);
	assign w_sys_tmp12246 = (r_run_copy1_j_298 * w_sys_tmp12247);
	assign w_sys_tmp12247 = 32'sh00000081;
	assign w_sys_tmp12248 = w_sub31_result_dataout;
	assign w_sys_tmp12249 = (w_sys_tmp12250 + r_run_k_35);
	assign w_sys_tmp12250 = (r_run_copy0_j_297 * w_sys_tmp12247);
	assign w_sys_tmp12252 = (r_run_copy0_j_297 + w_sys_intOne);
	assign w_sys_tmp12253 = (r_run_copy1_j_298 + w_sys_intOne);
	assign w_sys_tmp12254 = (r_run_j_36 + w_sys_intOne);
	assign w_sys_tmp12333 = w_fld_T_0_dataout_1;
	assign w_sys_tmp12334 = 32'sh00000514;


	sub19
		sub19_inst(
			.i_fld_T_0_addr_0 (w_sub19_T_addr),
			.i_fld_T_0_datain_0 (w_sub19_T_datain),
			.o_fld_T_0_dataout_0 (w_sub19_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub19_T_r_w),
			.i_fld_U_1_addr_0 (w_sub19_U_addr),
			.i_fld_U_1_datain_0 (w_sub19_U_datain),
			.o_fld_U_1_dataout_0 (w_sub19_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub19_U_r_w),
			.i_fld_result_2_addr_0 (w_sub19_result_addr),
			.i_fld_result_2_datain_0 (w_sub19_result_datain),
			.o_fld_result_2_dataout_0 (w_sub19_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub19_result_r_w),
			.o_run_busy (w_sub19_run_busy),
			.i_run_req (r_sub19_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub12
		sub12_inst(
			.i_fld_T_0_addr_0 (w_sub12_T_addr),
			.i_fld_T_0_datain_0 (w_sub12_T_datain),
			.o_fld_T_0_dataout_0 (w_sub12_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub12_T_r_w),
			.i_fld_U_1_addr_0 (w_sub12_U_addr),
			.i_fld_U_1_datain_0 (w_sub12_U_datain),
			.o_fld_U_1_dataout_0 (w_sub12_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub12_U_r_w),
			.i_fld_result_2_addr_0 (w_sub12_result_addr),
			.i_fld_result_2_datain_0 (w_sub12_result_datain),
			.o_fld_result_2_dataout_0 (w_sub12_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub12_result_r_w),
			.o_run_busy (w_sub12_run_busy),
			.i_run_req (r_sub12_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub11
		sub11_inst(
			.i_fld_T_0_addr_0 (w_sub11_T_addr),
			.i_fld_T_0_datain_0 (w_sub11_T_datain),
			.o_fld_T_0_dataout_0 (w_sub11_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub11_T_r_w),
			.i_fld_U_2_addr_0 (w_sub11_U_addr),
			.i_fld_U_2_datain_0 (w_sub11_U_datain),
			.o_fld_U_2_dataout_0 (w_sub11_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub11_U_r_w),
			.i_fld_V_1_addr_0 (w_sub11_V_addr),
			.i_fld_V_1_datain_0 (w_sub11_V_datain),
			.o_fld_V_1_dataout_0 (w_sub11_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub11_V_r_w),
			.i_fld_result_3_addr_0 (w_sub11_result_addr),
			.i_fld_result_3_datain_0 (w_sub11_result_datain),
			.o_fld_result_3_dataout_0 (w_sub11_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub11_result_r_w),
			.o_run_busy (w_sub11_run_busy),
			.i_run_req (r_sub11_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub14
		sub14_inst(
			.i_fld_T_0_addr_0 (w_sub14_T_addr),
			.i_fld_T_0_datain_0 (w_sub14_T_datain),
			.o_fld_T_0_dataout_0 (w_sub14_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub14_T_r_w),
			.i_fld_U_1_addr_0 (w_sub14_U_addr),
			.i_fld_U_1_datain_0 (w_sub14_U_datain),
			.o_fld_U_1_dataout_0 (w_sub14_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub14_U_r_w),
			.i_fld_result_2_addr_0 (w_sub14_result_addr),
			.i_fld_result_2_datain_0 (w_sub14_result_datain),
			.o_fld_result_2_dataout_0 (w_sub14_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub14_result_r_w),
			.o_run_busy (w_sub14_run_busy),
			.i_run_req (r_sub14_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub13
		sub13_inst(
			.i_fld_T_0_addr_0 (w_sub13_T_addr),
			.i_fld_T_0_datain_0 (w_sub13_T_datain),
			.o_fld_T_0_dataout_0 (w_sub13_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub13_T_r_w),
			.i_fld_U_1_addr_0 (w_sub13_U_addr),
			.i_fld_U_1_datain_0 (w_sub13_U_datain),
			.o_fld_U_1_dataout_0 (w_sub13_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub13_U_r_w),
			.i_fld_result_2_addr_0 (w_sub13_result_addr),
			.i_fld_result_2_datain_0 (w_sub13_result_datain),
			.o_fld_result_2_dataout_0 (w_sub13_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub13_result_r_w),
			.o_run_busy (w_sub13_run_busy),
			.i_run_req (r_sub13_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub16
		sub16_inst(
			.i_fld_T_0_addr_0 (w_sub16_T_addr),
			.i_fld_T_0_datain_0 (w_sub16_T_datain),
			.o_fld_T_0_dataout_0 (w_sub16_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub16_T_r_w),
			.i_fld_U_1_addr_0 (w_sub16_U_addr),
			.i_fld_U_1_datain_0 (w_sub16_U_datain),
			.o_fld_U_1_dataout_0 (w_sub16_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub16_U_r_w),
			.i_fld_result_2_addr_0 (w_sub16_result_addr),
			.i_fld_result_2_datain_0 (w_sub16_result_datain),
			.o_fld_result_2_dataout_0 (w_sub16_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub16_result_r_w),
			.o_run_busy (w_sub16_run_busy),
			.i_run_req (r_sub16_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub15
		sub15_inst(
			.i_fld_T_0_addr_0 (w_sub15_T_addr),
			.i_fld_T_0_datain_0 (w_sub15_T_datain),
			.o_fld_T_0_dataout_0 (w_sub15_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub15_T_r_w),
			.i_fld_U_1_addr_0 (w_sub15_U_addr),
			.i_fld_U_1_datain_0 (w_sub15_U_datain),
			.o_fld_U_1_dataout_0 (w_sub15_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub15_U_r_w),
			.i_fld_result_2_addr_0 (w_sub15_result_addr),
			.i_fld_result_2_datain_0 (w_sub15_result_datain),
			.o_fld_result_2_dataout_0 (w_sub15_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub15_result_r_w),
			.o_run_busy (w_sub15_run_busy),
			.i_run_req (r_sub15_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub18
		sub18_inst(
			.i_fld_T_0_addr_0 (w_sub18_T_addr),
			.i_fld_T_0_datain_0 (w_sub18_T_datain),
			.o_fld_T_0_dataout_0 (w_sub18_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub18_T_r_w),
			.i_fld_U_1_addr_0 (w_sub18_U_addr),
			.i_fld_U_1_datain_0 (w_sub18_U_datain),
			.o_fld_U_1_dataout_0 (w_sub18_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub18_U_r_w),
			.i_fld_result_2_addr_0 (w_sub18_result_addr),
			.i_fld_result_2_datain_0 (w_sub18_result_datain),
			.o_fld_result_2_dataout_0 (w_sub18_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub18_result_r_w),
			.o_run_busy (w_sub18_run_busy),
			.i_run_req (r_sub18_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub17
		sub17_inst(
			.i_fld_T_0_addr_0 (w_sub17_T_addr),
			.i_fld_T_0_datain_0 (w_sub17_T_datain),
			.o_fld_T_0_dataout_0 (w_sub17_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub17_T_r_w),
			.i_fld_U_1_addr_0 (w_sub17_U_addr),
			.i_fld_U_1_datain_0 (w_sub17_U_datain),
			.o_fld_U_1_dataout_0 (w_sub17_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub17_U_r_w),
			.i_fld_result_2_addr_0 (w_sub17_result_addr),
			.i_fld_result_2_datain_0 (w_sub17_result_datain),
			.o_fld_result_2_dataout_0 (w_sub17_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub17_result_r_w),
			.o_run_busy (w_sub17_run_busy),
			.i_run_req (r_sub17_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub20
		sub20_inst(
			.i_fld_T_0_addr_0 (w_sub20_T_addr),
			.i_fld_T_0_datain_0 (w_sub20_T_datain),
			.o_fld_T_0_dataout_0 (w_sub20_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub20_T_r_w),
			.i_fld_U_1_addr_0 (w_sub20_U_addr),
			.i_fld_U_1_datain_0 (w_sub20_U_datain),
			.o_fld_U_1_dataout_0 (w_sub20_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub20_U_r_w),
			.i_fld_result_2_addr_0 (w_sub20_result_addr),
			.i_fld_result_2_datain_0 (w_sub20_result_datain),
			.o_fld_result_2_dataout_0 (w_sub20_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub20_result_r_w),
			.o_run_busy (w_sub20_run_busy),
			.i_run_req (r_sub20_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub21
		sub21_inst(
			.i_fld_T_0_addr_0 (w_sub21_T_addr),
			.i_fld_T_0_datain_0 (w_sub21_T_datain),
			.o_fld_T_0_dataout_0 (w_sub21_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub21_T_r_w),
			.i_fld_U_1_addr_0 (w_sub21_U_addr),
			.i_fld_U_1_datain_0 (w_sub21_U_datain),
			.o_fld_U_1_dataout_0 (w_sub21_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub21_U_r_w),
			.i_fld_result_2_addr_0 (w_sub21_result_addr),
			.i_fld_result_2_datain_0 (w_sub21_result_datain),
			.o_fld_result_2_dataout_0 (w_sub21_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub21_result_r_w),
			.o_run_busy (w_sub21_run_busy),
			.i_run_req (r_sub21_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub28
		sub28_inst(
			.i_fld_T_0_addr_0 (w_sub28_T_addr),
			.i_fld_T_0_datain_0 (w_sub28_T_datain),
			.o_fld_T_0_dataout_0 (w_sub28_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub28_T_r_w),
			.i_fld_U_1_addr_0 (w_sub28_U_addr),
			.i_fld_U_1_datain_0 (w_sub28_U_datain),
			.o_fld_U_1_dataout_0 (w_sub28_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub28_U_r_w),
			.i_fld_result_2_addr_0 (w_sub28_result_addr),
			.i_fld_result_2_datain_0 (w_sub28_result_datain),
			.o_fld_result_2_dataout_0 (w_sub28_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub28_result_r_w),
			.o_run_busy (w_sub28_run_busy),
			.i_run_req (r_sub28_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub29
		sub29_inst(
			.i_fld_T_0_addr_0 (w_sub29_T_addr),
			.i_fld_T_0_datain_0 (w_sub29_T_datain),
			.o_fld_T_0_dataout_0 (w_sub29_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub29_T_r_w),
			.i_fld_U_1_addr_0 (w_sub29_U_addr),
			.i_fld_U_1_datain_0 (w_sub29_U_datain),
			.o_fld_U_1_dataout_0 (w_sub29_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub29_U_r_w),
			.i_fld_result_2_addr_0 (w_sub29_result_addr),
			.i_fld_result_2_datain_0 (w_sub29_result_datain),
			.o_fld_result_2_dataout_0 (w_sub29_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub29_result_r_w),
			.o_run_busy (w_sub29_run_busy),
			.i_run_req (r_sub29_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub26
		sub26_inst(
			.i_fld_T_0_addr_0 (w_sub26_T_addr),
			.i_fld_T_0_datain_0 (w_sub26_T_datain),
			.o_fld_T_0_dataout_0 (w_sub26_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub26_T_r_w),
			.i_fld_U_1_addr_0 (w_sub26_U_addr),
			.i_fld_U_1_datain_0 (w_sub26_U_datain),
			.o_fld_U_1_dataout_0 (w_sub26_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub26_U_r_w),
			.i_fld_result_2_addr_0 (w_sub26_result_addr),
			.i_fld_result_2_datain_0 (w_sub26_result_datain),
			.o_fld_result_2_dataout_0 (w_sub26_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub26_result_r_w),
			.o_run_busy (w_sub26_run_busy),
			.i_run_req (r_sub26_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub09
		sub09_inst(
			.i_fld_T_0_addr_0 (w_sub09_T_addr),
			.i_fld_T_0_datain_0 (w_sub09_T_datain),
			.o_fld_T_0_dataout_0 (w_sub09_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub09_T_r_w),
			.i_fld_U_1_addr_0 (w_sub09_U_addr),
			.i_fld_U_1_datain_0 (w_sub09_U_datain),
			.o_fld_U_1_dataout_0 (w_sub09_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub09_U_r_w),
			.i_fld_result_2_addr_0 (w_sub09_result_addr),
			.i_fld_result_2_datain_0 (w_sub09_result_datain),
			.o_fld_result_2_dataout_0 (w_sub09_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub09_result_r_w),
			.o_run_busy (w_sub09_run_busy),
			.i_run_req (r_sub09_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub27
		sub27_inst(
			.i_fld_T_0_addr_0 (w_sub27_T_addr),
			.i_fld_T_0_datain_0 (w_sub27_T_datain),
			.o_fld_T_0_dataout_0 (w_sub27_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub27_T_r_w),
			.i_fld_U_1_addr_0 (w_sub27_U_addr),
			.i_fld_U_1_datain_0 (w_sub27_U_datain),
			.o_fld_U_1_dataout_0 (w_sub27_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub27_U_r_w),
			.i_fld_result_2_addr_0 (w_sub27_result_addr),
			.i_fld_result_2_datain_0 (w_sub27_result_datain),
			.o_fld_result_2_dataout_0 (w_sub27_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub27_result_r_w),
			.o_run_busy (w_sub27_run_busy),
			.i_run_req (r_sub27_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub08
		sub08_inst(
			.i_fld_T_0_addr_0 (w_sub08_T_addr),
			.i_fld_T_0_datain_0 (w_sub08_T_datain),
			.o_fld_T_0_dataout_0 (w_sub08_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub08_T_r_w),
			.i_fld_U_1_addr_0 (w_sub08_U_addr),
			.i_fld_U_1_datain_0 (w_sub08_U_datain),
			.o_fld_U_1_dataout_0 (w_sub08_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub08_U_r_w),
			.i_fld_result_2_addr_0 (w_sub08_result_addr),
			.i_fld_result_2_datain_0 (w_sub08_result_datain),
			.o_fld_result_2_dataout_0 (w_sub08_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub08_result_r_w),
			.o_run_busy (w_sub08_run_busy),
			.i_run_req (r_sub08_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub24
		sub24_inst(
			.i_fld_T_0_addr_0 (w_sub24_T_addr),
			.i_fld_T_0_datain_0 (w_sub24_T_datain),
			.o_fld_T_0_dataout_0 (w_sub24_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub24_T_r_w),
			.i_fld_U_1_addr_0 (w_sub24_U_addr),
			.i_fld_U_1_datain_0 (w_sub24_U_datain),
			.o_fld_U_1_dataout_0 (w_sub24_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub24_U_r_w),
			.i_fld_result_2_addr_0 (w_sub24_result_addr),
			.i_fld_result_2_datain_0 (w_sub24_result_datain),
			.o_fld_result_2_dataout_0 (w_sub24_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub24_result_r_w),
			.o_run_busy (w_sub24_run_busy),
			.i_run_req (r_sub24_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub25
		sub25_inst(
			.i_fld_T_0_addr_0 (w_sub25_T_addr),
			.i_fld_T_0_datain_0 (w_sub25_T_datain),
			.o_fld_T_0_dataout_0 (w_sub25_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub25_T_r_w),
			.i_fld_U_1_addr_0 (w_sub25_U_addr),
			.i_fld_U_1_datain_0 (w_sub25_U_datain),
			.o_fld_U_1_dataout_0 (w_sub25_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub25_U_r_w),
			.i_fld_result_2_addr_0 (w_sub25_result_addr),
			.i_fld_result_2_datain_0 (w_sub25_result_datain),
			.o_fld_result_2_dataout_0 (w_sub25_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub25_result_r_w),
			.o_run_busy (w_sub25_run_busy),
			.i_run_req (r_sub25_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub22
		sub22_inst(
			.i_fld_T_0_addr_0 (w_sub22_T_addr),
			.i_fld_T_0_datain_0 (w_sub22_T_datain),
			.o_fld_T_0_dataout_0 (w_sub22_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub22_T_r_w),
			.i_fld_U_1_addr_0 (w_sub22_U_addr),
			.i_fld_U_1_datain_0 (w_sub22_U_datain),
			.o_fld_U_1_dataout_0 (w_sub22_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub22_U_r_w),
			.i_fld_result_2_addr_0 (w_sub22_result_addr),
			.i_fld_result_2_datain_0 (w_sub22_result_datain),
			.o_fld_result_2_dataout_0 (w_sub22_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub22_result_r_w),
			.o_run_busy (w_sub22_run_busy),
			.i_run_req (r_sub22_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub23
		sub23_inst(
			.i_fld_T_0_addr_0 (w_sub23_T_addr),
			.i_fld_T_0_datain_0 (w_sub23_T_datain),
			.o_fld_T_0_dataout_0 (w_sub23_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub23_T_r_w),
			.i_fld_U_1_addr_0 (w_sub23_U_addr),
			.i_fld_U_1_datain_0 (w_sub23_U_datain),
			.o_fld_U_1_dataout_0 (w_sub23_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub23_U_r_w),
			.i_fld_result_2_addr_0 (w_sub23_result_addr),
			.i_fld_result_2_datain_0 (w_sub23_result_datain),
			.o_fld_result_2_dataout_0 (w_sub23_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub23_result_r_w),
			.o_run_busy (w_sub23_run_busy),
			.i_run_req (r_sub23_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub03
		sub03_inst(
			.i_fld_T_0_addr_0 (w_sub03_T_addr),
			.i_fld_T_0_datain_0 (w_sub03_T_datain),
			.o_fld_T_0_dataout_0 (w_sub03_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub03_T_r_w),
			.i_fld_U_1_addr_0 (w_sub03_U_addr),
			.i_fld_U_1_datain_0 (w_sub03_U_datain),
			.o_fld_U_1_dataout_0 (w_sub03_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub03_U_r_w),
			.i_fld_result_2_addr_0 (w_sub03_result_addr),
			.i_fld_result_2_datain_0 (w_sub03_result_datain),
			.o_fld_result_2_dataout_0 (w_sub03_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub03_result_r_w),
			.o_run_busy (w_sub03_run_busy),
			.i_run_req (r_sub03_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub02
		sub02_inst(
			.i_fld_T_0_addr_0 (w_sub02_T_addr),
			.i_fld_T_0_datain_0 (w_sub02_T_datain),
			.o_fld_T_0_dataout_0 (w_sub02_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub02_T_r_w),
			.i_fld_U_1_addr_0 (w_sub02_U_addr),
			.i_fld_U_1_datain_0 (w_sub02_U_datain),
			.o_fld_U_1_dataout_0 (w_sub02_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub02_U_r_w),
			.i_fld_result_2_addr_0 (w_sub02_result_addr),
			.i_fld_result_2_datain_0 (w_sub02_result_datain),
			.o_fld_result_2_dataout_0 (w_sub02_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub02_result_r_w),
			.o_run_busy (w_sub02_run_busy),
			.i_run_req (r_sub02_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub01
		sub01_inst(
			.i_fld_T_0_addr_0 (w_sub01_T_addr),
			.i_fld_T_0_datain_0 (w_sub01_T_datain),
			.o_fld_T_0_dataout_0 (w_sub01_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub01_T_r_w),
			.i_fld_U_1_addr_0 (w_sub01_U_addr),
			.i_fld_U_1_datain_0 (w_sub01_U_datain),
			.o_fld_U_1_dataout_0 (w_sub01_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub01_U_r_w),
			.i_fld_result_2_addr_0 (w_sub01_result_addr),
			.i_fld_result_2_datain_0 (w_sub01_result_datain),
			.o_fld_result_2_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub01_result_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub00
		sub00_inst(
			.i_fld_T_0_addr_0 (w_sub00_T_addr),
			.i_fld_T_0_datain_0 (w_sub00_T_datain),
			.o_fld_T_0_dataout_0 (w_sub00_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub00_T_r_w),
			.i_fld_U_1_addr_0 (w_sub00_U_addr),
			.i_fld_U_1_datain_0 (w_sub00_U_datain),
			.o_fld_U_1_dataout_0 (w_sub00_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub00_U_r_w),
			.i_fld_result_2_addr_0 (w_sub00_result_addr),
			.i_fld_result_2_datain_0 (w_sub00_result_datain),
			.o_fld_result_2_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub00_result_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub07
		sub07_inst(
			.i_fld_T_0_addr_0 (w_sub07_T_addr),
			.i_fld_T_0_datain_0 (w_sub07_T_datain),
			.o_fld_T_0_dataout_0 (w_sub07_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub07_T_r_w),
			.i_fld_U_1_addr_0 (w_sub07_U_addr),
			.i_fld_U_1_datain_0 (w_sub07_U_datain),
			.o_fld_U_1_dataout_0 (w_sub07_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub07_U_r_w),
			.i_fld_result_2_addr_0 (w_sub07_result_addr),
			.i_fld_result_2_datain_0 (w_sub07_result_datain),
			.o_fld_result_2_dataout_0 (w_sub07_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub07_result_r_w),
			.o_run_busy (w_sub07_run_busy),
			.i_run_req (r_sub07_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub06
		sub06_inst(
			.i_fld_T_0_addr_0 (w_sub06_T_addr),
			.i_fld_T_0_datain_0 (w_sub06_T_datain),
			.o_fld_T_0_dataout_0 (w_sub06_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub06_T_r_w),
			.i_fld_U_1_addr_0 (w_sub06_U_addr),
			.i_fld_U_1_datain_0 (w_sub06_U_datain),
			.o_fld_U_1_dataout_0 (w_sub06_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub06_U_r_w),
			.i_fld_result_2_addr_0 (w_sub06_result_addr),
			.i_fld_result_2_datain_0 (w_sub06_result_datain),
			.o_fld_result_2_dataout_0 (w_sub06_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub06_result_r_w),
			.o_run_busy (w_sub06_run_busy),
			.i_run_req (r_sub06_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub05
		sub05_inst(
			.i_fld_T_0_addr_0 (w_sub05_T_addr),
			.i_fld_T_0_datain_0 (w_sub05_T_datain),
			.o_fld_T_0_dataout_0 (w_sub05_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub05_T_r_w),
			.i_fld_U_1_addr_0 (w_sub05_U_addr),
			.i_fld_U_1_datain_0 (w_sub05_U_datain),
			.o_fld_U_1_dataout_0 (w_sub05_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub05_U_r_w),
			.i_fld_result_2_addr_0 (w_sub05_result_addr),
			.i_fld_result_2_datain_0 (w_sub05_result_datain),
			.o_fld_result_2_dataout_0 (w_sub05_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub05_result_r_w),
			.o_run_busy (w_sub05_run_busy),
			.i_run_req (r_sub05_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub04
		sub04_inst(
			.i_fld_T_0_addr_0 (w_sub04_T_addr),
			.i_fld_T_0_datain_0 (w_sub04_T_datain),
			.o_fld_T_0_dataout_0 (w_sub04_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub04_T_r_w),
			.i_fld_U_1_addr_0 (w_sub04_U_addr),
			.i_fld_U_1_datain_0 (w_sub04_U_datain),
			.o_fld_U_1_dataout_0 (w_sub04_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub04_U_r_w),
			.i_fld_result_2_addr_0 (w_sub04_result_addr),
			.i_fld_result_2_datain_0 (w_sub04_result_datain),
			.o_fld_result_2_dataout_0 (w_sub04_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub04_result_r_w),
			.o_run_busy (w_sub04_run_busy),
			.i_run_req (r_sub04_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub10
		sub10_inst(
			.i_fld_T_0_addr_0 (w_sub10_T_addr),
			.i_fld_T_0_datain_0 (w_sub10_T_datain),
			.o_fld_T_0_dataout_0 (w_sub10_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub10_T_r_w),
			.i_fld_U_1_addr_0 (w_sub10_U_addr),
			.i_fld_U_1_datain_0 (w_sub10_U_datain),
			.o_fld_U_1_dataout_0 (w_sub10_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub10_U_r_w),
			.i_fld_result_2_addr_0 (w_sub10_result_addr),
			.i_fld_result_2_datain_0 (w_sub10_result_datain),
			.o_fld_result_2_dataout_0 (w_sub10_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub10_result_r_w),
			.o_run_busy (w_sub10_run_busy),
			.i_run_req (r_sub10_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub31
		sub31_inst(
			.i_fld_T_0_addr_0 (w_sub31_T_addr),
			.i_fld_T_0_datain_0 (w_sub31_T_datain),
			.o_fld_T_0_dataout_0 (w_sub31_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub31_T_r_w),
			.i_fld_U_1_addr_0 (w_sub31_U_addr),
			.i_fld_U_1_datain_0 (w_sub31_U_datain),
			.o_fld_U_1_dataout_0 (w_sub31_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub31_U_r_w),
			.i_fld_result_2_addr_0 (w_sub31_result_addr),
			.i_fld_result_2_datain_0 (w_sub31_result_datain),
			.o_fld_result_2_dataout_0 (w_sub31_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub31_result_r_w),
			.o_run_busy (w_sub31_run_busy),
			.i_run_req (r_sub31_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub30
		sub30_inst(
			.i_fld_T_0_addr_0 (w_sub30_T_addr),
			.i_fld_T_0_datain_0 (w_sub30_T_datain),
			.o_fld_T_0_dataout_0 (w_sub30_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub30_T_r_w),
			.i_fld_U_1_addr_0 (w_sub30_U_addr),
			.i_fld_U_1_datain_0 (w_sub30_U_datain),
			.o_fld_U_1_dataout_0 (w_sub30_U_dataout),
			.i_fld_U_1_r_w_0 (w_sub30_U_r_w),
			.i_fld_result_2_addr_0 (w_sub30_result_addr),
			.i_fld_result_2_datain_0 (w_sub30_result_datain),
			.o_fld_result_2_dataout_0 (w_sub30_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub30_result_r_w),
			.o_run_busy (w_sub30_run_busy),
			.i_run_req (r_sub30_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_T_0(
			.clk (clock),
			.ce_0 (w_fld_T_0_ce_0),
			.addr_0 (w_fld_T_0_addr_0),
			.datain_0 (w_fld_T_0_datain_0),
			.dataout_0 (w_fld_T_0_dataout_0),
			.r_w_0 (w_fld_T_0_r_w_0),
			.ce_1 (w_fld_T_0_ce_1),
			.addr_1 (r_fld_T_0_addr_1),
			.datain_1 (r_fld_T_0_datain_1),
			.dataout_1 (w_fld_T_0_dataout_1),
			.r_w_1 (r_fld_T_0_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_TT_1(
			.clk (clock),
			.ce_0 (w_fld_TT_1_ce_0),
			.addr_0 (w_fld_TT_1_addr_0),
			.datain_0 (w_fld_TT_1_datain_0),
			.dataout_0 (w_fld_TT_1_dataout_0),
			.r_w_0 (w_fld_TT_1_r_w_0),
			.ce_1 (w_fld_TT_1_ce_1),
			.addr_1 (r_fld_TT_1_addr_1),
			.datain_1 (r_fld_TT_1_datain_1),
			.dataout_1 (w_fld_TT_1_dataout_1),
			.r_w_1 (r_fld_TT_1_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_U_2(
			.clk (clock),
			.ce_0 (w_fld_U_2_ce_0),
			.addr_0 (w_fld_U_2_addr_0),
			.datain_0 (w_fld_U_2_datain_0),
			.dataout_0 (w_fld_U_2_dataout_0),
			.r_w_0 (w_fld_U_2_r_w_0),
			.ce_1 (w_fld_U_2_ce_1),
			.addr_1 (r_fld_U_2_addr_1),
			.datain_1 (r_fld_U_2_datain_1),
			.dataout_1 (w_fld_U_2_dataout_1),
			.r_w_1 (r_fld_U_2_r_w_1)
		);

	AddFloat
		AddFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_AddFloat_portA_0),
			.b (r_ip_AddFloat_portB_0),
			.result (w_ip_AddFloat_result_0)
		);

	MultFloat
		MultFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_MultFloat_multiplicand_0),
			.b (r_ip_MultFloat_multiplier_0),
			.result (w_ip_MultFloat_product_0)
		);

	FixedToFloat
		FixedToFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_FixedToFloat_fixed_0),
			.result (w_ip_FixedToFloat_floating_0)
		);

	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hc) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h14)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp38;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'he)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
									else
									if((r_sys_run_step==6'h14)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
									else
									if((r_sys_run_step==6'h10)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp110[31], w_sys_tmp110[30:0] };

									end
									else
									if((r_sys_run_step==6'h12)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
									else
									if((r_sys_run_step==6'hc)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
									else
									if((r_sys_run_step==6'h11)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp110[31], w_sys_tmp110[30:0] };

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h13) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp4_float;

									end
									else
									if((6'h7<=r_sys_run_step && r_sys_run_step<=6'hb) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'hf)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_dy_42;

									end
									else
									if((r_sys_run_step==6'h18)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h1b)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp18;

									end
									else
									if((r_sys_run_step==6'hc) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h16)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp36;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'hf)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'h15) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1b)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==6'h19)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp1_float;

									end
									else
									if((6'h7<=r_sys_run_step && r_sys_run_step<=6'hb)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp19;

									end
									else
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h16)) begin
										r_ip_MultFloat_multiplier_0 <= r_run_YY_47;

									end
									else
									if((r_sys_run_step==6'hc)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp37;

									end
									else
									if((r_sys_run_step==6'h13) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1a)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp3_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_ip_FixedToFloat_fixed_0 <= w_sys_tmp20;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						10'h21b: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_return <= 32'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h218: begin
							r_sys_run_return <= r_sys_tmp6_float;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 10'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h0: begin
							r_sys_run_phase <= 10'h2;
						end

						10'h2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h4;

									end
								end

							endcase
						end

						10'h4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h5;

									end
								end

							endcase
						end

						10'h5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp12) ? 10'h9 : 10'hf);

									end
								end

							endcase
						end

						10'h6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h5;

									end
								end

							endcase
						end

						10'h9: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'ha;

									end
								end

							endcase
						end

						10'ha: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp15) ? 10'hd : 10'h6);

									end
								end

							endcase
						end

						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h20)) begin
										r_sys_run_phase <= 10'ha;

									end
								end

							endcase
						end

						10'hf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h10;

									end
								end

							endcase
						end

						10'h10: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp184) ? 10'h13 : 10'h15);

									end
								end

							endcase
						end

						10'h13: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_run_phase <= 10'h10;

									end
								end

							endcase
						end

						10'h15: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h16;

									end
								end

							endcase
						end

						10'h16: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp202) ? 10'h19 : 10'h1b);

									end
								end

							endcase
						end

						10'h19: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_phase <= 10'h16;

									end
								end

							endcase
						end

						10'h1b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1c;

									end
								end

							endcase
						end

						10'h1c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp292) ? 10'h1f : 10'h21);

									end
								end

							endcase
						end

						10'h1f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sys_run_phase <= 10'h1c;

									end
								end

							endcase
						end

						10'h21: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h22;

									end
								end

							endcase
						end

						10'h22: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp339) ? 10'h26 : 10'h56);

									end
								end

							endcase
						end

						10'h23: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h22;

									end
								end

							endcase
						end

						10'h26: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h27;

									end
								end

							endcase
						end

						10'h27: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp343) ? 10'h2a : 10'h2c);

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h27;

									end
								end

							endcase
						end

						10'h2c: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h2d;

									end
								end

							endcase
						end

						10'h2d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp488) ? 10'h30 : 10'h32);

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h2d;

									end
								end

							endcase
						end

						10'h32: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h33;

									end
								end

							endcase
						end

						10'h33: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp633) ? 10'h36 : 10'h38);

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h33;

									end
								end

							endcase
						end

						10'h38: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h39;

									end
								end

							endcase
						end

						10'h39: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp778) ? 10'h3c : 10'h3e);

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h39;

									end
								end

							endcase
						end

						10'h3e: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h3f;

									end
								end

							endcase
						end

						10'h3f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp923) ? 10'h42 : 10'h44);

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h3f;

									end
								end

							endcase
						end

						10'h44: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h45;

									end
								end

							endcase
						end

						10'h45: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1068) ? 10'h48 : 10'h4a);

									end
								end

							endcase
						end

						10'h48: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h45;

									end
								end

							endcase
						end

						10'h4a: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h4b;

									end
								end

							endcase
						end

						10'h4b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1213) ? 10'h4e : 10'h50);

									end
								end

							endcase
						end

						10'h4e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h4b;

									end
								end

							endcase
						end

						10'h50: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h51;

									end
								end

							endcase
						end

						10'h51: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1358) ? 10'h54 : 10'h23);

									end
								end

							endcase
						end

						10'h54: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h51;

									end
								end

							endcase
						end

						10'h56: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h57;

									end
								end

							endcase
						end

						10'h57: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1502) ? 10'h5b : 10'h8b);

									end
								end

							endcase
						end

						10'h58: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h57;

									end
								end

							endcase
						end

						10'h5b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h5c;

									end
								end

							endcase
						end

						10'h5c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1506) ? 10'h5f : 10'h61);

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h5c;

									end
								end

							endcase
						end

						10'h61: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h62;

									end
								end

							endcase
						end

						10'h62: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1651) ? 10'h65 : 10'h67);

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h62;

									end
								end

							endcase
						end

						10'h67: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h68;

									end
								end

							endcase
						end

						10'h68: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1796) ? 10'h6b : 10'h6d);

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h68;

									end
								end

							endcase
						end

						10'h6d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h6e;

									end
								end

							endcase
						end

						10'h6e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1941) ? 10'h71 : 10'h73);

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h6e;

									end
								end

							endcase
						end

						10'h73: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h74;

									end
								end

							endcase
						end

						10'h74: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2086) ? 10'h77 : 10'h79);

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h74;

									end
								end

							endcase
						end

						10'h79: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h7a;

									end
								end

							endcase
						end

						10'h7a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2231) ? 10'h7d : 10'h7f);

									end
								end

							endcase
						end

						10'h7d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h7a;

									end
								end

							endcase
						end

						10'h7f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h80;

									end
								end

							endcase
						end

						10'h80: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2376) ? 10'h83 : 10'h85);

									end
								end

							endcase
						end

						10'h83: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h80;

									end
								end

							endcase
						end

						10'h85: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h86;

									end
								end

							endcase
						end

						10'h86: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2521) ? 10'h89 : 10'h58);

									end
								end

							endcase
						end

						10'h89: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h86;

									end
								end

							endcase
						end

						10'h8b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h8c;

									end
								end

							endcase
						end

						10'h8c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2665) ? 10'h90 : 10'hc0);

									end
								end

							endcase
						end

						10'h8d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h8c;

									end
								end

							endcase
						end

						10'h90: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h91;

									end
								end

							endcase
						end

						10'h91: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2669) ? 10'h94 : 10'h96);

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h91;

									end
								end

							endcase
						end

						10'h96: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h97;

									end
								end

							endcase
						end

						10'h97: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2814) ? 10'h9a : 10'h9c);

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h97;

									end
								end

							endcase
						end

						10'h9c: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h9d;

									end
								end

							endcase
						end

						10'h9d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2959) ? 10'ha0 : 10'ha2);

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h9d;

									end
								end

							endcase
						end

						10'ha2: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'ha3;

									end
								end

							endcase
						end

						10'ha3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3104) ? 10'ha6 : 10'ha8);

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'ha3;

									end
								end

							endcase
						end

						10'ha8: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'ha9;

									end
								end

							endcase
						end

						10'ha9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3249) ? 10'hac : 10'hae);

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'ha9;

									end
								end

							endcase
						end

						10'hae: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'haf;

									end
								end

							endcase
						end

						10'haf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3394) ? 10'hb2 : 10'hb4);

									end
								end

							endcase
						end

						10'hb2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'haf;

									end
								end

							endcase
						end

						10'hb4: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hb5;

									end
								end

							endcase
						end

						10'hb5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3539) ? 10'hb8 : 10'hba);

									end
								end

							endcase
						end

						10'hb8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'hb5;

									end
								end

							endcase
						end

						10'hba: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hbb;

									end
								end

							endcase
						end

						10'hbb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3684) ? 10'hbe : 10'h8d);

									end
								end

							endcase
						end

						10'hbe: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'hbb;

									end
								end

							endcase
						end

						10'hc0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hc1;

									end
								end

							endcase
						end

						10'hc1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3828) ? 10'hc5 : 10'hf5);

									end
								end

							endcase
						end

						10'hc2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hc1;

									end
								end

							endcase
						end

						10'hc5: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hc6;

									end
								end

							endcase
						end

						10'hc6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3832) ? 10'hc9 : 10'hcb);

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'hc6;

									end
								end

							endcase
						end

						10'hcb: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hcc;

									end
								end

							endcase
						end

						10'hcc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3977) ? 10'hcf : 10'hd1);

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'hcc;

									end
								end

							endcase
						end

						10'hd1: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hd2;

									end
								end

							endcase
						end

						10'hd2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4122) ? 10'hd5 : 10'hd7);

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'hd2;

									end
								end

							endcase
						end

						10'hd7: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hd8;

									end
								end

							endcase
						end

						10'hd8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4267) ? 10'hdb : 10'hdd);

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'hd8;

									end
								end

							endcase
						end

						10'hdd: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hde;

									end
								end

							endcase
						end

						10'hde: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4412) ? 10'he1 : 10'he3);

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'hde;

									end
								end

							endcase
						end

						10'he3: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'he4;

									end
								end

							endcase
						end

						10'he4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4557) ? 10'he7 : 10'he9);

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'he4;

									end
								end

							endcase
						end

						10'he9: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hea;

									end
								end

							endcase
						end

						10'hea: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4702) ? 10'hed : 10'hef);

									end
								end

							endcase
						end

						10'hed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'hea;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hf0;

									end
								end

							endcase
						end

						10'hf0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4847) ? 10'hf3 : 10'hc2);

									end
								end

							endcase
						end

						10'hf3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'hf0;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hf6;

									end
								end

							endcase
						end

						10'hf6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4991) ? 10'hf9 : 10'h145);

									end
								end

							endcase
						end

						10'hf7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hf6;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h1e: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_phase <= 10'hfb;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								6'h1f: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_phase <= 10'hfd;

									end
								end

							endcase
						end

						10'hfd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hfe;

									end
								end

							endcase
						end

						10'hfe: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4995) ? 10'h101 : 10'h103);

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_phase <= 10'hfe;

									end
								end

							endcase
						end

						10'h103: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h104;

									end
								end

							endcase
						end

						10'h104: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp5079) ? 10'h107 : 10'h109);

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_phase <= 10'h104;

									end
								end

							endcase
						end

						10'h109: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h10a;

									end
								end

							endcase
						end

						10'h10a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp5163) ? 10'h10d : 10'h10f);

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_phase <= 10'h10a;

									end
								end

							endcase
						end

						10'h10f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h110;

									end
								end

							endcase
						end

						10'h110: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp5247) ? 10'h113 : 10'h115);

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_phase <= 10'h110;

									end
								end

							endcase
						end

						10'h115: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h116;

									end
								end

							endcase
						end

						10'h116: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp5330) ? 10'h119 : 10'h11b);

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 10'h116;

									end
								end

							endcase
						end

						10'h11b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h11c;

									end
								end

							endcase
						end

						10'h11c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp5831) ? 10'h11f : 10'h121);

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 10'h11c;

									end
								end

							endcase
						end

						10'h121: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h122;

									end
								end

							endcase
						end

						10'h122: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6332) ? 10'h125 : 10'h127);

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 10'h122;

									end
								end

							endcase
						end

						10'h127: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h128;

									end
								end

							endcase
						end

						10'h128: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6833) ? 10'h12b : 10'h12d);

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 10'h128;

									end
								end

							endcase
						end

						10'h12d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h12e;

									end
								end

							endcase
						end

						10'h12e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7334) ? 10'h131 : 10'h133);

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 10'h12e;

									end
								end

							endcase
						end

						10'h133: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h134;

									end
								end

							endcase
						end

						10'h134: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7835) ? 10'h137 : 10'h139);

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 10'h134;

									end
								end

							endcase
						end

						10'h139: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h13a;

									end
								end

							endcase
						end

						10'h13a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp8336) ? 10'h13d : 10'h13f);

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 10'h13a;

									end
								end

							endcase
						end

						10'h13f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h140;

									end
								end

							endcase
						end

						10'h140: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp8837) ? 10'h143 : 10'hf7);

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3a)) begin
										r_sys_run_phase <= 10'h140;

									end
								end

							endcase
						end

						10'h145: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h146;

									end
								end

							endcase
						end

						10'h146: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp9326) ? 10'h14a : 10'h17a);

									end
								end

							endcase
						end

						10'h147: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h146;

									end
								end

							endcase
						end

						10'h14a: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h14b;

									end
								end

							endcase
						end

						10'h14b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp9331) ? 10'h14e : 10'h150);

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h14b;

									end
								end

							endcase
						end

						10'h150: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h151;

									end
								end

							endcase
						end

						10'h151: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp9406) ? 10'h154 : 10'h156);

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h151;

									end
								end

							endcase
						end

						10'h156: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h157;

									end
								end

							endcase
						end

						10'h157: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp9502) ? 10'h15a : 10'h15c);

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h157;

									end
								end

							endcase
						end

						10'h15c: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h15d;

									end
								end

							endcase
						end

						10'h15d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp9598) ? 10'h160 : 10'h162);

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h15d;

									end
								end

							endcase
						end

						10'h162: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h163;

									end
								end

							endcase
						end

						10'h163: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp9694) ? 10'h166 : 10'h168);

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h163;

									end
								end

							endcase
						end

						10'h168: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h169;

									end
								end

							endcase
						end

						10'h169: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp9790) ? 10'h16c : 10'h16e);

									end
								end

							endcase
						end

						10'h16c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h169;

									end
								end

							endcase
						end

						10'h16e: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h16f;

									end
								end

							endcase
						end

						10'h16f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp9886) ? 10'h172 : 10'h174);

									end
								end

							endcase
						end

						10'h172: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h16f;

									end
								end

							endcase
						end

						10'h174: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h175;

									end
								end

							endcase
						end

						10'h175: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp9982) ? 10'h178 : 10'h147);

									end
								end

							endcase
						end

						10'h178: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h175;

									end
								end

							endcase
						end

						10'h17a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h17b;

									end
								end

							endcase
						end

						10'h17b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp10078) ? 10'h17f : 10'h1af);

									end
								end

							endcase
						end

						10'h17c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h17b;

									end
								end

							endcase
						end

						10'h17f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h180;

									end
								end

							endcase
						end

						10'h180: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp10083) ? 10'h183 : 10'h185);

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h180;

									end
								end

							endcase
						end

						10'h185: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h186;

									end
								end

							endcase
						end

						10'h186: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp10158) ? 10'h189 : 10'h18b);

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h186;

									end
								end

							endcase
						end

						10'h18b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h18c;

									end
								end

							endcase
						end

						10'h18c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp10254) ? 10'h18f : 10'h191);

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h18c;

									end
								end

							endcase
						end

						10'h191: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h192;

									end
								end

							endcase
						end

						10'h192: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp10350) ? 10'h195 : 10'h197);

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h192;

									end
								end

							endcase
						end

						10'h197: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h198;

									end
								end

							endcase
						end

						10'h198: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp10446) ? 10'h19b : 10'h19d);

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h198;

									end
								end

							endcase
						end

						10'h19d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h19e;

									end
								end

							endcase
						end

						10'h19e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp10542) ? 10'h1a1 : 10'h1a3);

									end
								end

							endcase
						end

						10'h1a1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h19e;

									end
								end

							endcase
						end

						10'h1a3: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1a4;

									end
								end

							endcase
						end

						10'h1a4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp10638) ? 10'h1a7 : 10'h1a9);

									end
								end

							endcase
						end

						10'h1a7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1a4;

									end
								end

							endcase
						end

						10'h1a9: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1aa;

									end
								end

							endcase
						end

						10'h1aa: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp10734) ? 10'h1ad : 10'h17c);

									end
								end

							endcase
						end

						10'h1ad: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1aa;

									end
								end

							endcase
						end

						10'h1af: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1b0;

									end
								end

							endcase
						end

						10'h1b0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp10830) ? 10'h1b4 : 10'h1e4);

									end
								end

							endcase
						end

						10'h1b1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1b0;

									end
								end

							endcase
						end

						10'h1b4: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1b5;

									end
								end

							endcase
						end

						10'h1b5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp10835) ? 10'h1b8 : 10'h1ba);

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1b5;

									end
								end

							endcase
						end

						10'h1ba: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1bb;

									end
								end

							endcase
						end

						10'h1bb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp10910) ? 10'h1be : 10'h1c0);

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1bb;

									end
								end

							endcase
						end

						10'h1c0: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1c1;

									end
								end

							endcase
						end

						10'h1c1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp11006) ? 10'h1c4 : 10'h1c6);

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1c1;

									end
								end

							endcase
						end

						10'h1c6: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1c7;

									end
								end

							endcase
						end

						10'h1c7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp11102) ? 10'h1ca : 10'h1cc);

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1c7;

									end
								end

							endcase
						end

						10'h1cc: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1cd;

									end
								end

							endcase
						end

						10'h1cd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp11198) ? 10'h1d0 : 10'h1d2);

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1cd;

									end
								end

							endcase
						end

						10'h1d2: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1d3;

									end
								end

							endcase
						end

						10'h1d3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp11294) ? 10'h1d6 : 10'h1d8);

									end
								end

							endcase
						end

						10'h1d6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1d3;

									end
								end

							endcase
						end

						10'h1d8: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1d9;

									end
								end

							endcase
						end

						10'h1d9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp11390) ? 10'h1dc : 10'h1de);

									end
								end

							endcase
						end

						10'h1dc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1d9;

									end
								end

							endcase
						end

						10'h1de: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1df;

									end
								end

							endcase
						end

						10'h1df: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp11486) ? 10'h1e2 : 10'h1b1);

									end
								end

							endcase
						end

						10'h1e2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1df;

									end
								end

							endcase
						end

						10'h1e4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1e5;

									end
								end

							endcase
						end

						10'h1e5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp11582) ? 10'h1e9 : 10'h219);

									end
								end

							endcase
						end

						10'h1e6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1e5;

									end
								end

							endcase
						end

						10'h1e9: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1ea;

									end
								end

							endcase
						end

						10'h1ea: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp11587) ? 10'h1ed : 10'h1ef);

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1ea;

									end
								end

							endcase
						end

						10'h1ef: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1f0;

									end
								end

							endcase
						end

						10'h1f0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp11662) ? 10'h1f3 : 10'h1f5);

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1f0;

									end
								end

							endcase
						end

						10'h1f5: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1f6;

									end
								end

							endcase
						end

						10'h1f6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp11758) ? 10'h1f9 : 10'h1fb);

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1f6;

									end
								end

							endcase
						end

						10'h1fb: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1fc;

									end
								end

							endcase
						end

						10'h1fc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp11854) ? 10'h1ff : 10'h201);

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1fc;

									end
								end

							endcase
						end

						10'h201: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h202;

									end
								end

							endcase
						end

						10'h202: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp11950) ? 10'h205 : 10'h207);

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h202;

									end
								end

							endcase
						end

						10'h207: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h208;

									end
								end

							endcase
						end

						10'h208: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp12046) ? 10'h20b : 10'h20d);

									end
								end

							endcase
						end

						10'h20b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h208;

									end
								end

							endcase
						end

						10'h20d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h20e;

									end
								end

							endcase
						end

						10'h20e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp12142) ? 10'h211 : 10'h213);

									end
								end

							endcase
						end

						10'h211: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h20e;

									end
								end

							endcase
						end

						10'h213: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h214;

									end
								end

							endcase
						end

						10'h214: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp12238) ? 10'h217 : 10'h1e6);

									end
								end

							endcase
						end

						10'h217: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h214;

									end
								end

							endcase
						end

						10'h218: begin
							r_sys_run_phase <= 10'h21b;
						end

						10'h219: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_run_phase <= 10'h218;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sys_run_phase <= 10'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 6'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'ha: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h20)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h10: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h13: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h15: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h16: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h19: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h21: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h22: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h23: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h26: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h27: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h2c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h2d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h32: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h33: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h38: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h39: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h3e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h3f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h44: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h45: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h48: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h4a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h4b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h4e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h50: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h51: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h54: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h56: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h57: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h58: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h5b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h5c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h61: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h62: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h67: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h68: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h6d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h6e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h73: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h74: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h79: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h7a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h7d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h7f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h80: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h83: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h85: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h86: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h89: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h8b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h8c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h8d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h90: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h91: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h96: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h97: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h9c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h9d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'ha2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'ha3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'ha8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'ha9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hae: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'haf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hb2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hb4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hb5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hb8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hba: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hbb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hbe: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hc0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hc1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hc2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hc5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hc6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hcb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hcc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hd1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hd2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hd7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hd8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hdd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hde: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'he3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'he4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'he9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hea: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hf0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hf3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hf6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hf7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1f: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hfd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hfe: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h103: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h104: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h109: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h10a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h10f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h110: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h115: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h116: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h11b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h11c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h121: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h122: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h127: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h128: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h12d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h12e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h133: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h134: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h139: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h13a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h13f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h140: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3a)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h145: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h146: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h147: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h14a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h14b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h150: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h151: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h156: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h157: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h15c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h15d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h162: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h163: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h168: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h169: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h16c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h16e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h16f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h172: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h174: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h175: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h178: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h17a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h17b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h17c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h17f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h180: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h185: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h186: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h18b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h18c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h191: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h192: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h197: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h198: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h19d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h19e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1a1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1a3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1a4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1a7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1a9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1aa: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1ad: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1af: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1b0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1b1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1b4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1b5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1ba: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1bb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1c0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1c1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1c6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1c7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1cc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1cd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1d2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1d3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1d6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1d8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1d9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1dc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1de: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1df: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1e2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1e4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1e5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1e6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1e9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1ea: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1ef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1f0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1f5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1f6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1fb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1fc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h201: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h202: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h207: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h208: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h20b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h20d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h20e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h211: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h213: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h214: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h217: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h219: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 6'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'ha: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h20)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h1f)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'hf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h10: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h13: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h3)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h15: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h16: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h19: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'hc)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h1b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h5)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h21: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h22: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h23: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h26: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h27: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h2c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h2d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h32: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h33: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h38: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h39: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h3e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h3f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h44: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h45: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h48: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h4a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h4b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h4e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h50: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h51: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h54: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h56: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h57: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h58: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h5b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h5c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h61: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h62: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h67: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h68: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h6d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h6e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h73: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h74: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h79: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h7a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h7d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h7f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h80: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h83: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h85: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h86: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h89: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h8b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h8c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h8d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h90: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h91: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h96: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h97: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h9c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h9d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'ha2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'ha3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'ha8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'ha9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'hae: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'haf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hb2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hb4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hb5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hb8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hba: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hbb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hbe: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hc0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hc1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hc2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hc5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hc6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hcb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hcc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hd1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hd2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hd7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hd8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'hdd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hde: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'he3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'he4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'he9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hea: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hf0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hf3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hf6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hf7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub00_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub01_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub02_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub03_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub04_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub05_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub06_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub07_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub08_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub09_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub10_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub11_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub12_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub13_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub14_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub15_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub16_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub17_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub18_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub19_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub20_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub21_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub22_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub23_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub24_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub25_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub26_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub27_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub28_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub29_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub30_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'h1f: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub31_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hfd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hfe: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h1c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h103: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h104: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h1c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h109: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h10a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h1c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h10f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h110: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h1c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h115: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h116: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h11b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h11c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h121: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h122: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h127: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h128: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h12d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h12e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h133: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h134: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h139: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h13a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h13f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h140: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h39)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h3a)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h145: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h146: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h147: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h14a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h14b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h150: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h151: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h156: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h157: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h15c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h15d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h162: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h163: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h168: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h169: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h16c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h16e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h16f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h172: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h174: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h175: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h178: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h17a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h17b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h17c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h17f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h180: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h185: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h186: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h18b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h18c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h191: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h192: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h197: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h198: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h19d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h19e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1a1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h1a3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1a4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1a7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1a9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1aa: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1ad: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h1af: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1b0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1b1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1b4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1b5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h1ba: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1bb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1c0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1c1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1c6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1c7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h1cc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1cd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1d2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1d3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1d6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1d8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1d9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1dc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1de: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1df: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1e2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1e4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1e5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1e6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1e9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1ea: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1ef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1f0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1f5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1f6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1fb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1fc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h201: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h202: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h207: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h208: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h20b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h20d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h20e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h211: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h213: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h214: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h217: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h219: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						10'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						10'h21b: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_T_0_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp22[14:0] );

									end
								end

							endcase
						end

						10'h13: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp193[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp189[14:0] );

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp197[14:0] );

									end
								end

							endcase
						end

						10'h19: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h2) || (r_sys_run_step==6'h4) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'hc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp207[14:0] );

									end
									else
									if((r_sys_run_step==6'h1) || (r_sys_run_step==6'h3) || (r_sys_run_step==6'h5) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h9) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp212[14:0] );

									end
								end

							endcase
						end

						10'h1f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp298[14:0] );

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp360[14:0] );

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp505[14:0] );

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp650[14:0] );

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp795[14:0] );

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp940[14:0] );

									end
								end

							endcase
						end

						10'h48: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1085[14:0] );

									end
								end

							endcase
						end

						10'h4e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1230[14:0] );

									end
								end

							endcase
						end

						10'h54: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1375[14:0] );

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1523[14:0] );

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1668[14:0] );

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1813[14:0] );

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1958[14:0] );

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2103[14:0] );

									end
								end

							endcase
						end

						10'h7d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2248[14:0] );

									end
								end

							endcase
						end

						10'h83: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2393[14:0] );

									end
								end

							endcase
						end

						10'h89: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2538[14:0] );

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2686[14:0] );

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2831[14:0] );

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2976[14:0] );

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3121[14:0] );

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3266[14:0] );

									end
								end

							endcase
						end

						10'hb2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3411[14:0] );

									end
								end

							endcase
						end

						10'hb8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3556[14:0] );

									end
								end

							endcase
						end

						10'hbe: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3701[14:0] );

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3849[14:0] );

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3994[14:0] );

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4139[14:0] );

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4284[14:0] );

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4429[14:0] );

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4574[14:0] );

									end
								end

							endcase
						end

						10'hed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4719[14:0] );

									end
								end

							endcase
						end

						10'hf3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4864[14:0] );

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9336[14:0] );

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9413[14:0] );

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9509[14:0] );

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9605[14:0] );

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9701[14:0] );

									end
								end

							endcase
						end

						10'h16c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9797[14:0] );

									end
								end

							endcase
						end

						10'h172: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9893[14:0] );

									end
								end

							endcase
						end

						10'h178: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9989[14:0] );

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10088[14:0] );

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10165[14:0] );

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10261[14:0] );

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10357[14:0] );

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10453[14:0] );

									end
								end

							endcase
						end

						10'h1a1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10549[14:0] );

									end
								end

							endcase
						end

						10'h1a7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10645[14:0] );

									end
								end

							endcase
						end

						10'h1ad: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10741[14:0] );

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10840[14:0] );

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10917[14:0] );

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11013[14:0] );

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11109[14:0] );

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11205[14:0] );

									end
								end

							endcase
						end

						10'h1d6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11301[14:0] );

									end
								end

							endcase
						end

						10'h1dc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11397[14:0] );

									end
								end

							endcase
						end

						10'h1e2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11493[14:0] );

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11592[14:0] );

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11669[14:0] );

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11765[14:0] );

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11861[14:0] );

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11957[14:0] );

									end
								end

							endcase
						end

						10'h20b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12053[14:0] );

									end
								end

							endcase
						end

						10'h211: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12149[14:0] );

									end
								end

							endcase
						end

						10'h217: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12245[14:0] );

									end
								end

							endcase
						end

						10'h219: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12334[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp25;

									end
								end

							endcase
						end

						10'h13: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp196;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp191;

									end
								end

							endcase
						end

						10'h19: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'hd)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp210;

									end
								end

							endcase
						end

						10'h1f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp301;

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp9339;

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp9416;

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp9512;

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp9608;

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp9704;

									end
								end

							endcase
						end

						10'h16c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp9800;

									end
								end

							endcase
						end

						10'h172: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp9896;

									end
								end

							endcase
						end

						10'h178: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp9992;

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp10091;

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp10168;

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp10264;

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp10360;

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp10456;

									end
								end

							endcase
						end

						10'h1a1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp10552;

									end
								end

							endcase
						end

						10'h1a7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp10648;

									end
								end

							endcase
						end

						10'h1ad: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp10744;

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp10843;

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp10920;

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp11016;

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp11112;

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp11208;

									end
								end

							endcase
						end

						10'h1d6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp11304;

									end
								end

							endcase
						end

						10'h1dc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp11400;

									end
								end

							endcase
						end

						10'h1e2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp11496;

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp11595;

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp11672;

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp11768;

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp11864;

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp11960;

									end
								end

							endcase
						end

						10'h20b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp12056;

									end
								end

							endcase
						end

						10'h211: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp12152;

									end
								end

							endcase
						end

						10'h217: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp12248;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_T_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h13: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h3)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h19: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'hd)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h48: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h4e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h54: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h7d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h83: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h89: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hb2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hb8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hbe: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hf3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h16c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h172: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h178: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1a1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1a7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1ad: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1d6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1dc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1e2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h20b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h211: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h217: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h219: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_fld_T_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_TT_1_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_TT_1_addr_1 <= $signed( w_sys_tmp27[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_TT_1_datain_1 <= w_sys_tmp25;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_TT_1_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_TT_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h21b: begin
							r_fld_TT_1_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_U_2_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h18) || (r_sys_run_step==6'h1a) || (6'h1c<=r_sys_run_step && r_sys_run_step<=6'h20)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp32[14:0] );

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp352[14:0] );

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp497[14:0] );

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp642[14:0] );

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp787[14:0] );

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp932[14:0] );

									end
								end

							endcase
						end

						10'h48: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1077[14:0] );

									end
								end

							endcase
						end

						10'h4e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1222[14:0] );

									end
								end

							endcase
						end

						10'h54: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1367[14:0] );

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1515[14:0] );

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1660[14:0] );

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1805[14:0] );

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1950[14:0] );

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2095[14:0] );

									end
								end

							endcase
						end

						10'h7d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2240[14:0] );

									end
								end

							endcase
						end

						10'h83: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2385[14:0] );

									end
								end

							endcase
						end

						10'h89: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2530[14:0] );

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2678[14:0] );

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2823[14:0] );

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2968[14:0] );

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3113[14:0] );

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3258[14:0] );

									end
								end

							endcase
						end

						10'hb2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3403[14:0] );

									end
								end

							endcase
						end

						10'hb8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3548[14:0] );

									end
								end

							endcase
						end

						10'hbe: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3693[14:0] );

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3841[14:0] );

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3986[14:0] );

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4131[14:0] );

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4276[14:0] );

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4421[14:0] );

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4566[14:0] );

									end
								end

							endcase
						end

						10'hed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4711[14:0] );

									end
								end

							endcase
						end

						10'hf3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4856[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h18) || (r_sys_run_step==6'h1a) || (6'h1c<=r_sys_run_step && r_sys_run_step<=6'h20)) begin
										r_fld_U_2_datain_1 <= w_sys_tmp18;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_U_2_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h18) || (r_sys_run_step==6'h1a) || (6'h1c<=r_sys_run_step && r_sys_run_step<=6'h20)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h48: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h4e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h54: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h7d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h83: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h89: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hb2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hb8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hbe: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hf3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_fld_U_2_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_35 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'h6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_35 <= w_sys_tmp14;

									end
								end

							endcase
						end

						10'hf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_35 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'h13: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_run_k_35 <= w_sys_tmp201;

									end
								end

							endcase
						end

						10'h21: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_35 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'h23: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_35 <= w_sys_tmp342;

									end
								end

							endcase
						end

						10'h56: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_35 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'h58: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_35 <= w_sys_tmp1505;

									end
								end

							endcase
						end

						10'h8b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_35 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'h8d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_35 <= w_sys_tmp2668;

									end
								end

							endcase
						end

						10'hc0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_35 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'hc2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_35 <= w_sys_tmp3831;

									end
								end

							endcase
						end

						10'hfd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_35 <= w_sys_tmp4994;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_run_k_35 <= w_sys_tmp5077;

									end
								end

							endcase
						end

						10'h103: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_35 <= w_sys_tmp5078;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_run_k_35 <= w_sys_tmp5161;

									end
								end

							endcase
						end

						10'h109: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_35 <= w_sys_tmp5162;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_run_k_35 <= w_sys_tmp5245;

									end
								end

							endcase
						end

						10'h10f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_35 <= w_sys_tmp5246;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_run_k_35 <= w_sys_tmp5329;

									end
								end

							endcase
						end

						10'h145: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_35 <= w_sys_tmp9325;

									end
								end

							endcase
						end

						10'h147: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_35 <= w_sys_tmp9329;

									end
								end

							endcase
						end

						10'h17a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_35 <= w_sys_tmp10077;

									end
								end

							endcase
						end

						10'h17c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_35 <= w_sys_tmp10081;

									end
								end

							endcase
						end

						10'h1af: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_35 <= w_sys_tmp10829;

									end
								end

							endcase
						end

						10'h1b1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_35 <= w_sys_tmp10833;

									end
								end

							endcase
						end

						10'h1e4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_35 <= w_sys_tmp11581;

									end
								end

							endcase
						end

						10'h1e6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_35 <= w_sys_tmp11585;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp42;

									end
								end

							endcase
						end

						10'h15: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'h19: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h2) || (r_sys_run_step==6'h4) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'hc)) begin
										r_run_j_36 <= w_sys_tmp217;

									end
								end

							endcase
						end

						10'h1b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp290;

									end
								end

							endcase
						end

						10'h1f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp302;

									end
								end

							endcase
						end

						10'h26: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp366;

									end
								end

							endcase
						end

						10'h2c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp487;

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp511;

									end
								end

							endcase
						end

						10'h32: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp632;

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp656;

									end
								end

							endcase
						end

						10'h38: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp777;

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp801;

									end
								end

							endcase
						end

						10'h3e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp922;

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp946;

									end
								end

							endcase
						end

						10'h44: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp1067;

									end
								end

							endcase
						end

						10'h48: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp1091;

									end
								end

							endcase
						end

						10'h4a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp1212;

									end
								end

							endcase
						end

						10'h4e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp1236;

									end
								end

							endcase
						end

						10'h50: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp1357;

									end
								end

							endcase
						end

						10'h54: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp1381;

									end
								end

							endcase
						end

						10'h5b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp1529;

									end
								end

							endcase
						end

						10'h61: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp1650;

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp1674;

									end
								end

							endcase
						end

						10'h67: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp1795;

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp1819;

									end
								end

							endcase
						end

						10'h6d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp1940;

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp1964;

									end
								end

							endcase
						end

						10'h73: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp2085;

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp2109;

									end
								end

							endcase
						end

						10'h79: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp2230;

									end
								end

							endcase
						end

						10'h7d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp2254;

									end
								end

							endcase
						end

						10'h7f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp2375;

									end
								end

							endcase
						end

						10'h83: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp2399;

									end
								end

							endcase
						end

						10'h85: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp2520;

									end
								end

							endcase
						end

						10'h89: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp2544;

									end
								end

							endcase
						end

						10'h90: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp2692;

									end
								end

							endcase
						end

						10'h96: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp2813;

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp2837;

									end
								end

							endcase
						end

						10'h9c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp2958;

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp2982;

									end
								end

							endcase
						end

						10'ha2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp3103;

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp3127;

									end
								end

							endcase
						end

						10'ha8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp3248;

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp3272;

									end
								end

							endcase
						end

						10'hae: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp3393;

									end
								end

							endcase
						end

						10'hb2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp3417;

									end
								end

							endcase
						end

						10'hb4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp3538;

									end
								end

							endcase
						end

						10'hb8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp3562;

									end
								end

							endcase
						end

						10'hba: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp3683;

									end
								end

							endcase
						end

						10'hbe: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp3707;

									end
								end

							endcase
						end

						10'hc5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp3855;

									end
								end

							endcase
						end

						10'hcb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp3976;

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp4000;

									end
								end

							endcase
						end

						10'hd1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp4121;

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp4145;

									end
								end

							endcase
						end

						10'hd7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp4266;

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp4290;

									end
								end

							endcase
						end

						10'hdd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp4411;

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp4435;

									end
								end

							endcase
						end

						10'he3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp4556;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp4580;

									end
								end

							endcase
						end

						10'he9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp4701;

									end
								end

							endcase
						end

						10'hed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp4725;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp4846;

									end
								end

							endcase
						end

						10'hf3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp4870;

									end
								end

							endcase
						end

						10'h115: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_36 <= w_sys_tmp5403;

									end
								end

							endcase
						end

						10'h11b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp5830;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_36 <= w_sys_tmp5904;

									end
								end

							endcase
						end

						10'h121: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp6331;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_36 <= w_sys_tmp6405;

									end
								end

							endcase
						end

						10'h127: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp6832;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_36 <= w_sys_tmp6906;

									end
								end

							endcase
						end

						10'h12d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp7333;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_36 <= w_sys_tmp7407;

									end
								end

							endcase
						end

						10'h133: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp7834;

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_36 <= w_sys_tmp7908;

									end
								end

							endcase
						end

						10'h139: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp8335;

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_36 <= w_sys_tmp8409;

									end
								end

							endcase
						end

						10'h13f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp8836;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_36 <= w_sys_tmp8910;

									end
								end

							endcase
						end

						10'h14a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp9330;

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp9344;

									end
								end

							endcase
						end

						10'h150: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp9405;

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp9422;

									end
								end

							endcase
						end

						10'h156: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp9501;

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp9518;

									end
								end

							endcase
						end

						10'h15c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp9597;

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp9614;

									end
								end

							endcase
						end

						10'h162: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp9693;

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp9710;

									end
								end

							endcase
						end

						10'h168: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp9789;

									end
								end

							endcase
						end

						10'h16c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp9806;

									end
								end

							endcase
						end

						10'h16e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp9885;

									end
								end

							endcase
						end

						10'h172: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp9902;

									end
								end

							endcase
						end

						10'h174: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp9981;

									end
								end

							endcase
						end

						10'h178: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp9998;

									end
								end

							endcase
						end

						10'h17f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp10082;

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp10096;

									end
								end

							endcase
						end

						10'h185: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp10157;

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp10174;

									end
								end

							endcase
						end

						10'h18b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp10253;

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp10270;

									end
								end

							endcase
						end

						10'h191: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp10349;

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp10366;

									end
								end

							endcase
						end

						10'h197: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp10445;

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp10462;

									end
								end

							endcase
						end

						10'h19d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp10541;

									end
								end

							endcase
						end

						10'h1a1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp10558;

									end
								end

							endcase
						end

						10'h1a3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp10637;

									end
								end

							endcase
						end

						10'h1a7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp10654;

									end
								end

							endcase
						end

						10'h1a9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp10733;

									end
								end

							endcase
						end

						10'h1ad: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp10750;

									end
								end

							endcase
						end

						10'h1b4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp10834;

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp10848;

									end
								end

							endcase
						end

						10'h1ba: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp10909;

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp10926;

									end
								end

							endcase
						end

						10'h1c0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp11005;

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp11022;

									end
								end

							endcase
						end

						10'h1c6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp11101;

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp11118;

									end
								end

							endcase
						end

						10'h1cc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp11197;

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp11214;

									end
								end

							endcase
						end

						10'h1d2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp11293;

									end
								end

							endcase
						end

						10'h1d6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp11310;

									end
								end

							endcase
						end

						10'h1d8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp11389;

									end
								end

							endcase
						end

						10'h1dc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp11406;

									end
								end

							endcase
						end

						10'h1de: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp11485;

									end
								end

							endcase
						end

						10'h1e2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp11502;

									end
								end

							endcase
						end

						10'h1e9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp11586;

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_36 <= w_sys_tmp11600;

									end
								end

							endcase
						end

						10'h1ef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp11661;

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp11678;

									end
								end

							endcase
						end

						10'h1f5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp11757;

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp11774;

									end
								end

							endcase
						end

						10'h1fb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp11853;

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp11870;

									end
								end

							endcase
						end

						10'h201: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp11949;

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp11966;

									end
								end

							endcase
						end

						10'h207: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp12045;

									end
								end

							endcase
						end

						10'h20b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp12062;

									end
								end

							endcase
						end

						10'h20d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp12141;

									end
								end

							endcase
						end

						10'h211: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp12158;

									end
								end

							endcase
						end

						10'h213: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_36 <= w_sys_tmp12237;

									end
								end

							endcase
						end

						10'h217: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_36 <= w_sys_tmp12254;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_n_37 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'hf7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_n_37 <= w_sys_tmp4993;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_mx_38 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_my_39 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_dt_40 <= w_sys_tmp5;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_dx_41 <= w_sys_tmp6;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_dy_42 <= w_sys_tmp7;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_r1_43 <= w_sys_tmp8;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_r2_44 <= w_sys_tmp9;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_r3_45 <= w_sys_tmp10;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_r4_46 <= w_sys_tmp11;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h10) || (r_sys_run_step==6'h11)) begin
										r_run_YY_47 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'hc) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h14)) begin
										r_run_YY_47 <= w_sys_tmp18;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_kx_48 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_ky_49 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_nlast_50 <= w_sys_intOne;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h154: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_51 <= w_sys_tmp9410;

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_51 <= w_sys_tmp9506;

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_51 <= w_sys_tmp9602;

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_51 <= w_sys_tmp9698;

									end
								end

							endcase
						end

						10'h16c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_51 <= w_sys_tmp9794;

									end
								end

							endcase
						end

						10'h172: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_51 <= w_sys_tmp9890;

									end
								end

							endcase
						end

						10'h178: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_51 <= w_sys_tmp9986;

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_51 <= w_sys_tmp10162;

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_51 <= w_sys_tmp10258;

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_51 <= w_sys_tmp10354;

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_51 <= w_sys_tmp10450;

									end
								end

							endcase
						end

						10'h1a1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_51 <= w_sys_tmp10546;

									end
								end

							endcase
						end

						10'h1a7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_51 <= w_sys_tmp10642;

									end
								end

							endcase
						end

						10'h1ad: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_51 <= w_sys_tmp10738;

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_51 <= w_sys_tmp10914;

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_51 <= w_sys_tmp11010;

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_51 <= w_sys_tmp11106;

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_51 <= w_sys_tmp11202;

									end
								end

							endcase
						end

						10'h1d6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_51 <= w_sys_tmp11298;

									end
								end

							endcase
						end

						10'h1dc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_51 <= w_sys_tmp11394;

									end
								end

							endcase
						end

						10'h1e2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_51 <= w_sys_tmp11490;

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_51 <= w_sys_tmp11666;

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_51 <= w_sys_tmp11762;

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_51 <= w_sys_tmp11858;

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_51 <= w_sys_tmp11954;

									end
								end

							endcase
						end

						10'h20b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_51 <= w_sys_tmp12050;

									end
								end

							endcase
						end

						10'h211: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_51 <= w_sys_tmp12146;

									end
								end

							endcase
						end

						10'h217: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_51 <= w_sys_tmp12242;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_52 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h18) || (r_sys_run_step==6'h1a) || (6'h1c<=r_sys_run_step && r_sys_run_step<=6'h20)) begin
										r_run_copy0_j_52 <= w_sys_tmp40;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_53 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy1_j_53 <= w_sys_tmp41;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h15: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_54 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h19: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1) || (r_sys_run_step==6'h3) || (r_sys_run_step==6'h5) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h9) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hd)) begin
										r_run_copy0_j_54 <= w_sys_tmp216;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h26: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_55 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_55 <= w_sys_tmp363;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h26: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_56 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_56 <= w_sys_tmp364;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h26: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_57 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_57 <= w_sys_tmp365;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2c: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_58 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_58 <= w_sys_tmp508;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2c: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_59 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_59 <= w_sys_tmp509;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2c: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_60 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_60 <= w_sys_tmp510;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h32: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_61 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_61 <= w_sys_tmp653;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h32: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_62 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_62 <= w_sys_tmp654;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h32: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_63 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_63 <= w_sys_tmp655;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h38: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_64 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_64 <= w_sys_tmp798;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h38: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_65 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_65 <= w_sys_tmp799;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h38: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_66 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_66 <= w_sys_tmp800;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h3e: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_67 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_67 <= w_sys_tmp943;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h3e: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_68 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_68 <= w_sys_tmp944;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h3e: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_69 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_69 <= w_sys_tmp945;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h44: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_70 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h48: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_70 <= w_sys_tmp1088;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h44: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_71 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h48: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_71 <= w_sys_tmp1089;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h44: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_72 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h48: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_72 <= w_sys_tmp1090;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4a: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_73 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h4e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_73 <= w_sys_tmp1233;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4a: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_74 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h4e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_74 <= w_sys_tmp1234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4a: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_75 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h4e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_75 <= w_sys_tmp1235;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h50: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_76 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h54: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_76 <= w_sys_tmp1378;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h50: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_77 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h54: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_77 <= w_sys_tmp1379;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h50: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_78 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h54: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_78 <= w_sys_tmp1380;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h5b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_79 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_79 <= w_sys_tmp1526;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h5b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_80 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_80 <= w_sys_tmp1527;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h5b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_81 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_81 <= w_sys_tmp1528;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h61: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_82 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_82 <= w_sys_tmp1671;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h61: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_83 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_83 <= w_sys_tmp1672;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h61: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_84 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_84 <= w_sys_tmp1673;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h67: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_85 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_85 <= w_sys_tmp1816;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h67: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_86 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_86 <= w_sys_tmp1817;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h67: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_87 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_87 <= w_sys_tmp1818;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h6d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_88 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_88 <= w_sys_tmp1961;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h6d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_89 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_89 <= w_sys_tmp1962;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h6d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_90 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_90 <= w_sys_tmp1963;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h73: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_91 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_91 <= w_sys_tmp2106;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h73: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_92 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_92 <= w_sys_tmp2107;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h73: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_93 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_93 <= w_sys_tmp2108;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h79: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_94 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h7d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_94 <= w_sys_tmp2251;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h79: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_95 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h7d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_95 <= w_sys_tmp2252;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h79: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_96 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h7d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_96 <= w_sys_tmp2253;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h7f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_97 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h83: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_97 <= w_sys_tmp2396;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h7f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_98 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h83: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_98 <= w_sys_tmp2397;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h7f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_99 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h83: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_99 <= w_sys_tmp2398;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h85: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_100 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h89: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_100 <= w_sys_tmp2541;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h85: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_101 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h89: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_101 <= w_sys_tmp2542;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h85: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_102 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h89: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_102 <= w_sys_tmp2543;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h90: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_103 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_103 <= w_sys_tmp2689;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h90: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_104 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_104 <= w_sys_tmp2690;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h90: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_105 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_105 <= w_sys_tmp2691;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h96: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_106 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_106 <= w_sys_tmp2834;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h96: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_107 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_107 <= w_sys_tmp2835;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h96: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_108 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_108 <= w_sys_tmp2836;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9c: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_109 <= r_run_j_36;

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_109 <= w_sys_tmp2979;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9c: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_110 <= r_run_j_36;

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_110 <= w_sys_tmp2980;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9c: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_111 <= r_run_j_36;

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_111 <= w_sys_tmp2981;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha2: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_112 <= r_run_j_36;

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_112 <= w_sys_tmp3124;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha2: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_113 <= r_run_j_36;

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_113 <= w_sys_tmp3125;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha2: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_114 <= r_run_j_36;

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_114 <= w_sys_tmp3126;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha8: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_115 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_115 <= w_sys_tmp3269;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha8: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_116 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_116 <= w_sys_tmp3270;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha8: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_117 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_117 <= w_sys_tmp3271;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hae: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_118 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hb2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_118 <= w_sys_tmp3414;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hae: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_119 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hb2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_119 <= w_sys_tmp3415;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hae: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_120 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hb2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_120 <= w_sys_tmp3416;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb4: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_121 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hb8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_121 <= w_sys_tmp3559;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb4: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_122 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hb8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_122 <= w_sys_tmp3560;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb4: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_123 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hb8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_123 <= w_sys_tmp3561;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hba: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_124 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hbe: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_124 <= w_sys_tmp3704;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hba: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_125 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hbe: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_125 <= w_sys_tmp3705;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hba: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_126 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hbe: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_126 <= w_sys_tmp3706;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc5: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_127 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_127 <= w_sys_tmp3852;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc5: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_128 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_128 <= w_sys_tmp3853;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc5: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_129 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_129 <= w_sys_tmp3854;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hcb: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_130 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_130 <= w_sys_tmp3997;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hcb: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_131 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_131 <= w_sys_tmp3998;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hcb: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_132 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_132 <= w_sys_tmp3999;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd1: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_133 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_133 <= w_sys_tmp4142;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd1: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_134 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_134 <= w_sys_tmp4143;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd1: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_135 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_135 <= w_sys_tmp4144;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd7: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_136 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_136 <= w_sys_tmp4287;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd7: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_137 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_137 <= w_sys_tmp4288;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd7: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_138 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_138 <= w_sys_tmp4289;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hdd: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_139 <= r_run_j_36;

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_139 <= w_sys_tmp4432;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hdd: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_140 <= r_run_j_36;

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_140 <= w_sys_tmp4433;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hdd: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_141 <= r_run_j_36;

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_141 <= w_sys_tmp4434;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he3: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_142 <= r_run_j_36;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_142 <= w_sys_tmp4577;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he3: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_143 <= r_run_j_36;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_143 <= w_sys_tmp4578;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he3: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_144 <= r_run_j_36;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_144 <= w_sys_tmp4579;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he9: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_145 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_145 <= w_sys_tmp4722;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he9: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_146 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_146 <= w_sys_tmp4723;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he9: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_147 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_147 <= w_sys_tmp4724;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_148 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hf3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_148 <= w_sys_tmp4867;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_149 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hf3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_149 <= w_sys_tmp4868;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_150 <= r_run_j_36;

									end
								end

							endcase
						end

						10'hf3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_150 <= w_sys_tmp4869;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_151 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_151 <= w_sys_tmp5392;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_152 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_152 <= w_sys_tmp5393;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_153 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_153 <= w_sys_tmp5394;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_154 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_154 <= w_sys_tmp5395;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_155 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_155 <= w_sys_tmp5396;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_156 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_156 <= w_sys_tmp5397;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_157 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_157 <= w_sys_tmp5398;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_158 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_158 <= w_sys_tmp5399;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_159 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_159 <= w_sys_tmp5400;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_160 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_160 <= w_sys_tmp5401;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_161 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_161 <= w_sys_tmp5402;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_162 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_162 <= w_sys_tmp5893;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_163 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_163 <= w_sys_tmp5894;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_164 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_164 <= w_sys_tmp5895;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_165 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_165 <= w_sys_tmp5896;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_166 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_166 <= w_sys_tmp5897;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_167 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_167 <= w_sys_tmp5898;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_168 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_168 <= w_sys_tmp5899;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_169 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_169 <= w_sys_tmp5900;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_170 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_170 <= w_sys_tmp5901;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_171 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_171 <= w_sys_tmp5902;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_172 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_172 <= w_sys_tmp5903;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_173 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_173 <= w_sys_tmp6394;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_174 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_174 <= w_sys_tmp6395;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_175 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_175 <= w_sys_tmp6396;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_176 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_176 <= w_sys_tmp6397;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_177 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_177 <= w_sys_tmp6398;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_178 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_178 <= w_sys_tmp6399;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_179 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_179 <= w_sys_tmp6400;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_180 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_180 <= w_sys_tmp6401;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_181 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_181 <= w_sys_tmp6402;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_182 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_182 <= w_sys_tmp6403;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_183 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_183 <= w_sys_tmp6404;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_184 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_184 <= w_sys_tmp6895;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_185 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_185 <= w_sys_tmp6896;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_186 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_186 <= w_sys_tmp6897;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_187 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_187 <= w_sys_tmp6898;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_188 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_188 <= w_sys_tmp6899;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_189 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_189 <= w_sys_tmp6900;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_190 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_190 <= w_sys_tmp6901;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_191 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_191 <= w_sys_tmp6902;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_192 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_192 <= w_sys_tmp6903;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_193 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_193 <= w_sys_tmp6904;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_194 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_194 <= w_sys_tmp6905;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_195 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_195 <= w_sys_tmp7396;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_196 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_196 <= w_sys_tmp7397;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_197 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_197 <= w_sys_tmp7398;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_198 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_198 <= w_sys_tmp7399;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_199 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_199 <= w_sys_tmp7400;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_200 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_200 <= w_sys_tmp7401;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_201 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_201 <= w_sys_tmp7402;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_202 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_202 <= w_sys_tmp7403;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_203 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_203 <= w_sys_tmp7404;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_204 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_204 <= w_sys_tmp7405;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_205 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_205 <= w_sys_tmp7406;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h133: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_206 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_206 <= w_sys_tmp7897;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h133: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_207 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_207 <= w_sys_tmp7898;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h133: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_208 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_208 <= w_sys_tmp7899;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h133: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_209 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_209 <= w_sys_tmp7900;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h133: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_210 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_210 <= w_sys_tmp7901;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h133: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_211 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_211 <= w_sys_tmp7902;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h133: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_212 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_212 <= w_sys_tmp7903;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h133: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_213 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_213 <= w_sys_tmp7904;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h133: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_214 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_214 <= w_sys_tmp7905;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h133: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_215 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_215 <= w_sys_tmp7906;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h133: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_216 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_216 <= w_sys_tmp7907;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h139: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_217 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_217 <= w_sys_tmp8398;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h139: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_218 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_218 <= w_sys_tmp8399;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h139: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_219 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_219 <= w_sys_tmp8400;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h139: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_220 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_220 <= w_sys_tmp8401;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h139: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_221 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_221 <= w_sys_tmp8402;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h139: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_222 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_222 <= w_sys_tmp8403;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h139: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_223 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_223 <= w_sys_tmp8404;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h139: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_224 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_224 <= w_sys_tmp8405;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h139: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_225 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_225 <= w_sys_tmp8406;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h139: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_226 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_226 <= w_sys_tmp8407;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h139: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_227 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_227 <= w_sys_tmp8408;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h13f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_228 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_228 <= w_sys_tmp8899;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h13f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_229 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h4) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'he)) begin
										r_run_copy1_j_229 <= w_sys_tmp8900;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h13f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_230 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h3) || (r_sys_run_step==6'h5) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h9) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hd)) begin
										r_run_copy2_j_230 <= w_sys_tmp8901;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h13f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_231 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_231 <= w_sys_tmp8902;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h13f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_232 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_232 <= w_sys_tmp8903;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h13f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_233 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_233 <= w_sys_tmp8904;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h13f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_234 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy6_j_234 <= w_sys_tmp8905;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h13f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_235 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_235 <= w_sys_tmp8906;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h13f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_236 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_236 <= w_sys_tmp8907;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h13f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_237 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_237 <= w_sys_tmp8908;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h13f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_238 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_238 <= w_sys_tmp8909;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h14a: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_239 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_239 <= w_sys_tmp9343;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h150: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_240 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_240 <= w_sys_tmp9420;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h150: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_241 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_241 <= w_sys_tmp9421;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h156: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_242 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_242 <= w_sys_tmp9516;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h156: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_243 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_243 <= w_sys_tmp9517;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h15c: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_244 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_244 <= w_sys_tmp9612;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h15c: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_245 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_245 <= w_sys_tmp9613;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h162: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_246 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_246 <= w_sys_tmp9708;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h162: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_247 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_247 <= w_sys_tmp9709;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h168: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_248 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h16c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_248 <= w_sys_tmp9804;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h168: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_249 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h16c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_249 <= w_sys_tmp9805;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h16e: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_250 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h172: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_250 <= w_sys_tmp9900;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h16e: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_251 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h172: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_251 <= w_sys_tmp9901;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h174: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_252 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h178: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_252 <= w_sys_tmp9996;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h174: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_253 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h178: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_253 <= w_sys_tmp9997;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h17f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_254 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_254 <= w_sys_tmp10095;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h185: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_255 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_255 <= w_sys_tmp10172;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h185: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_256 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_256 <= w_sys_tmp10173;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h18b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_257 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_257 <= w_sys_tmp10268;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h18b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_258 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_258 <= w_sys_tmp10269;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h191: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_259 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_259 <= w_sys_tmp10364;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h191: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_260 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_260 <= w_sys_tmp10365;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h197: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_261 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_261 <= w_sys_tmp10460;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h197: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_262 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_262 <= w_sys_tmp10461;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h19d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_263 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h1a1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_263 <= w_sys_tmp10556;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h19d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_264 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h1a1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_264 <= w_sys_tmp10557;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1a3: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_265 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h1a7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_265 <= w_sys_tmp10652;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1a3: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_266 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h1a7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_266 <= w_sys_tmp10653;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1a9: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_267 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h1ad: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_267 <= w_sys_tmp10748;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1a9: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_268 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h1ad: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_268 <= w_sys_tmp10749;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1b4: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_269 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_269 <= w_sys_tmp10847;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1ba: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_270 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_270 <= w_sys_tmp10924;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1ba: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_271 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_271 <= w_sys_tmp10925;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1c0: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_272 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_272 <= w_sys_tmp11020;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1c0: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_273 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_273 <= w_sys_tmp11021;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1c6: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_274 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_274 <= w_sys_tmp11116;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1c6: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_275 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_275 <= w_sys_tmp11117;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1cc: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_276 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_276 <= w_sys_tmp11212;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1cc: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_277 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_277 <= w_sys_tmp11213;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1d2: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_278 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h1d6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_278 <= w_sys_tmp11308;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1d2: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_279 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h1d6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_279 <= w_sys_tmp11309;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1d8: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_280 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h1dc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_280 <= w_sys_tmp11404;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1d8: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_281 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h1dc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_281 <= w_sys_tmp11405;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1de: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_282 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h1e2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_282 <= w_sys_tmp11500;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1de: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_283 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h1e2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_283 <= w_sys_tmp11501;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1e9: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_284 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_284 <= w_sys_tmp11599;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1ef: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_285 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_285 <= w_sys_tmp11676;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1ef: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_286 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_286 <= w_sys_tmp11677;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1f5: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_287 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_287 <= w_sys_tmp11772;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1f5: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_288 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_288 <= w_sys_tmp11773;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1fb: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_289 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_289 <= w_sys_tmp11868;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1fb: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_290 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_290 <= w_sys_tmp11869;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h201: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_291 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_291 <= w_sys_tmp11964;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h201: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_292 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_292 <= w_sys_tmp11965;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h207: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_293 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h20b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_293 <= w_sys_tmp12060;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h207: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_294 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h20b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_294 <= w_sys_tmp12061;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h20d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_295 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h211: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_295 <= w_sys_tmp12156;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h20d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_296 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h211: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_296 <= w_sys_tmp12157;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h213: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_297 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h217: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_297 <= w_sys_tmp12252;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h213: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_298 <= r_run_j_36;

									end
								end

							endcase
						end

						10'h217: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_298 <= w_sys_tmp12253;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub19_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp3117[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub19_T_datain <= w_sys_tmp3120;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub19_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub19_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp3109[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub19_U_datain <= w_sys_tmp3112;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub19_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub19_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hf)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp5168[11:0] );

									end
									else
									if((r_sys_run_step==6'he)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp5180[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp5171[11:0] );

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp5174[11:0] );

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp6862[11:0] );

									end
									else
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp6891[11:0] );

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp6877[11:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp6867[11:0] );

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp11113[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'he)) begin
										r_sub19_result_datain <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_sub19_result_datain <= w_sys_tmp5198;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub19_result_datain <= w_sys_tmp6842;

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub19_result_datain <= r_sys_tmp3_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'he)) begin
										r_sub19_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'hf)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub19_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub19_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub12_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h77: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp2099[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h77: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_T_datain <= w_sys_tmp2102;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h77: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub12_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h77: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp2091[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h77: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_U_datain <= w_sys_tmp2094;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h77: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub12_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h12)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5096[11:0] );

									end
									else
									if((r_sys_run_step==6'h11)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5090[11:0] );

									end
									else
									if((r_sys_run_step==6'h13)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5084[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5087[11:0] );

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp7349[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp7344[11:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp7359[11:0] );

									end
									else
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp7373[11:0] );

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp10457[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h11)) begin
										r_sub12_result_datain <= w_sys_tmp5125;

									end
									else
									if((r_sys_run_step==6'h12)) begin
										r_sub12_result_datain <= r_sys_tmp1_float;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub12_result_datain <= w_sys_tmp7353;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub12_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub12_result_datain <= w_sys_tmp7391;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h11) || (r_sys_run_step==6'h12)) begin
										r_sub12_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h13)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub12_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub12_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub11_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h71: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp1954[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h71: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_T_datain <= w_sys_tmp1957;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h71: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub11_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_V_addr <= 12'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub11_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h71: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp1946[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h71: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_U_datain <= w_sys_tmp1949;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h71: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub11_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'he)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5096[11:0] );

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5090[11:0] );

									end
									else
									if((r_sys_run_step==6'hf)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5084[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5087[11:0] );

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp6848[11:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp6858[11:0] );

									end
									else
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp6872[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp6843[11:0] );

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp10361[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'he)) begin
										r_sub11_result_datain <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_sub11_result_datain <= w_sys_tmp5114;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub11_result_datain <= w_sys_tmp6890;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub11_result_datain <= w_sys_tmp6852;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub11_result_datain <= r_sys_tmp1_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'he)) begin
										r_sub11_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hf)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub11_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub11_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub14_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h83: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp2389[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h83: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_T_datain <= w_sys_tmp2392;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h83: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub14_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h83: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp2381[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h83: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_U_datain <= w_sys_tmp2384;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h83: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub14_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1a)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5096[11:0] );

									end
									else
									if((r_sys_run_step==6'h19)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5090[11:0] );

									end
									else
									if((r_sys_run_step==6'h1b)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5084[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5087[11:0] );

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp8351[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp8346[11:0] );

									end
									else
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp8375[11:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp8361[11:0] );

									end
								end

							endcase
						end

						10'h1a7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp10649[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1a)) begin
										r_sub14_result_datain <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==6'h19)) begin
										r_sub14_result_datain <= w_sys_tmp5147;

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub14_result_datain <= w_sys_tmp8393;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub14_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub14_result_datain <= w_sys_tmp8355;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a)) begin
										r_sub14_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1b)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub14_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h1a7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub14_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub13_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h7d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp2244[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h7d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_T_datain <= w_sys_tmp2247;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h7d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub13_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h7d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp2236[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h7d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_U_datain <= w_sys_tmp2239;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h7d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub13_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h16)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5096[11:0] );

									end
									else
									if((r_sys_run_step==6'h15)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5090[11:0] );

									end
									else
									if((r_sys_run_step==6'h17)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5084[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5087[11:0] );

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp7850[11:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp7860[11:0] );

									end
									else
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp7874[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp7845[11:0] );

									end
								end

							endcase
						end

						10'h1a1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp10553[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h15)) begin
										r_sub13_result_datain <= w_sys_tmp5136;

									end
									else
									if((r_sys_run_step==6'h16)) begin
										r_sub13_result_datain <= r_sys_tmp3_float;

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub13_result_datain <= w_sys_tmp7854;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub13_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub13_result_datain <= w_sys_tmp7892;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h15) || (r_sys_run_step==6'h16)) begin
										r_sub13_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h17)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub13_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h1a1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub13_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub16_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h94: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp2682[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h94: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub16_T_datain <= w_sys_tmp2685;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h94: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub16_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub16_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h94: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp2674[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h94: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub16_U_datain <= w_sys_tmp2677;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h94: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub16_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub16_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp5168[11:0] );

									end
									else
									if((r_sys_run_step==6'h3)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp5177[11:0] );

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp5359[11:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp5364[11:0] );

									end
									else
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp5388[11:0] );

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp5374[11:0] );

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp8895[11:0] );

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp10844[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub16_result_datain <= w_sys_tmp5170;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub16_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub16_result_datain <= w_sys_tmp5339;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub16_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h3)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub16_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub16_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub15_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h89: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp2534[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h89: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_T_datain <= w_sys_tmp2537;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h89: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub15_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h89: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp2526[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h89: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_U_datain <= w_sys_tmp2529;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h89: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub15_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp5090[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp5087[11:0] );

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp8847[11:0] );

									end
									else
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp8876[11:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp8862[11:0] );

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp8852[11:0] );

									end
								end

							endcase
						end

						10'h1ad: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp10745[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sub15_result_datain <= w_sys_tmp5158;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub15_result_datain <= w_sys_tmp8856;

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub15_result_datain <= r_sys_tmp7_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sub15_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub15_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h1ad: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub15_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub18_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp2972[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub18_T_datain <= w_sys_tmp2975;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub18_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub18_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp2964[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub18_U_datain <= w_sys_tmp2967;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub18_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub18_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hb)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp5168[11:0] );

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp5180[11:0] );

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp5174[11:0] );

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp6366[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp6361[11:0] );

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp6376[11:0] );

									end
									else
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp6390[11:0] );

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp11017[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9)) begin
										r_sub18_result_datain <= w_sys_tmp5170;

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_sub18_result_datain <= r_sys_tmp5_float;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub18_result_datain <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub18_result_datain <= w_sys_tmp6341;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha)) begin
										r_sub18_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'hb)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub18_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub18_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub17_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp2827[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub17_T_datain <= w_sys_tmp2830;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub17_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub17_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp2819[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub17_U_datain <= w_sys_tmp2822;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub17_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub17_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h7)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp5168[11:0] );

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp5180[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp5171[11:0] );

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp5174[11:0] );

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp5889[11:0] );

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp5875[11:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp5865[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp5860[11:0] );

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp10921[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub17_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub17_result_datain <= w_sys_tmp5176;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub17_result_datain <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub17_result_datain <= w_sys_tmp5840;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6)) begin
										r_sub17_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub17_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub17_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub20_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp3262[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub20_T_datain <= w_sys_tmp3265;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub20_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub20_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp3254[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub20_U_datain <= w_sys_tmp3257;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub20_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub20_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h13)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp5168[11:0] );

									end
									else
									if((r_sys_run_step==6'h12)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp5180[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp5171[11:0] );

									end
									else
									if((r_sys_run_step==6'h11)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp5174[11:0] );

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp7392[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp7363[11:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp7368[11:0] );

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp7378[11:0] );

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp11209[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h12)) begin
										r_sub20_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h11)) begin
										r_sub20_result_datain <= w_sys_tmp5209;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub20_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub20_result_datain <= w_sys_tmp7343;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h11) || (r_sys_run_step==6'h12)) begin
										r_sub20_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h13)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub20_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub20_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub21_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp3407[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub21_T_datain <= w_sys_tmp3410;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub21_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub21_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp3399[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub21_U_datain <= w_sys_tmp3402;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub21_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub21_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h17)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp5168[11:0] );

									end
									else
									if((r_sys_run_step==6'h16)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp5180[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp5171[11:0] );

									end
									else
									if((r_sys_run_step==6'h15)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp5174[11:0] );

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp7879[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp7864[11:0] );

									end
									else
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp7893[11:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp7869[11:0] );

									end
								end

							endcase
						end

						10'h1d6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp11305[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h15)) begin
										r_sub21_result_datain <= w_sys_tmp5220;

									end
									else
									if((r_sys_run_step==6'h16)) begin
										r_sub21_result_datain <= r_sys_tmp3_float;

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub21_result_datain <= w_sys_tmp7844;

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub21_result_datain <= r_sys_tmp5_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h15) || (r_sys_run_step==6'h16)) begin
										r_sub21_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h17)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub21_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h1d6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub21_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub28_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub28_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub28_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub28_T_addr <= $signed( w_sys_tmp4425[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub28_T_datain <= w_sys_tmp4428;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub28_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub28_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub28_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub28_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub28_U_addr <= $signed( w_sys_tmp4417[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub28_U_datain <= w_sys_tmp4420;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub28_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub28_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub28_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub28_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h11)) begin
										r_sub28_result_addr <= $signed( w_sys_tmp5258[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_addr <= $signed( w_sys_tmp5255[11:0] );

									end
									else
									if((r_sys_run_step==6'h13)) begin
										r_sub28_result_addr <= $signed( w_sys_tmp5252[11:0] );

									end
									else
									if((r_sys_run_step==6'h12)) begin
										r_sub28_result_addr <= $signed( w_sys_tmp5264[11:0] );

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub28_result_addr <= $signed( w_sys_tmp7387[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub28_result_addr <= $signed( w_sys_tmp7382[11:0] );

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub28_result_addr <= $signed( w_sys_tmp11961[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h12)) begin
										r_sub28_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h11)) begin
										r_sub28_result_datain <= w_sys_tmp5293;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub28_result_datain <= w_sys_tmp7391;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub28_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h11) || (r_sys_run_step==6'h12)) begin
										r_sub28_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h13)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub28_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub28_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub29_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub29_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub29_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub29_T_addr <= $signed( w_sys_tmp4570[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub29_T_datain <= w_sys_tmp4573;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub29_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub29_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub29_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub29_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub29_U_addr <= $signed( w_sys_tmp4562[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub29_U_datain <= w_sys_tmp4565;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub29_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub29_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub29_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub29_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h15)) begin
										r_sub29_result_addr <= $signed( w_sys_tmp5258[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_addr <= $signed( w_sys_tmp5255[11:0] );

									end
									else
									if((r_sys_run_step==6'h17)) begin
										r_sub29_result_addr <= $signed( w_sys_tmp5252[11:0] );

									end
									else
									if((r_sys_run_step==6'h16)) begin
										r_sub29_result_addr <= $signed( w_sys_tmp5264[11:0] );

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub29_result_addr <= $signed( w_sys_tmp7888[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub29_result_addr <= $signed( w_sys_tmp7883[11:0] );

									end
								end

							endcase
						end

						10'h20b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub29_result_addr <= $signed( w_sys_tmp12057[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h15)) begin
										r_sub29_result_datain <= w_sys_tmp5304;

									end
									else
									if((r_sys_run_step==6'h16)) begin
										r_sub29_result_datain <= r_sys_tmp3_float;

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub29_result_datain <= w_sys_tmp7892;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub29_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h15) || (r_sys_run_step==6'h16)) begin
										r_sub29_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h17)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub29_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h20b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub29_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub26_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub26_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub26_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub26_T_addr <= $signed( w_sys_tmp4135[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub26_T_datain <= w_sys_tmp4138;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub26_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub26_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub26_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub26_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub26_U_addr <= $signed( w_sys_tmp4127[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub26_U_datain <= w_sys_tmp4130;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub26_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub26_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub26_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub26_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9)) begin
										r_sub26_result_addr <= $signed( w_sys_tmp5258[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_addr <= $signed( w_sys_tmp5255[11:0] );

									end
									else
									if((r_sys_run_step==6'hb)) begin
										r_sub26_result_addr <= $signed( w_sys_tmp5252[11:0] );

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_sub26_result_addr <= $signed( w_sys_tmp5264[11:0] );

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub26_result_addr <= $signed( w_sys_tmp6380[11:0] );

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub26_result_addr <= $signed( w_sys_tmp6385[11:0] );

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub26_result_addr <= $signed( w_sys_tmp11769[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9)) begin
										r_sub26_result_datain <= w_sys_tmp5254;

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_sub26_result_datain <= r_sys_tmp0_float;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub26_result_datain <= w_sys_tmp6389;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub26_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha)) begin
										r_sub26_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub26_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub26_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub09_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h65: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp1664[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h65: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_T_datain <= w_sys_tmp1667;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h65: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub09_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h65: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp1656[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h65: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_U_datain <= w_sys_tmp1659;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h65: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub09_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5096[11:0] );

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5090[11:0] );

									end
									else
									if((r_sys_run_step==6'h7)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5084[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5087[11:0] );

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5846[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5841[11:0] );

									end
									else
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5870[11:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5856[11:0] );

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp10169[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub09_result_datain <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub09_result_datain <= w_sys_tmp5092;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub09_result_datain <= w_sys_tmp5850;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub09_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub09_result_datain <= w_sys_tmp5888;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6)) begin
										r_sub09_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub09_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub09_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub27_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub27_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub27_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hdb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub27_T_addr <= $signed( w_sys_tmp4280[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hdb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub27_T_datain <= w_sys_tmp4283;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub27_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hdb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub27_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub27_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub27_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hdb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub27_U_addr <= $signed( w_sys_tmp4272[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hdb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub27_U_datain <= w_sys_tmp4275;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub27_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hdb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub27_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub27_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub27_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub27_result_addr <= $signed( w_sys_tmp5258[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_addr <= $signed( w_sys_tmp5255[11:0] );

									end
									else
									if((r_sys_run_step==6'hf)) begin
										r_sub27_result_addr <= $signed( w_sys_tmp5252[11:0] );

									end
									else
									if((r_sys_run_step==6'he)) begin
										r_sub27_result_addr <= $signed( w_sys_tmp5264[11:0] );

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub27_result_addr <= $signed( w_sys_tmp6886[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub27_result_addr <= $signed( w_sys_tmp6881[11:0] );

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub27_result_addr <= $signed( w_sys_tmp11865[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'he)) begin
										r_sub27_result_datain <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_sub27_result_datain <= w_sys_tmp5282;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub27_result_datain <= w_sys_tmp6890;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub27_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'he)) begin
										r_sub27_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hf)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub27_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub27_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h5f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp1519[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h5f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_T_datain <= w_sys_tmp1522;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h5f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub08_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h5f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp1511[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h5f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_U_datain <= w_sys_tmp1514;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h5f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub08_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp5093[11:0] );

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp5084[11:0] );

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp5340[11:0] );

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp5345[11:0] );

									end
									else
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp5369[11:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp5355[11:0] );

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp10092[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub08_result_datain <= w_sys_tmp5086;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub08_result_datain <= w_sys_tmp5387;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub08_result_datain <= w_sys_tmp5349;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub08_result_datain <= r_sys_tmp5_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub08_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h3)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub08_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub08_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub24_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp3845[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub24_T_datain <= w_sys_tmp3848;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub24_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub24_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp3837[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub24_U_datain <= w_sys_tmp3840;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub24_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub24_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp5252[11:0] );

									end
									else
									if((r_sys_run_step==6'h3)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp5261[11:0] );

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp5378[11:0] );

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp5383[11:0] );

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp11596[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub24_result_datain <= w_sys_tmp5254;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub24_result_datain <= w_sys_tmp5387;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub24_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h3)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub24_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub24_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub25_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub25_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub25_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hcf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub25_T_addr <= $signed( w_sys_tmp3990[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hcf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub25_T_datain <= w_sys_tmp3993;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub25_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hcf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub25_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub25_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub25_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hcf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub25_U_addr <= $signed( w_sys_tmp3982[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hcf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub25_U_datain <= w_sys_tmp3985;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub25_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hcf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub25_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub25_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub25_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5)) begin
										r_sub25_result_addr <= $signed( w_sys_tmp5258[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_addr <= $signed( w_sys_tmp5255[11:0] );

									end
									else
									if((r_sys_run_step==6'h7)) begin
										r_sub25_result_addr <= $signed( w_sys_tmp5252[11:0] );

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub25_result_addr <= $signed( w_sys_tmp5264[11:0] );

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub25_result_addr <= $signed( w_sys_tmp5879[11:0] );

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub25_result_addr <= $signed( w_sys_tmp5884[11:0] );

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub25_result_addr <= $signed( w_sys_tmp11673[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5)) begin
										r_sub25_result_datain <= w_sys_tmp5260;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub25_result_datain <= r_sys_tmp5_float;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub25_result_datain <= w_sys_tmp5888;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub25_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6)) begin
										r_sub25_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub25_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub25_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub22_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp3552[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub22_T_datain <= w_sys_tmp3555;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub22_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub22_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp3544[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub22_U_datain <= w_sys_tmp3547;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub22_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub22_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1b)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp5168[11:0] );

									end
									else
									if((r_sys_run_step==6'h1a)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp5180[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp5171[11:0] );

									end
									else
									if((r_sys_run_step==6'h19)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp5174[11:0] );

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp8380[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp8365[11:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp8370[11:0] );

									end
									else
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp8394[11:0] );

									end
								end

							endcase
						end

						10'h1dc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp11401[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1a)) begin
										r_sub22_result_datain <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==6'h19)) begin
										r_sub22_result_datain <= w_sys_tmp5231;

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub22_result_datain <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub22_result_datain <= w_sys_tmp8345;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a)) begin
										r_sub22_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1b)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub22_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h1dc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub22_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub23_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hbe: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp3697[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hbe: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub23_T_datain <= w_sys_tmp3700;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hbe: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub23_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub23_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hbe: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp3689[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hbe: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub23_U_datain <= w_sys_tmp3692;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hbe: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub23_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub23_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp5171[11:0] );

									end
									else
									if((r_sys_run_step==6'h1d)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp5174[11:0] );

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp8866[11:0] );

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp8881[11:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp8871[11:0] );

									end
								end

							endcase
						end

						10'h1e2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp11497[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sub23_result_datain <= w_sys_tmp5242;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h2a)) begin
										r_sub23_result_datain <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'h3a)) begin
										r_sub23_result_datain <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==6'h22)) begin
										r_sub23_result_datain <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==6'h12)) begin
										r_sub23_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h32)) begin
										r_sub23_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub23_result_datain <= w_sys_tmp8846;

									end
									else
									if((r_sys_run_step==6'h1a)) begin
										r_sub23_result_datain <= r_sys_tmp3_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sub23_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub23_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h1e2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub23_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h3c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp791[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h3c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_T_datain <= w_sys_tmp794;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h3c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub03_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h3c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp783[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h3c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_U_datain <= w_sys_tmp786;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h3c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub03_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp5006[11:0] );

									end
									else
									if((r_sys_run_step==6'he)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp5012[11:0] );

									end
									else
									if((r_sys_run_step==6'hf)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp5000[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp5003[11:0] );

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp6838[11:0] );

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp6853[11:0] );

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp9609[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub03_result_datain <= w_sys_tmp5030;

									end
									else
									if((r_sys_run_step==6'he)) begin
										r_sub03_result_datain <= r_sys_tmp5_float;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub03_result_datain <= w_sys_tmp6842;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'he)) begin
										r_sub03_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hf)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub03_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub03_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h36: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp646[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h36: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_T_datain <= w_sys_tmp649;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h36: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub02_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h36: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp638[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h36: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_U_datain <= w_sys_tmp641;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h36: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub02_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp5006[11:0] );

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp5012[11:0] );

									end
									else
									if((r_sys_run_step==6'hb)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp5000[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp5003[11:0] );

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp6337[11:0] );

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp6352[11:0] );

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp9513[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha)) begin
										r_sub02_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_sub02_result_datain <= w_sys_tmp5002;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub02_result_datain <= w_sys_tmp6341;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha)) begin
										r_sub02_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub02_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub02_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h30: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp501[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h30: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_T_datain <= w_sys_tmp504;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h30: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub01_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h30: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp493[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h30: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_U_datain <= w_sys_tmp496;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h30: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub01_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp5006[11:0] );

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp5012[11:0] );

									end
									else
									if((r_sys_run_step==6'h7)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp5000[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp5003[11:0] );

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp5851[11:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp5836[11:0] );

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp9417[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub01_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub01_result_datain <= w_sys_tmp5008;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub01_result_datain <= w_sys_tmp5840;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6)) begin
										r_sub01_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub01_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp356[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_T_datain <= w_sys_tmp359;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub00_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp348[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_U_datain <= w_sys_tmp351;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub00_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp5000[11:0] );

									end
									else
									if((r_sys_run_step==6'h3)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp5009[11:0] );

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp5350[11:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp5335[11:0] );

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp9340[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub00_result_datain <= w_sys_tmp5002;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub00_result_datain <= w_sys_tmp5339;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub00_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h3)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub00_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub07_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h54: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp1371[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h54: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_T_datain <= w_sys_tmp1374;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h54: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub07_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h54: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp1363[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h54: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_U_datain <= w_sys_tmp1366;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h54: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub07_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp5006[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp5003[11:0] );

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp8857[11:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp8842[11:0] );

									end
								end

							endcase
						end

						10'h178: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp9993[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sub07_result_datain <= w_sys_tmp5074;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub07_result_datain <= w_sys_tmp8846;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sub07_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub07_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h178: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub07_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub06_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp1226[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_T_datain <= w_sys_tmp1229;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub06_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp1218[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_U_datain <= w_sys_tmp1221;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub06_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h19)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp5006[11:0] );

									end
									else
									if((r_sys_run_step==6'h1a)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp5012[11:0] );

									end
									else
									if((r_sys_run_step==6'h1b)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp5000[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp5003[11:0] );

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp8356[11:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp8341[11:0] );

									end
								end

							endcase
						end

						10'h172: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp9897[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1a)) begin
										r_sub06_result_datain <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==6'h19)) begin
										r_sub06_result_datain <= w_sys_tmp5063;

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub06_result_datain <= w_sys_tmp8345;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a)) begin
										r_sub06_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1b)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub06_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h172: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub06_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub05_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h48: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp1081[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h48: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_T_datain <= w_sys_tmp1084;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h48: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub05_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h48: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp1073[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h48: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_U_datain <= w_sys_tmp1076;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h48: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub05_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h15)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp5006[11:0] );

									end
									else
									if((r_sys_run_step==6'h16)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp5012[11:0] );

									end
									else
									if((r_sys_run_step==6'h17)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp5000[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp5003[11:0] );

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp7840[11:0] );

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp7855[11:0] );

									end
								end

							endcase
						end

						10'h16c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp9801[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h16)) begin
										r_sub05_result_datain <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'h15)) begin
										r_sub05_result_datain <= w_sys_tmp5052;

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub05_result_datain <= w_sys_tmp7844;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h15) || (r_sys_run_step==6'h16)) begin
										r_sub05_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h17)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub05_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h16c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub05_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub04_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h42: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp936[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h42: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_T_datain <= w_sys_tmp939;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h42: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub04_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h42: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp928[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h42: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_U_datain <= w_sys_tmp931;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h42: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub04_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h11)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp5006[11:0] );

									end
									else
									if((r_sys_run_step==6'h12)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp5012[11:0] );

									end
									else
									if((r_sys_run_step==6'h13)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp5000[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp5003[11:0] );

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp7354[11:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp7339[11:0] );

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp9705[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h12)) begin
										r_sub04_result_datain <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==6'h11)) begin
										r_sub04_result_datain <= w_sys_tmp5041;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub04_result_datain <= w_sys_tmp7343;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h11) || (r_sys_run_step==6'h12)) begin
										r_sub04_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h13)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub04_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub04_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub10_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h6b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp1809[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h6b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_T_datain <= w_sys_tmp1812;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h6b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub10_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h6b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp1801[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h6b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_U_datain <= w_sys_tmp1804;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h6b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub10_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5096[11:0] );

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5090[11:0] );

									end
									else
									if((r_sys_run_step==6'hb)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5084[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5087[11:0] );

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp6371[11:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp6357[11:0] );

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp6347[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp6342[11:0] );

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp10265[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha)) begin
										r_sub10_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_sub10_result_datain <= w_sys_tmp5086;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub10_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub10_result_datain <= w_sys_tmp6389;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub10_result_datain <= w_sys_tmp6351;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha)) begin
										r_sub10_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub10_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub10_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub31_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub31_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub31_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub31_T_addr <= $signed( w_sys_tmp4860[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub31_T_datain <= w_sys_tmp4863;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub31_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub31_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub31_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub31_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub31_U_addr <= $signed( w_sys_tmp4852[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub31_U_datain <= w_sys_tmp4855;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub31_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub31_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub31_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub31_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sub31_result_addr <= $signed( w_sys_tmp5258[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_addr <= $signed( w_sys_tmp5255[11:0] );

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h3) || (r_sys_run_step==6'h5) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h9) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hd)) begin
										r_sub31_result_addr <= $signed( w_sys_tmp8885[11:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h4) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'he)) begin
										r_sub31_result_addr <= $signed( w_sys_tmp8890[11:0] );

									end
								end

							endcase
						end

						10'h217: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub31_result_addr <= $signed( w_sys_tmp12249[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sub31_result_datain <= w_sys_tmp5326;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h4) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'ha)) begin
										r_sub31_result_datain <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==6'hc)) begin
										r_sub31_result_datain <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub31_result_datain <= w_sys_tmp8894;

									end
									else
									if((r_sys_run_step==6'h8) || (r_sys_run_step==6'he)) begin
										r_sub31_result_datain <= r_sys_tmp5_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub31_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sub31_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h4) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'he)) begin
										r_sub31_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h3) || (r_sys_run_step==6'h5) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h9) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hd)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h217: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub31_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub30_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub30_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub30_T_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub30_T_addr <= $signed( w_sys_tmp4715[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub30_T_datain <= w_sys_tmp4718;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub30_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub30_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub30_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub30_U_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub30_U_addr <= $signed( w_sys_tmp4707[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub30_U_datain <= w_sys_tmp4710;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub30_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub30_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub30_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub30_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h19)) begin
										r_sub30_result_addr <= $signed( w_sys_tmp5258[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_addr <= $signed( w_sys_tmp5255[11:0] );

									end
									else
									if((r_sys_run_step==6'h1b)) begin
										r_sub30_result_addr <= $signed( w_sys_tmp5252[11:0] );

									end
									else
									if((r_sys_run_step==6'h1a)) begin
										r_sub30_result_addr <= $signed( w_sys_tmp5264[11:0] );

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub30_result_addr <= $signed( w_sys_tmp8389[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub30_result_addr <= $signed( w_sys_tmp8384[11:0] );

									end
								end

							endcase
						end

						10'h211: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub30_result_addr <= $signed( w_sys_tmp12153[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1a)) begin
										r_sub30_result_datain <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==6'h19)) begin
										r_sub30_result_datain <= w_sys_tmp5315;

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub30_result_datain <= w_sys_tmp8393;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub30_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a)) begin
										r_sub30_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1b)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub30_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h211: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h21b: begin
							r_sub30_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h16)) begin
										r_sys_tmp0_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_sub27_result_dataout;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp0_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp0_float <= w_sub28_result_dataout;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5)) begin
										r_sys_tmp0_float <= w_sub31_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h16)) begin
										r_sys_tmp1_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub29_result_dataout;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub20_result_dataout;

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_tmp1_float <= w_sub31_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h12) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h19)) begin
										r_sys_tmp2_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp2_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp2_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp2_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp2_float <= w_sub31_result_dataout;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp2_float <= w_sub26_result_dataout;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9)) begin
										r_sys_tmp2_float <= w_sub31_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h11) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h17)) begin
										r_sys_tmp3_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp3_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp3_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp3_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp3_float <= w_sub30_result_dataout;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp3_float <= w_sub27_result_dataout;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h7)) begin
										r_sys_tmp3_float <= w_sub31_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hc) || (r_sys_run_step==6'hd)) begin
										r_sys_tmp4_float <= w_ip_FixedToFloat_floating_0;

									end
									else
									if((r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h19)) begin
										r_sys_tmp4_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp4_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp4_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp4_float <= w_sub20_result_dataout;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp4_float <= w_sub28_result_dataout;

									end
								end

							endcase
						end

						10'h13d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp4_float <= w_sub30_result_dataout;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'hb)) begin
										r_sys_tmp4_float <= w_sub31_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp5_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp5_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp5_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp5_float <= w_sub26_result_dataout;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp5_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp5_float <= w_sub25_result_dataout;

									end
								end

							endcase
						end

						10'h137: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp5_float <= w_sub29_result_dataout;

									end
								end

							endcase
						end

						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h8)) begin
										r_sys_tmp5_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hf)) begin
										r_sys_tmp6_float <= w_sub31_result_dataout;

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h4) || (r_sys_run_step==6'h6)) begin
										r_sys_tmp6_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

						10'h219: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp6_float <= w_sys_tmp12333;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h143: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sys_tmp7_float <= w_sub23_result_dataout;

									end
									else
									if((r_sys_run_step==6'h7)) begin
										r_sys_tmp7_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
