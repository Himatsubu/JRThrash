/*
TimeStamp:	2016/9/29		13:0
*/


module c1(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy	
);

	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 7:0] r_sys_run_phase;
	reg         [ 4:0] r_sys_run_stage;
	reg         [ 8:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 4:0] w_sys_run_stage_p1;
	wire        [ 8:0] w_sys_run_step_p1;
	wire signed [14:0] w_fld_u_0_addr_0;
	wire        [31:0] w_fld_u_0_datain_0;
	wire        [31:0] w_fld_u_0_dataout_0;
	wire               w_fld_u_0_r_w_0;
	wire               w_fld_u_0_ce_0;
	reg  signed [14:0] r_fld_u_0_addr_1;
	reg         [31:0] r_fld_u_0_datain_1;
	wire        [31:0] w_fld_u_0_dataout_1;
	reg                r_fld_u_0_r_w_1;
	wire               w_fld_u_0_ce_1;
	reg  signed [31:0] r_run_k_17;
	reg  signed [31:0] r_run_j_18;
	reg  signed [31:0] r_run_n_19;
	reg  signed [31:0] r_run_mx_20;
	reg  signed [31:0] r_run_my_21;
	reg  signed [31:0] r_run_nlast_22;
	reg  signed [31:0] r_run_copy0_j_23;
	reg  signed [31:0] r_run_copy1_j_24;
	reg  signed [31:0] r_run_copy2_j_25;
	reg  signed [31:0] r_run_copy0_j_26;
	reg  signed [31:0] r_run_copy0_j_27;
	reg  signed [31:0] r_run_copy0_j_28;
	reg  signed [31:0] r_run_copy0_j_29;
	reg  signed [31:0] r_run_copy0_j_30;
	reg  signed [31:0] r_run_copy0_j_31;
	reg  signed [31:0] r_run_copy0_j_32;
	reg  signed [31:0] r_run_copy0_j_33;
	reg  signed [31:0] r_run_copy0_j_34;
	reg  signed [31:0] r_run_copy0_j_35;
	reg  signed [31:0] r_run_copy0_j_36;
	reg  signed [31:0] r_run_copy0_j_37;
	reg  signed [31:0] r_run_copy0_j_38;
	reg  signed [31:0] r_run_copy0_j_39;
	reg  signed [31:0] r_run_copy0_j_40;
	reg  signed [31:0] r_run_copy0_j_41;
	reg                r_sub09_run_req;
	wire               w_sub09_run_busy;
	wire signed [12:0] w_sub09_u_addr;
	reg  signed [12:0] r_sub09_u_addr;
	wire        [31:0] w_sub09_u_datain;
	reg         [31:0] r_sub09_u_datain;
	wire        [31:0] w_sub09_u_dataout;
	wire               w_sub09_u_r_w;
	reg                r_sub09_u_r_w;
	wire signed [12:0] w_sub09_result_addr;
	reg  signed [12:0] r_sub09_result_addr;
	wire        [31:0] w_sub09_result_datain;
	reg         [31:0] r_sub09_result_datain;
	wire        [31:0] w_sub09_result_dataout;
	wire               w_sub09_result_r_w;
	reg                r_sub09_result_r_w;
	reg                r_sub08_run_req;
	wire               w_sub08_run_busy;
	wire signed [12:0] w_sub08_u_addr;
	reg  signed [12:0] r_sub08_u_addr;
	wire        [31:0] w_sub08_u_datain;
	reg         [31:0] r_sub08_u_datain;
	wire        [31:0] w_sub08_u_dataout;
	wire               w_sub08_u_r_w;
	reg                r_sub08_u_r_w;
	wire signed [12:0] w_sub08_result_addr;
	reg  signed [12:0] r_sub08_result_addr;
	wire        [31:0] w_sub08_result_datain;
	reg         [31:0] r_sub08_result_datain;
	wire        [31:0] w_sub08_result_dataout;
	wire               w_sub08_result_r_w;
	reg                r_sub08_result_r_w;
	reg                r_sub12_run_req;
	wire               w_sub12_run_busy;
	wire signed [12:0] w_sub12_u_addr;
	reg  signed [12:0] r_sub12_u_addr;
	wire        [31:0] w_sub12_u_datain;
	reg         [31:0] r_sub12_u_datain;
	wire        [31:0] w_sub12_u_dataout;
	wire               w_sub12_u_r_w;
	reg                r_sub12_u_r_w;
	wire signed [12:0] w_sub12_result_addr;
	reg  signed [12:0] r_sub12_result_addr;
	wire        [31:0] w_sub12_result_datain;
	reg         [31:0] r_sub12_result_datain;
	wire        [31:0] w_sub12_result_dataout;
	wire               w_sub12_result_r_w;
	reg                r_sub12_result_r_w;
	reg                r_sub03_run_req;
	wire               w_sub03_run_busy;
	wire signed [12:0] w_sub03_u_addr;
	reg  signed [12:0] r_sub03_u_addr;
	wire        [31:0] w_sub03_u_datain;
	reg         [31:0] r_sub03_u_datain;
	wire        [31:0] w_sub03_u_dataout;
	wire               w_sub03_u_r_w;
	reg                r_sub03_u_r_w;
	wire signed [12:0] w_sub03_result_addr;
	reg  signed [12:0] r_sub03_result_addr;
	wire        [31:0] w_sub03_result_datain;
	reg         [31:0] r_sub03_result_datain;
	wire        [31:0] w_sub03_result_dataout;
	wire               w_sub03_result_r_w;
	reg                r_sub03_result_r_w;
	reg                r_sub02_run_req;
	wire               w_sub02_run_busy;
	wire signed [12:0] w_sub02_u_addr;
	reg  signed [12:0] r_sub02_u_addr;
	wire        [31:0] w_sub02_u_datain;
	reg         [31:0] r_sub02_u_datain;
	wire        [31:0] w_sub02_u_dataout;
	wire               w_sub02_u_r_w;
	reg                r_sub02_u_r_w;
	wire signed [12:0] w_sub02_result_addr;
	reg  signed [12:0] r_sub02_result_addr;
	wire        [31:0] w_sub02_result_datain;
	reg         [31:0] r_sub02_result_datain;
	wire        [31:0] w_sub02_result_dataout;
	wire               w_sub02_result_r_w;
	reg                r_sub02_result_r_w;
	reg                r_sub11_run_req;
	wire               w_sub11_run_busy;
	wire signed [12:0] w_sub11_u_addr;
	reg  signed [12:0] r_sub11_u_addr;
	wire        [31:0] w_sub11_u_datain;
	reg         [31:0] r_sub11_u_datain;
	wire        [31:0] w_sub11_u_dataout;
	wire               w_sub11_u_r_w;
	reg                r_sub11_u_r_w;
	wire signed [12:0] w_sub11_result_addr;
	reg  signed [12:0] r_sub11_result_addr;
	wire        [31:0] w_sub11_result_datain;
	reg         [31:0] r_sub11_result_datain;
	wire        [31:0] w_sub11_result_dataout;
	wire               w_sub11_result_r_w;
	reg                r_sub11_result_r_w;
	reg                r_sub14_run_req;
	wire               w_sub14_run_busy;
	wire signed [12:0] w_sub14_u_addr;
	reg  signed [12:0] r_sub14_u_addr;
	wire        [31:0] w_sub14_u_datain;
	reg         [31:0] r_sub14_u_datain;
	wire        [31:0] w_sub14_u_dataout;
	wire               w_sub14_u_r_w;
	reg                r_sub14_u_r_w;
	wire signed [12:0] w_sub14_result_addr;
	reg  signed [12:0] r_sub14_result_addr;
	wire        [31:0] w_sub14_result_datain;
	reg         [31:0] r_sub14_result_datain;
	wire        [31:0] w_sub14_result_dataout;
	wire               w_sub14_result_r_w;
	reg                r_sub14_result_r_w;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [12:0] w_sub01_u_addr;
	reg  signed [12:0] r_sub01_u_addr;
	wire        [31:0] w_sub01_u_datain;
	reg         [31:0] r_sub01_u_datain;
	wire        [31:0] w_sub01_u_dataout;
	wire               w_sub01_u_r_w;
	reg                r_sub01_u_r_w;
	wire signed [12:0] w_sub01_result_addr;
	reg  signed [12:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub13_run_req;
	wire               w_sub13_run_busy;
	wire signed [12:0] w_sub13_u_addr;
	reg  signed [12:0] r_sub13_u_addr;
	wire        [31:0] w_sub13_u_datain;
	reg         [31:0] r_sub13_u_datain;
	wire        [31:0] w_sub13_u_dataout;
	wire               w_sub13_u_r_w;
	reg                r_sub13_u_r_w;
	wire signed [12:0] w_sub13_result_addr;
	reg  signed [12:0] r_sub13_result_addr;
	wire        [31:0] w_sub13_result_datain;
	reg         [31:0] r_sub13_result_datain;
	wire        [31:0] w_sub13_result_dataout;
	wire               w_sub13_result_r_w;
	reg                r_sub13_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [12:0] w_sub00_u_addr;
	reg  signed [12:0] r_sub00_u_addr;
	wire        [31:0] w_sub00_u_datain;
	reg         [31:0] r_sub00_u_datain;
	wire        [31:0] w_sub00_u_dataout;
	wire               w_sub00_u_r_w;
	reg                r_sub00_u_r_w;
	wire signed [12:0] w_sub00_result_addr;
	reg  signed [12:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	reg                r_sub07_run_req;
	wire               w_sub07_run_busy;
	wire signed [12:0] w_sub07_u_addr;
	reg  signed [12:0] r_sub07_u_addr;
	wire        [31:0] w_sub07_u_datain;
	reg         [31:0] r_sub07_u_datain;
	wire        [31:0] w_sub07_u_dataout;
	wire               w_sub07_u_r_w;
	reg                r_sub07_u_r_w;
	wire signed [12:0] w_sub07_result_addr;
	reg  signed [12:0] r_sub07_result_addr;
	wire        [31:0] w_sub07_result_datain;
	reg         [31:0] r_sub07_result_datain;
	wire        [31:0] w_sub07_result_dataout;
	wire               w_sub07_result_r_w;
	reg                r_sub07_result_r_w;
	reg                r_sub06_run_req;
	wire               w_sub06_run_busy;
	wire signed [12:0] w_sub06_u_addr;
	reg  signed [12:0] r_sub06_u_addr;
	wire        [31:0] w_sub06_u_datain;
	reg         [31:0] r_sub06_u_datain;
	wire        [31:0] w_sub06_u_dataout;
	wire               w_sub06_u_r_w;
	reg                r_sub06_u_r_w;
	wire signed [12:0] w_sub06_result_addr;
	reg  signed [12:0] r_sub06_result_addr;
	wire        [31:0] w_sub06_result_datain;
	reg         [31:0] r_sub06_result_datain;
	wire        [31:0] w_sub06_result_dataout;
	wire               w_sub06_result_r_w;
	reg                r_sub06_result_r_w;
	reg                r_sub15_run_req;
	wire               w_sub15_run_busy;
	wire signed [12:0] w_sub15_u_addr;
	reg  signed [12:0] r_sub15_u_addr;
	wire        [31:0] w_sub15_u_datain;
	reg         [31:0] r_sub15_u_datain;
	wire        [31:0] w_sub15_u_dataout;
	wire               w_sub15_u_r_w;
	reg                r_sub15_u_r_w;
	wire signed [12:0] w_sub15_result_addr;
	reg  signed [12:0] r_sub15_result_addr;
	wire        [31:0] w_sub15_result_datain;
	reg         [31:0] r_sub15_result_datain;
	wire        [31:0] w_sub15_result_dataout;
	wire               w_sub15_result_r_w;
	reg                r_sub15_result_r_w;
	reg                r_sub05_run_req;
	wire               w_sub05_run_busy;
	wire signed [12:0] w_sub05_u_addr;
	reg  signed [12:0] r_sub05_u_addr;
	wire        [31:0] w_sub05_u_datain;
	reg         [31:0] r_sub05_u_datain;
	wire        [31:0] w_sub05_u_dataout;
	wire               w_sub05_u_r_w;
	reg                r_sub05_u_r_w;
	wire signed [12:0] w_sub05_result_addr;
	reg  signed [12:0] r_sub05_result_addr;
	wire        [31:0] w_sub05_result_datain;
	reg         [31:0] r_sub05_result_datain;
	wire        [31:0] w_sub05_result_dataout;
	wire               w_sub05_result_r_w;
	reg                r_sub05_result_r_w;
	reg                r_sub04_run_req;
	wire               w_sub04_run_busy;
	wire signed [12:0] w_sub04_u_addr;
	reg  signed [12:0] r_sub04_u_addr;
	wire        [31:0] w_sub04_u_datain;
	reg         [31:0] r_sub04_u_datain;
	wire        [31:0] w_sub04_u_dataout;
	wire               w_sub04_u_r_w;
	reg                r_sub04_u_r_w;
	wire signed [12:0] w_sub04_result_addr;
	reg  signed [12:0] r_sub04_result_addr;
	wire        [31:0] w_sub04_result_datain;
	reg         [31:0] r_sub04_result_datain;
	wire        [31:0] w_sub04_result_dataout;
	wire               w_sub04_result_r_w;
	reg                r_sub04_result_r_w;
	reg                r_sub10_run_req;
	wire               w_sub10_run_busy;
	wire signed [12:0] w_sub10_u_addr;
	reg  signed [12:0] r_sub10_u_addr;
	wire        [31:0] w_sub10_u_datain;
	reg         [31:0] r_sub10_u_datain;
	wire        [31:0] w_sub10_u_dataout;
	wire               w_sub10_u_r_w;
	reg                r_sub10_u_r_w;
	wire signed [12:0] w_sub10_result_addr;
	reg  signed [12:0] r_sub10_result_addr;
	wire        [31:0] w_sub10_result_datain;
	reg         [31:0] r_sub10_result_datain;
	wire        [31:0] w_sub10_result_dataout;
	wire               w_sub10_result_r_w;
	reg                r_sub10_result_r_w;
	wire signed [31:0] w_sys_tmp1;
	wire               w_sys_tmp3;
	wire               w_sys_tmp4;
	wire signed [31:0] w_sys_tmp5;
	wire               w_sys_tmp6;
	wire               w_sys_tmp7;
	wire signed [31:0] w_sys_tmp10;
	wire signed [31:0] w_sys_tmp11;
	wire signed [31:0] w_sys_tmp12;
	wire        [31:0] w_sys_tmp13;
	wire signed [31:0] w_sys_tmp14;
	wire               w_sys_tmp51;
	wire               w_sys_tmp52;
	wire signed [31:0] w_sys_tmp53;
	wire               w_sys_tmp54;
	wire               w_sys_tmp55;
	wire signed [31:0] w_sys_tmp58;
	wire signed [31:0] w_sys_tmp59;
	wire        [31:0] w_sys_tmp60;
	wire signed [31:0] w_sys_tmp62;
	wire signed [31:0] w_sys_tmp63;
	wire        [31:0] w_sys_tmp64;
	wire signed [31:0] w_sys_tmp66;
	wire signed [31:0] w_sys_tmp67;
	wire        [31:0] w_sys_tmp69;
	wire signed [31:0] w_sys_tmp71;
	wire signed [31:0] w_sys_tmp72;
	wire signed [31:0] w_sys_tmp75;
	wire signed [31:0] w_sys_tmp76;
	wire signed [31:0] w_sys_tmp77;
	wire signed [31:0] w_sys_tmp78;
	wire               w_sys_tmp211;
	wire               w_sys_tmp212;
	wire signed [31:0] w_sys_tmp213;
	wire signed [31:0] w_sys_tmp216;
	wire signed [31:0] w_sys_tmp217;
	wire        [31:0] w_sys_tmp218;
	wire signed [31:0] w_sys_tmp222;
	wire signed [31:0] w_sys_tmp223;
	wire signed [31:0] w_sys_tmp228;
	wire signed [31:0] w_sys_tmp229;
	wire signed [31:0] w_sys_tmp234;
	wire signed [31:0] w_sys_tmp235;
	wire signed [31:0] w_sys_tmp240;
	wire signed [31:0] w_sys_tmp241;
	wire signed [31:0] w_sys_tmp246;
	wire signed [31:0] w_sys_tmp247;
	wire signed [31:0] w_sys_tmp252;
	wire signed [31:0] w_sys_tmp253;
	wire signed [31:0] w_sys_tmp258;
	wire signed [31:0] w_sys_tmp259;
	wire signed [31:0] w_sys_tmp264;
	wire signed [31:0] w_sys_tmp265;
	wire signed [31:0] w_sys_tmp270;
	wire signed [31:0] w_sys_tmp271;
	wire signed [31:0] w_sys_tmp276;
	wire signed [31:0] w_sys_tmp277;
	wire signed [31:0] w_sys_tmp282;
	wire signed [31:0] w_sys_tmp283;
	wire signed [31:0] w_sys_tmp288;
	wire signed [31:0] w_sys_tmp289;
	wire signed [31:0] w_sys_tmp294;
	wire signed [31:0] w_sys_tmp295;
	wire signed [31:0] w_sys_tmp300;
	wire signed [31:0] w_sys_tmp301;
	wire signed [31:0] w_sys_tmp306;
	wire signed [31:0] w_sys_tmp307;
	wire signed [31:0] w_sys_tmp312;
	wire signed [31:0] w_sys_tmp313;
	wire signed [31:0] w_sys_tmp318;
	wire signed [31:0] w_sys_tmp319;
	wire signed [31:0] w_sys_tmp324;
	wire signed [31:0] w_sys_tmp325;
	wire signed [31:0] w_sys_tmp330;
	wire signed [31:0] w_sys_tmp331;
	wire signed [31:0] w_sys_tmp336;
	wire signed [31:0] w_sys_tmp337;
	wire signed [31:0] w_sys_tmp342;
	wire signed [31:0] w_sys_tmp343;
	wire signed [31:0] w_sys_tmp348;
	wire signed [31:0] w_sys_tmp349;
	wire signed [31:0] w_sys_tmp354;
	wire signed [31:0] w_sys_tmp355;
	wire signed [31:0] w_sys_tmp360;
	wire signed [31:0] w_sys_tmp361;
	wire signed [31:0] w_sys_tmp366;
	wire signed [31:0] w_sys_tmp367;
	wire signed [31:0] w_sys_tmp372;
	wire signed [31:0] w_sys_tmp373;
	wire signed [31:0] w_sys_tmp378;
	wire signed [31:0] w_sys_tmp379;
	wire signed [31:0] w_sys_tmp384;
	wire signed [31:0] w_sys_tmp385;
	wire signed [31:0] w_sys_tmp390;
	wire signed [31:0] w_sys_tmp391;
	wire signed [31:0] w_sys_tmp396;
	wire signed [31:0] w_sys_tmp397;
	wire signed [31:0] w_sys_tmp402;
	wire signed [31:0] w_sys_tmp403;
	wire signed [31:0] w_sys_tmp408;
	wire signed [31:0] w_sys_tmp409;
	wire signed [31:0] w_sys_tmp429;
	wire signed [31:0] w_sys_tmp430;
	wire signed [31:0] w_sys_tmp435;
	wire signed [31:0] w_sys_tmp436;
	wire signed [31:0] w_sys_tmp441;
	wire signed [31:0] w_sys_tmp442;
	wire signed [31:0] w_sys_tmp447;
	wire signed [31:0] w_sys_tmp448;
	wire signed [31:0] w_sys_tmp453;
	wire signed [31:0] w_sys_tmp454;
	wire signed [31:0] w_sys_tmp459;
	wire signed [31:0] w_sys_tmp460;
	wire signed [31:0] w_sys_tmp465;
	wire signed [31:0] w_sys_tmp466;
	wire signed [31:0] w_sys_tmp471;
	wire signed [31:0] w_sys_tmp472;
	wire signed [31:0] w_sys_tmp477;
	wire signed [31:0] w_sys_tmp478;
	wire signed [31:0] w_sys_tmp483;
	wire signed [31:0] w_sys_tmp484;
	wire signed [31:0] w_sys_tmp489;
	wire signed [31:0] w_sys_tmp490;
	wire signed [31:0] w_sys_tmp495;
	wire signed [31:0] w_sys_tmp496;
	wire signed [31:0] w_sys_tmp501;
	wire signed [31:0] w_sys_tmp502;
	wire signed [31:0] w_sys_tmp507;
	wire signed [31:0] w_sys_tmp508;
	wire signed [31:0] w_sys_tmp513;
	wire signed [31:0] w_sys_tmp514;
	wire signed [31:0] w_sys_tmp519;
	wire signed [31:0] w_sys_tmp520;
	wire signed [31:0] w_sys_tmp525;
	wire signed [31:0] w_sys_tmp526;
	wire signed [31:0] w_sys_tmp531;
	wire signed [31:0] w_sys_tmp532;
	wire signed [31:0] w_sys_tmp537;
	wire signed [31:0] w_sys_tmp538;
	wire signed [31:0] w_sys_tmp543;
	wire signed [31:0] w_sys_tmp544;
	wire signed [31:0] w_sys_tmp549;
	wire signed [31:0] w_sys_tmp550;
	wire signed [31:0] w_sys_tmp555;
	wire signed [31:0] w_sys_tmp556;
	wire signed [31:0] w_sys_tmp561;
	wire signed [31:0] w_sys_tmp562;
	wire signed [31:0] w_sys_tmp567;
	wire signed [31:0] w_sys_tmp568;
	wire signed [31:0] w_sys_tmp573;
	wire signed [31:0] w_sys_tmp574;
	wire signed [31:0] w_sys_tmp579;
	wire signed [31:0] w_sys_tmp580;
	wire signed [31:0] w_sys_tmp585;
	wire signed [31:0] w_sys_tmp586;
	wire signed [31:0] w_sys_tmp591;
	wire signed [31:0] w_sys_tmp592;
	wire signed [31:0] w_sys_tmp597;
	wire signed [31:0] w_sys_tmp598;
	wire signed [31:0] w_sys_tmp603;
	wire signed [31:0] w_sys_tmp604;
	wire signed [31:0] w_sys_tmp609;
	wire signed [31:0] w_sys_tmp610;
	wire signed [31:0] w_sys_tmp615;
	wire signed [31:0] w_sys_tmp616;
	wire signed [31:0] w_sys_tmp633;
	wire signed [31:0] w_sys_tmp634;
	wire signed [31:0] w_sys_tmp639;
	wire signed [31:0] w_sys_tmp640;
	wire signed [31:0] w_sys_tmp645;
	wire signed [31:0] w_sys_tmp646;
	wire signed [31:0] w_sys_tmp651;
	wire signed [31:0] w_sys_tmp652;
	wire signed [31:0] w_sys_tmp657;
	wire signed [31:0] w_sys_tmp658;
	wire signed [31:0] w_sys_tmp663;
	wire signed [31:0] w_sys_tmp664;
	wire signed [31:0] w_sys_tmp669;
	wire signed [31:0] w_sys_tmp670;
	wire signed [31:0] w_sys_tmp675;
	wire signed [31:0] w_sys_tmp676;
	wire signed [31:0] w_sys_tmp681;
	wire signed [31:0] w_sys_tmp682;
	wire signed [31:0] w_sys_tmp687;
	wire signed [31:0] w_sys_tmp688;
	wire signed [31:0] w_sys_tmp693;
	wire signed [31:0] w_sys_tmp694;
	wire signed [31:0] w_sys_tmp699;
	wire signed [31:0] w_sys_tmp700;
	wire signed [31:0] w_sys_tmp705;
	wire signed [31:0] w_sys_tmp706;
	wire signed [31:0] w_sys_tmp711;
	wire signed [31:0] w_sys_tmp712;
	wire signed [31:0] w_sys_tmp717;
	wire signed [31:0] w_sys_tmp718;
	wire signed [31:0] w_sys_tmp723;
	wire signed [31:0] w_sys_tmp724;
	wire signed [31:0] w_sys_tmp729;
	wire signed [31:0] w_sys_tmp730;
	wire signed [31:0] w_sys_tmp735;
	wire signed [31:0] w_sys_tmp736;
	wire signed [31:0] w_sys_tmp741;
	wire signed [31:0] w_sys_tmp742;
	wire signed [31:0] w_sys_tmp747;
	wire signed [31:0] w_sys_tmp748;
	wire signed [31:0] w_sys_tmp753;
	wire signed [31:0] w_sys_tmp754;
	wire signed [31:0] w_sys_tmp759;
	wire signed [31:0] w_sys_tmp760;
	wire signed [31:0] w_sys_tmp765;
	wire signed [31:0] w_sys_tmp766;
	wire signed [31:0] w_sys_tmp771;
	wire signed [31:0] w_sys_tmp772;
	wire signed [31:0] w_sys_tmp777;
	wire signed [31:0] w_sys_tmp778;
	wire signed [31:0] w_sys_tmp783;
	wire signed [31:0] w_sys_tmp784;
	wire signed [31:0] w_sys_tmp789;
	wire signed [31:0] w_sys_tmp790;
	wire signed [31:0] w_sys_tmp795;
	wire signed [31:0] w_sys_tmp796;
	wire signed [31:0] w_sys_tmp801;
	wire signed [31:0] w_sys_tmp802;
	wire signed [31:0] w_sys_tmp807;
	wire signed [31:0] w_sys_tmp808;
	wire signed [31:0] w_sys_tmp813;
	wire signed [31:0] w_sys_tmp814;
	wire signed [31:0] w_sys_tmp819;
	wire signed [31:0] w_sys_tmp820;
	wire signed [31:0] w_sys_tmp837;
	wire signed [31:0] w_sys_tmp838;
	wire signed [31:0] w_sys_tmp843;
	wire signed [31:0] w_sys_tmp844;
	wire signed [31:0] w_sys_tmp849;
	wire signed [31:0] w_sys_tmp850;
	wire signed [31:0] w_sys_tmp855;
	wire signed [31:0] w_sys_tmp856;
	wire signed [31:0] w_sys_tmp861;
	wire signed [31:0] w_sys_tmp862;
	wire signed [31:0] w_sys_tmp867;
	wire signed [31:0] w_sys_tmp868;
	wire signed [31:0] w_sys_tmp873;
	wire signed [31:0] w_sys_tmp874;
	wire signed [31:0] w_sys_tmp879;
	wire signed [31:0] w_sys_tmp880;
	wire signed [31:0] w_sys_tmp885;
	wire signed [31:0] w_sys_tmp886;
	wire signed [31:0] w_sys_tmp891;
	wire signed [31:0] w_sys_tmp892;
	wire signed [31:0] w_sys_tmp897;
	wire signed [31:0] w_sys_tmp898;
	wire signed [31:0] w_sys_tmp903;
	wire signed [31:0] w_sys_tmp904;
	wire signed [31:0] w_sys_tmp909;
	wire signed [31:0] w_sys_tmp910;
	wire signed [31:0] w_sys_tmp915;
	wire signed [31:0] w_sys_tmp916;
	wire signed [31:0] w_sys_tmp921;
	wire signed [31:0] w_sys_tmp922;
	wire signed [31:0] w_sys_tmp927;
	wire signed [31:0] w_sys_tmp928;
	wire signed [31:0] w_sys_tmp933;
	wire signed [31:0] w_sys_tmp934;
	wire signed [31:0] w_sys_tmp939;
	wire signed [31:0] w_sys_tmp940;
	wire signed [31:0] w_sys_tmp945;
	wire signed [31:0] w_sys_tmp946;
	wire signed [31:0] w_sys_tmp951;
	wire signed [31:0] w_sys_tmp952;
	wire signed [31:0] w_sys_tmp957;
	wire signed [31:0] w_sys_tmp958;
	wire signed [31:0] w_sys_tmp963;
	wire signed [31:0] w_sys_tmp964;
	wire signed [31:0] w_sys_tmp969;
	wire signed [31:0] w_sys_tmp970;
	wire signed [31:0] w_sys_tmp975;
	wire signed [31:0] w_sys_tmp976;
	wire signed [31:0] w_sys_tmp981;
	wire signed [31:0] w_sys_tmp982;
	wire signed [31:0] w_sys_tmp987;
	wire signed [31:0] w_sys_tmp988;
	wire signed [31:0] w_sys_tmp993;
	wire signed [31:0] w_sys_tmp994;
	wire signed [31:0] w_sys_tmp999;
	wire signed [31:0] w_sys_tmp1000;
	wire signed [31:0] w_sys_tmp1005;
	wire signed [31:0] w_sys_tmp1006;
	wire signed [31:0] w_sys_tmp1011;
	wire signed [31:0] w_sys_tmp1012;
	wire signed [31:0] w_sys_tmp1017;
	wire signed [31:0] w_sys_tmp1018;
	wire signed [31:0] w_sys_tmp1023;
	wire signed [31:0] w_sys_tmp1024;
	wire signed [31:0] w_sys_tmp1025;
	wire signed [31:0] w_sys_tmp1026;
	wire               w_sys_tmp1027;
	wire               w_sys_tmp1028;
	wire signed [31:0] w_sys_tmp1029;
	wire signed [31:0] w_sys_tmp1032;
	wire signed [31:0] w_sys_tmp1033;
	wire        [31:0] w_sys_tmp1034;
	wire signed [31:0] w_sys_tmp1038;
	wire signed [31:0] w_sys_tmp1039;
	wire signed [31:0] w_sys_tmp1044;
	wire signed [31:0] w_sys_tmp1045;
	wire signed [31:0] w_sys_tmp1050;
	wire signed [31:0] w_sys_tmp1051;
	wire signed [31:0] w_sys_tmp1056;
	wire signed [31:0] w_sys_tmp1057;
	wire signed [31:0] w_sys_tmp1062;
	wire signed [31:0] w_sys_tmp1063;
	wire signed [31:0] w_sys_tmp1068;
	wire signed [31:0] w_sys_tmp1069;
	wire signed [31:0] w_sys_tmp1074;
	wire signed [31:0] w_sys_tmp1075;
	wire signed [31:0] w_sys_tmp1080;
	wire signed [31:0] w_sys_tmp1081;
	wire signed [31:0] w_sys_tmp1086;
	wire signed [31:0] w_sys_tmp1087;
	wire signed [31:0] w_sys_tmp1092;
	wire signed [31:0] w_sys_tmp1093;
	wire signed [31:0] w_sys_tmp1098;
	wire signed [31:0] w_sys_tmp1099;
	wire signed [31:0] w_sys_tmp1104;
	wire signed [31:0] w_sys_tmp1105;
	wire signed [31:0] w_sys_tmp1110;
	wire signed [31:0] w_sys_tmp1111;
	wire signed [31:0] w_sys_tmp1116;
	wire signed [31:0] w_sys_tmp1117;
	wire signed [31:0] w_sys_tmp1122;
	wire signed [31:0] w_sys_tmp1123;
	wire signed [31:0] w_sys_tmp1128;
	wire signed [31:0] w_sys_tmp1129;
	wire signed [31:0] w_sys_tmp1134;
	wire signed [31:0] w_sys_tmp1135;
	wire signed [31:0] w_sys_tmp1140;
	wire signed [31:0] w_sys_tmp1141;
	wire signed [31:0] w_sys_tmp1146;
	wire signed [31:0] w_sys_tmp1147;
	wire signed [31:0] w_sys_tmp1152;
	wire signed [31:0] w_sys_tmp1153;
	wire signed [31:0] w_sys_tmp1158;
	wire signed [31:0] w_sys_tmp1159;
	wire signed [31:0] w_sys_tmp1164;
	wire signed [31:0] w_sys_tmp1165;
	wire signed [31:0] w_sys_tmp1170;
	wire signed [31:0] w_sys_tmp1171;
	wire signed [31:0] w_sys_tmp1176;
	wire signed [31:0] w_sys_tmp1177;
	wire signed [31:0] w_sys_tmp1182;
	wire signed [31:0] w_sys_tmp1183;
	wire signed [31:0] w_sys_tmp1188;
	wire signed [31:0] w_sys_tmp1189;
	wire signed [31:0] w_sys_tmp1194;
	wire signed [31:0] w_sys_tmp1195;
	wire signed [31:0] w_sys_tmp1200;
	wire signed [31:0] w_sys_tmp1201;
	wire signed [31:0] w_sys_tmp1206;
	wire signed [31:0] w_sys_tmp1207;
	wire signed [31:0] w_sys_tmp1212;
	wire signed [31:0] w_sys_tmp1213;
	wire signed [31:0] w_sys_tmp1218;
	wire signed [31:0] w_sys_tmp1219;
	wire signed [31:0] w_sys_tmp1224;
	wire signed [31:0] w_sys_tmp1225;
	wire signed [31:0] w_sys_tmp1245;
	wire signed [31:0] w_sys_tmp1246;
	wire signed [31:0] w_sys_tmp1251;
	wire signed [31:0] w_sys_tmp1252;
	wire signed [31:0] w_sys_tmp1257;
	wire signed [31:0] w_sys_tmp1258;
	wire signed [31:0] w_sys_tmp1263;
	wire signed [31:0] w_sys_tmp1264;
	wire signed [31:0] w_sys_tmp1269;
	wire signed [31:0] w_sys_tmp1270;
	wire signed [31:0] w_sys_tmp1275;
	wire signed [31:0] w_sys_tmp1276;
	wire signed [31:0] w_sys_tmp1281;
	wire signed [31:0] w_sys_tmp1282;
	wire signed [31:0] w_sys_tmp1287;
	wire signed [31:0] w_sys_tmp1288;
	wire signed [31:0] w_sys_tmp1293;
	wire signed [31:0] w_sys_tmp1294;
	wire signed [31:0] w_sys_tmp1299;
	wire signed [31:0] w_sys_tmp1300;
	wire signed [31:0] w_sys_tmp1305;
	wire signed [31:0] w_sys_tmp1306;
	wire signed [31:0] w_sys_tmp1311;
	wire signed [31:0] w_sys_tmp1312;
	wire signed [31:0] w_sys_tmp1317;
	wire signed [31:0] w_sys_tmp1318;
	wire signed [31:0] w_sys_tmp1323;
	wire signed [31:0] w_sys_tmp1324;
	wire signed [31:0] w_sys_tmp1329;
	wire signed [31:0] w_sys_tmp1330;
	wire signed [31:0] w_sys_tmp1335;
	wire signed [31:0] w_sys_tmp1336;
	wire signed [31:0] w_sys_tmp1341;
	wire signed [31:0] w_sys_tmp1342;
	wire signed [31:0] w_sys_tmp1347;
	wire signed [31:0] w_sys_tmp1348;
	wire signed [31:0] w_sys_tmp1353;
	wire signed [31:0] w_sys_tmp1354;
	wire signed [31:0] w_sys_tmp1359;
	wire signed [31:0] w_sys_tmp1360;
	wire signed [31:0] w_sys_tmp1365;
	wire signed [31:0] w_sys_tmp1366;
	wire signed [31:0] w_sys_tmp1371;
	wire signed [31:0] w_sys_tmp1372;
	wire signed [31:0] w_sys_tmp1377;
	wire signed [31:0] w_sys_tmp1378;
	wire signed [31:0] w_sys_tmp1383;
	wire signed [31:0] w_sys_tmp1384;
	wire signed [31:0] w_sys_tmp1389;
	wire signed [31:0] w_sys_tmp1390;
	wire signed [31:0] w_sys_tmp1395;
	wire signed [31:0] w_sys_tmp1396;
	wire signed [31:0] w_sys_tmp1401;
	wire signed [31:0] w_sys_tmp1402;
	wire signed [31:0] w_sys_tmp1407;
	wire signed [31:0] w_sys_tmp1408;
	wire signed [31:0] w_sys_tmp1413;
	wire signed [31:0] w_sys_tmp1414;
	wire signed [31:0] w_sys_tmp1419;
	wire signed [31:0] w_sys_tmp1420;
	wire signed [31:0] w_sys_tmp1425;
	wire signed [31:0] w_sys_tmp1426;
	wire signed [31:0] w_sys_tmp1431;
	wire signed [31:0] w_sys_tmp1432;
	wire signed [31:0] w_sys_tmp1449;
	wire signed [31:0] w_sys_tmp1450;
	wire signed [31:0] w_sys_tmp1455;
	wire signed [31:0] w_sys_tmp1456;
	wire signed [31:0] w_sys_tmp1461;
	wire signed [31:0] w_sys_tmp1462;
	wire signed [31:0] w_sys_tmp1467;
	wire signed [31:0] w_sys_tmp1468;
	wire signed [31:0] w_sys_tmp1473;
	wire signed [31:0] w_sys_tmp1474;
	wire signed [31:0] w_sys_tmp1479;
	wire signed [31:0] w_sys_tmp1480;
	wire signed [31:0] w_sys_tmp1485;
	wire signed [31:0] w_sys_tmp1486;
	wire signed [31:0] w_sys_tmp1491;
	wire signed [31:0] w_sys_tmp1492;
	wire signed [31:0] w_sys_tmp1497;
	wire signed [31:0] w_sys_tmp1498;
	wire signed [31:0] w_sys_tmp1503;
	wire signed [31:0] w_sys_tmp1504;
	wire signed [31:0] w_sys_tmp1509;
	wire signed [31:0] w_sys_tmp1510;
	wire signed [31:0] w_sys_tmp1515;
	wire signed [31:0] w_sys_tmp1516;
	wire signed [31:0] w_sys_tmp1521;
	wire signed [31:0] w_sys_tmp1522;
	wire signed [31:0] w_sys_tmp1527;
	wire signed [31:0] w_sys_tmp1528;
	wire signed [31:0] w_sys_tmp1533;
	wire signed [31:0] w_sys_tmp1534;
	wire signed [31:0] w_sys_tmp1539;
	wire signed [31:0] w_sys_tmp1540;
	wire signed [31:0] w_sys_tmp1545;
	wire signed [31:0] w_sys_tmp1546;
	wire signed [31:0] w_sys_tmp1551;
	wire signed [31:0] w_sys_tmp1552;
	wire signed [31:0] w_sys_tmp1557;
	wire signed [31:0] w_sys_tmp1558;
	wire signed [31:0] w_sys_tmp1563;
	wire signed [31:0] w_sys_tmp1564;
	wire signed [31:0] w_sys_tmp1569;
	wire signed [31:0] w_sys_tmp1570;
	wire signed [31:0] w_sys_tmp1575;
	wire signed [31:0] w_sys_tmp1576;
	wire signed [31:0] w_sys_tmp1581;
	wire signed [31:0] w_sys_tmp1582;
	wire signed [31:0] w_sys_tmp1587;
	wire signed [31:0] w_sys_tmp1588;
	wire signed [31:0] w_sys_tmp1593;
	wire signed [31:0] w_sys_tmp1594;
	wire signed [31:0] w_sys_tmp1599;
	wire signed [31:0] w_sys_tmp1600;
	wire signed [31:0] w_sys_tmp1605;
	wire signed [31:0] w_sys_tmp1606;
	wire signed [31:0] w_sys_tmp1611;
	wire signed [31:0] w_sys_tmp1612;
	wire signed [31:0] w_sys_tmp1617;
	wire signed [31:0] w_sys_tmp1618;
	wire signed [31:0] w_sys_tmp1623;
	wire signed [31:0] w_sys_tmp1624;
	wire signed [31:0] w_sys_tmp1629;
	wire signed [31:0] w_sys_tmp1630;
	wire signed [31:0] w_sys_tmp1635;
	wire signed [31:0] w_sys_tmp1636;
	wire signed [31:0] w_sys_tmp1653;
	wire signed [31:0] w_sys_tmp1654;
	wire signed [31:0] w_sys_tmp1659;
	wire signed [31:0] w_sys_tmp1660;
	wire signed [31:0] w_sys_tmp1665;
	wire signed [31:0] w_sys_tmp1666;
	wire signed [31:0] w_sys_tmp1671;
	wire signed [31:0] w_sys_tmp1672;
	wire signed [31:0] w_sys_tmp1677;
	wire signed [31:0] w_sys_tmp1678;
	wire signed [31:0] w_sys_tmp1683;
	wire signed [31:0] w_sys_tmp1684;
	wire signed [31:0] w_sys_tmp1689;
	wire signed [31:0] w_sys_tmp1690;
	wire signed [31:0] w_sys_tmp1695;
	wire signed [31:0] w_sys_tmp1696;
	wire signed [31:0] w_sys_tmp1701;
	wire signed [31:0] w_sys_tmp1702;
	wire signed [31:0] w_sys_tmp1707;
	wire signed [31:0] w_sys_tmp1708;
	wire signed [31:0] w_sys_tmp1713;
	wire signed [31:0] w_sys_tmp1714;
	wire signed [31:0] w_sys_tmp1719;
	wire signed [31:0] w_sys_tmp1720;
	wire signed [31:0] w_sys_tmp1725;
	wire signed [31:0] w_sys_tmp1726;
	wire signed [31:0] w_sys_tmp1731;
	wire signed [31:0] w_sys_tmp1732;
	wire signed [31:0] w_sys_tmp1737;
	wire signed [31:0] w_sys_tmp1738;
	wire signed [31:0] w_sys_tmp1743;
	wire signed [31:0] w_sys_tmp1744;
	wire signed [31:0] w_sys_tmp1749;
	wire signed [31:0] w_sys_tmp1750;
	wire signed [31:0] w_sys_tmp1755;
	wire signed [31:0] w_sys_tmp1756;
	wire signed [31:0] w_sys_tmp1761;
	wire signed [31:0] w_sys_tmp1762;
	wire signed [31:0] w_sys_tmp1767;
	wire signed [31:0] w_sys_tmp1768;
	wire signed [31:0] w_sys_tmp1773;
	wire signed [31:0] w_sys_tmp1774;
	wire signed [31:0] w_sys_tmp1779;
	wire signed [31:0] w_sys_tmp1780;
	wire signed [31:0] w_sys_tmp1785;
	wire signed [31:0] w_sys_tmp1786;
	wire signed [31:0] w_sys_tmp1791;
	wire signed [31:0] w_sys_tmp1792;
	wire signed [31:0] w_sys_tmp1797;
	wire signed [31:0] w_sys_tmp1798;
	wire signed [31:0] w_sys_tmp1803;
	wire signed [31:0] w_sys_tmp1804;
	wire signed [31:0] w_sys_tmp1809;
	wire signed [31:0] w_sys_tmp1810;
	wire signed [31:0] w_sys_tmp1815;
	wire signed [31:0] w_sys_tmp1816;
	wire signed [31:0] w_sys_tmp1821;
	wire signed [31:0] w_sys_tmp1822;
	wire signed [31:0] w_sys_tmp1827;
	wire signed [31:0] w_sys_tmp1828;
	wire signed [31:0] w_sys_tmp1833;
	wire signed [31:0] w_sys_tmp1834;
	wire signed [31:0] w_sys_tmp1839;
	wire signed [31:0] w_sys_tmp1840;
	wire signed [31:0] w_sys_tmp1842;
	wire signed [31:0] w_sys_tmp1843;
	wire signed [31:0] w_sys_tmp1848;
	wire signed [31:0] w_sys_tmp1849;
	wire signed [31:0] w_sys_tmp1854;
	wire signed [31:0] w_sys_tmp1855;
	wire signed [31:0] w_sys_tmp1860;
	wire signed [31:0] w_sys_tmp1861;
	wire signed [31:0] w_sys_tmp1866;
	wire signed [31:0] w_sys_tmp1867;
	wire signed [31:0] w_sys_tmp1872;
	wire signed [31:0] w_sys_tmp1873;
	wire signed [31:0] w_sys_tmp1878;
	wire signed [31:0] w_sys_tmp1879;
	wire signed [31:0] w_sys_tmp1884;
	wire signed [31:0] w_sys_tmp1885;
	wire signed [31:0] w_sys_tmp1890;
	wire signed [31:0] w_sys_tmp1891;
	wire signed [31:0] w_sys_tmp1896;
	wire signed [31:0] w_sys_tmp1897;
	wire signed [31:0] w_sys_tmp1902;
	wire signed [31:0] w_sys_tmp1903;
	wire signed [31:0] w_sys_tmp1908;
	wire signed [31:0] w_sys_tmp1909;
	wire signed [31:0] w_sys_tmp1914;
	wire signed [31:0] w_sys_tmp1915;
	wire signed [31:0] w_sys_tmp1920;
	wire signed [31:0] w_sys_tmp1921;
	wire signed [31:0] w_sys_tmp1926;
	wire signed [31:0] w_sys_tmp1927;
	wire signed [31:0] w_sys_tmp1932;
	wire signed [31:0] w_sys_tmp1933;
	wire signed [31:0] w_sys_tmp1938;
	wire signed [31:0] w_sys_tmp1939;
	wire signed [31:0] w_sys_tmp1944;
	wire signed [31:0] w_sys_tmp1945;
	wire signed [31:0] w_sys_tmp1950;
	wire signed [31:0] w_sys_tmp1951;
	wire signed [31:0] w_sys_tmp1956;
	wire signed [31:0] w_sys_tmp1957;
	wire signed [31:0] w_sys_tmp1962;
	wire signed [31:0] w_sys_tmp1963;
	wire signed [31:0] w_sys_tmp1968;
	wire signed [31:0] w_sys_tmp1969;
	wire signed [31:0] w_sys_tmp1974;
	wire signed [31:0] w_sys_tmp1975;
	wire signed [31:0] w_sys_tmp1980;
	wire signed [31:0] w_sys_tmp1981;
	wire signed [31:0] w_sys_tmp1986;
	wire signed [31:0] w_sys_tmp1987;
	wire signed [31:0] w_sys_tmp1992;
	wire signed [31:0] w_sys_tmp1993;
	wire signed [31:0] w_sys_tmp1998;
	wire signed [31:0] w_sys_tmp1999;
	wire signed [31:0] w_sys_tmp2004;
	wire signed [31:0] w_sys_tmp2005;
	wire signed [31:0] w_sys_tmp2010;
	wire signed [31:0] w_sys_tmp2011;
	wire signed [31:0] w_sys_tmp2016;
	wire signed [31:0] w_sys_tmp2017;
	wire signed [31:0] w_sys_tmp2022;
	wire signed [31:0] w_sys_tmp2023;
	wire signed [31:0] w_sys_tmp2028;
	wire signed [31:0] w_sys_tmp2029;
	wire signed [31:0] w_sys_tmp2034;
	wire signed [31:0] w_sys_tmp2035;
	wire signed [31:0] w_sys_tmp2055;
	wire signed [31:0] w_sys_tmp2056;
	wire signed [31:0] w_sys_tmp2061;
	wire signed [31:0] w_sys_tmp2062;
	wire signed [31:0] w_sys_tmp2067;
	wire signed [31:0] w_sys_tmp2068;
	wire signed [31:0] w_sys_tmp2073;
	wire signed [31:0] w_sys_tmp2074;
	wire signed [31:0] w_sys_tmp2079;
	wire signed [31:0] w_sys_tmp2080;
	wire signed [31:0] w_sys_tmp2085;
	wire signed [31:0] w_sys_tmp2086;
	wire signed [31:0] w_sys_tmp2091;
	wire signed [31:0] w_sys_tmp2092;
	wire signed [31:0] w_sys_tmp2097;
	wire signed [31:0] w_sys_tmp2098;
	wire signed [31:0] w_sys_tmp2103;
	wire signed [31:0] w_sys_tmp2104;
	wire signed [31:0] w_sys_tmp2109;
	wire signed [31:0] w_sys_tmp2110;
	wire signed [31:0] w_sys_tmp2115;
	wire signed [31:0] w_sys_tmp2116;
	wire signed [31:0] w_sys_tmp2121;
	wire signed [31:0] w_sys_tmp2122;
	wire signed [31:0] w_sys_tmp2127;
	wire signed [31:0] w_sys_tmp2128;
	wire signed [31:0] w_sys_tmp2133;
	wire signed [31:0] w_sys_tmp2134;
	wire signed [31:0] w_sys_tmp2139;
	wire signed [31:0] w_sys_tmp2140;
	wire signed [31:0] w_sys_tmp2145;
	wire signed [31:0] w_sys_tmp2146;
	wire signed [31:0] w_sys_tmp2151;
	wire signed [31:0] w_sys_tmp2152;
	wire signed [31:0] w_sys_tmp2157;
	wire signed [31:0] w_sys_tmp2158;
	wire signed [31:0] w_sys_tmp2163;
	wire signed [31:0] w_sys_tmp2164;
	wire signed [31:0] w_sys_tmp2169;
	wire signed [31:0] w_sys_tmp2170;
	wire signed [31:0] w_sys_tmp2175;
	wire signed [31:0] w_sys_tmp2176;
	wire signed [31:0] w_sys_tmp2181;
	wire signed [31:0] w_sys_tmp2182;
	wire signed [31:0] w_sys_tmp2187;
	wire signed [31:0] w_sys_tmp2188;
	wire signed [31:0] w_sys_tmp2193;
	wire signed [31:0] w_sys_tmp2194;
	wire signed [31:0] w_sys_tmp2199;
	wire signed [31:0] w_sys_tmp2200;
	wire signed [31:0] w_sys_tmp2205;
	wire signed [31:0] w_sys_tmp2206;
	wire signed [31:0] w_sys_tmp2211;
	wire signed [31:0] w_sys_tmp2212;
	wire signed [31:0] w_sys_tmp2217;
	wire signed [31:0] w_sys_tmp2218;
	wire signed [31:0] w_sys_tmp2223;
	wire signed [31:0] w_sys_tmp2224;
	wire signed [31:0] w_sys_tmp2229;
	wire signed [31:0] w_sys_tmp2230;
	wire signed [31:0] w_sys_tmp2235;
	wire signed [31:0] w_sys_tmp2236;
	wire signed [31:0] w_sys_tmp2241;
	wire signed [31:0] w_sys_tmp2242;
	wire signed [31:0] w_sys_tmp2259;
	wire signed [31:0] w_sys_tmp2260;
	wire signed [31:0] w_sys_tmp2265;
	wire signed [31:0] w_sys_tmp2266;
	wire signed [31:0] w_sys_tmp2271;
	wire signed [31:0] w_sys_tmp2272;
	wire signed [31:0] w_sys_tmp2277;
	wire signed [31:0] w_sys_tmp2278;
	wire signed [31:0] w_sys_tmp2283;
	wire signed [31:0] w_sys_tmp2284;
	wire signed [31:0] w_sys_tmp2289;
	wire signed [31:0] w_sys_tmp2290;
	wire signed [31:0] w_sys_tmp2295;
	wire signed [31:0] w_sys_tmp2296;
	wire signed [31:0] w_sys_tmp2301;
	wire signed [31:0] w_sys_tmp2302;
	wire signed [31:0] w_sys_tmp2307;
	wire signed [31:0] w_sys_tmp2308;
	wire signed [31:0] w_sys_tmp2313;
	wire signed [31:0] w_sys_tmp2314;
	wire signed [31:0] w_sys_tmp2319;
	wire signed [31:0] w_sys_tmp2320;
	wire signed [31:0] w_sys_tmp2325;
	wire signed [31:0] w_sys_tmp2326;
	wire signed [31:0] w_sys_tmp2331;
	wire signed [31:0] w_sys_tmp2332;
	wire signed [31:0] w_sys_tmp2337;
	wire signed [31:0] w_sys_tmp2338;
	wire signed [31:0] w_sys_tmp2343;
	wire signed [31:0] w_sys_tmp2344;
	wire signed [31:0] w_sys_tmp2349;
	wire signed [31:0] w_sys_tmp2350;
	wire signed [31:0] w_sys_tmp2355;
	wire signed [31:0] w_sys_tmp2356;
	wire signed [31:0] w_sys_tmp2361;
	wire signed [31:0] w_sys_tmp2362;
	wire signed [31:0] w_sys_tmp2367;
	wire signed [31:0] w_sys_tmp2368;
	wire signed [31:0] w_sys_tmp2373;
	wire signed [31:0] w_sys_tmp2374;
	wire signed [31:0] w_sys_tmp2379;
	wire signed [31:0] w_sys_tmp2380;
	wire signed [31:0] w_sys_tmp2385;
	wire signed [31:0] w_sys_tmp2386;
	wire signed [31:0] w_sys_tmp2391;
	wire signed [31:0] w_sys_tmp2392;
	wire signed [31:0] w_sys_tmp2397;
	wire signed [31:0] w_sys_tmp2398;
	wire signed [31:0] w_sys_tmp2403;
	wire signed [31:0] w_sys_tmp2404;
	wire signed [31:0] w_sys_tmp2409;
	wire signed [31:0] w_sys_tmp2410;
	wire signed [31:0] w_sys_tmp2415;
	wire signed [31:0] w_sys_tmp2416;
	wire signed [31:0] w_sys_tmp2421;
	wire signed [31:0] w_sys_tmp2422;
	wire signed [31:0] w_sys_tmp2427;
	wire signed [31:0] w_sys_tmp2428;
	wire signed [31:0] w_sys_tmp2433;
	wire signed [31:0] w_sys_tmp2434;
	wire signed [31:0] w_sys_tmp2439;
	wire signed [31:0] w_sys_tmp2440;
	wire signed [31:0] w_sys_tmp2445;
	wire signed [31:0] w_sys_tmp2446;
	wire signed [31:0] w_sys_tmp2463;
	wire signed [31:0] w_sys_tmp2464;
	wire signed [31:0] w_sys_tmp2469;
	wire signed [31:0] w_sys_tmp2470;
	wire signed [31:0] w_sys_tmp2475;
	wire signed [31:0] w_sys_tmp2476;
	wire signed [31:0] w_sys_tmp2481;
	wire signed [31:0] w_sys_tmp2482;
	wire signed [31:0] w_sys_tmp2487;
	wire signed [31:0] w_sys_tmp2488;
	wire signed [31:0] w_sys_tmp2493;
	wire signed [31:0] w_sys_tmp2494;
	wire signed [31:0] w_sys_tmp2499;
	wire signed [31:0] w_sys_tmp2500;
	wire signed [31:0] w_sys_tmp2505;
	wire signed [31:0] w_sys_tmp2506;
	wire signed [31:0] w_sys_tmp2511;
	wire signed [31:0] w_sys_tmp2512;
	wire signed [31:0] w_sys_tmp2517;
	wire signed [31:0] w_sys_tmp2518;
	wire signed [31:0] w_sys_tmp2523;
	wire signed [31:0] w_sys_tmp2524;
	wire signed [31:0] w_sys_tmp2529;
	wire signed [31:0] w_sys_tmp2530;
	wire signed [31:0] w_sys_tmp2535;
	wire signed [31:0] w_sys_tmp2536;
	wire signed [31:0] w_sys_tmp2541;
	wire signed [31:0] w_sys_tmp2542;
	wire signed [31:0] w_sys_tmp2547;
	wire signed [31:0] w_sys_tmp2548;
	wire signed [31:0] w_sys_tmp2553;
	wire signed [31:0] w_sys_tmp2554;
	wire signed [31:0] w_sys_tmp2559;
	wire signed [31:0] w_sys_tmp2560;
	wire signed [31:0] w_sys_tmp2565;
	wire signed [31:0] w_sys_tmp2566;
	wire signed [31:0] w_sys_tmp2571;
	wire signed [31:0] w_sys_tmp2572;
	wire signed [31:0] w_sys_tmp2577;
	wire signed [31:0] w_sys_tmp2578;
	wire signed [31:0] w_sys_tmp2583;
	wire signed [31:0] w_sys_tmp2584;
	wire signed [31:0] w_sys_tmp2589;
	wire signed [31:0] w_sys_tmp2590;
	wire signed [31:0] w_sys_tmp2595;
	wire signed [31:0] w_sys_tmp2596;
	wire signed [31:0] w_sys_tmp2601;
	wire signed [31:0] w_sys_tmp2602;
	wire signed [31:0] w_sys_tmp2607;
	wire signed [31:0] w_sys_tmp2608;
	wire signed [31:0] w_sys_tmp2613;
	wire signed [31:0] w_sys_tmp2614;
	wire signed [31:0] w_sys_tmp2619;
	wire signed [31:0] w_sys_tmp2620;
	wire signed [31:0] w_sys_tmp2625;
	wire signed [31:0] w_sys_tmp2626;
	wire signed [31:0] w_sys_tmp2631;
	wire signed [31:0] w_sys_tmp2632;
	wire signed [31:0] w_sys_tmp2637;
	wire signed [31:0] w_sys_tmp2638;
	wire signed [31:0] w_sys_tmp2643;
	wire signed [31:0] w_sys_tmp2644;
	wire signed [31:0] w_sys_tmp2649;
	wire signed [31:0] w_sys_tmp2650;
	wire signed [31:0] w_sys_tmp2652;
	wire signed [31:0] w_sys_tmp2653;
	wire signed [31:0] w_sys_tmp2658;
	wire signed [31:0] w_sys_tmp2659;
	wire signed [31:0] w_sys_tmp2664;
	wire signed [31:0] w_sys_tmp2665;
	wire signed [31:0] w_sys_tmp2670;
	wire signed [31:0] w_sys_tmp2671;
	wire signed [31:0] w_sys_tmp2676;
	wire signed [31:0] w_sys_tmp2677;
	wire signed [31:0] w_sys_tmp2682;
	wire signed [31:0] w_sys_tmp2683;
	wire signed [31:0] w_sys_tmp2688;
	wire signed [31:0] w_sys_tmp2689;
	wire signed [31:0] w_sys_tmp2694;
	wire signed [31:0] w_sys_tmp2695;
	wire signed [31:0] w_sys_tmp2700;
	wire signed [31:0] w_sys_tmp2701;
	wire signed [31:0] w_sys_tmp2706;
	wire signed [31:0] w_sys_tmp2707;
	wire signed [31:0] w_sys_tmp2712;
	wire signed [31:0] w_sys_tmp2713;
	wire signed [31:0] w_sys_tmp2718;
	wire signed [31:0] w_sys_tmp2719;
	wire signed [31:0] w_sys_tmp2724;
	wire signed [31:0] w_sys_tmp2725;
	wire signed [31:0] w_sys_tmp2730;
	wire signed [31:0] w_sys_tmp2731;
	wire signed [31:0] w_sys_tmp2736;
	wire signed [31:0] w_sys_tmp2737;
	wire signed [31:0] w_sys_tmp2742;
	wire signed [31:0] w_sys_tmp2743;
	wire signed [31:0] w_sys_tmp2748;
	wire signed [31:0] w_sys_tmp2749;
	wire signed [31:0] w_sys_tmp2754;
	wire signed [31:0] w_sys_tmp2755;
	wire signed [31:0] w_sys_tmp2760;
	wire signed [31:0] w_sys_tmp2761;
	wire signed [31:0] w_sys_tmp2766;
	wire signed [31:0] w_sys_tmp2767;
	wire signed [31:0] w_sys_tmp2772;
	wire signed [31:0] w_sys_tmp2773;
	wire signed [31:0] w_sys_tmp2778;
	wire signed [31:0] w_sys_tmp2779;
	wire signed [31:0] w_sys_tmp2784;
	wire signed [31:0] w_sys_tmp2785;
	wire signed [31:0] w_sys_tmp2790;
	wire signed [31:0] w_sys_tmp2791;
	wire signed [31:0] w_sys_tmp2796;
	wire signed [31:0] w_sys_tmp2797;
	wire signed [31:0] w_sys_tmp2802;
	wire signed [31:0] w_sys_tmp2803;
	wire signed [31:0] w_sys_tmp2808;
	wire signed [31:0] w_sys_tmp2809;
	wire signed [31:0] w_sys_tmp2814;
	wire signed [31:0] w_sys_tmp2815;
	wire signed [31:0] w_sys_tmp2820;
	wire signed [31:0] w_sys_tmp2821;
	wire signed [31:0] w_sys_tmp2826;
	wire signed [31:0] w_sys_tmp2827;
	wire signed [31:0] w_sys_tmp2832;
	wire signed [31:0] w_sys_tmp2833;
	wire signed [31:0] w_sys_tmp2838;
	wire signed [31:0] w_sys_tmp2839;
	wire signed [31:0] w_sys_tmp2844;
	wire signed [31:0] w_sys_tmp2845;
	wire signed [31:0] w_sys_tmp2865;
	wire signed [31:0] w_sys_tmp2866;
	wire signed [31:0] w_sys_tmp2871;
	wire signed [31:0] w_sys_tmp2872;
	wire signed [31:0] w_sys_tmp2877;
	wire signed [31:0] w_sys_tmp2878;
	wire signed [31:0] w_sys_tmp2883;
	wire signed [31:0] w_sys_tmp2884;
	wire signed [31:0] w_sys_tmp2889;
	wire signed [31:0] w_sys_tmp2890;
	wire signed [31:0] w_sys_tmp2895;
	wire signed [31:0] w_sys_tmp2896;
	wire signed [31:0] w_sys_tmp2901;
	wire signed [31:0] w_sys_tmp2902;
	wire signed [31:0] w_sys_tmp2907;
	wire signed [31:0] w_sys_tmp2908;
	wire signed [31:0] w_sys_tmp2913;
	wire signed [31:0] w_sys_tmp2914;
	wire signed [31:0] w_sys_tmp2919;
	wire signed [31:0] w_sys_tmp2920;
	wire signed [31:0] w_sys_tmp2925;
	wire signed [31:0] w_sys_tmp2926;
	wire signed [31:0] w_sys_tmp2931;
	wire signed [31:0] w_sys_tmp2932;
	wire signed [31:0] w_sys_tmp2937;
	wire signed [31:0] w_sys_tmp2938;
	wire signed [31:0] w_sys_tmp2943;
	wire signed [31:0] w_sys_tmp2944;
	wire signed [31:0] w_sys_tmp2949;
	wire signed [31:0] w_sys_tmp2950;
	wire signed [31:0] w_sys_tmp2955;
	wire signed [31:0] w_sys_tmp2956;
	wire signed [31:0] w_sys_tmp2961;
	wire signed [31:0] w_sys_tmp2962;
	wire signed [31:0] w_sys_tmp2967;
	wire signed [31:0] w_sys_tmp2968;
	wire signed [31:0] w_sys_tmp2973;
	wire signed [31:0] w_sys_tmp2974;
	wire signed [31:0] w_sys_tmp2979;
	wire signed [31:0] w_sys_tmp2980;
	wire signed [31:0] w_sys_tmp2985;
	wire signed [31:0] w_sys_tmp2986;
	wire signed [31:0] w_sys_tmp2991;
	wire signed [31:0] w_sys_tmp2992;
	wire signed [31:0] w_sys_tmp2997;
	wire signed [31:0] w_sys_tmp2998;
	wire signed [31:0] w_sys_tmp3003;
	wire signed [31:0] w_sys_tmp3004;
	wire signed [31:0] w_sys_tmp3009;
	wire signed [31:0] w_sys_tmp3010;
	wire signed [31:0] w_sys_tmp3015;
	wire signed [31:0] w_sys_tmp3016;
	wire signed [31:0] w_sys_tmp3021;
	wire signed [31:0] w_sys_tmp3022;
	wire signed [31:0] w_sys_tmp3027;
	wire signed [31:0] w_sys_tmp3028;
	wire signed [31:0] w_sys_tmp3033;
	wire signed [31:0] w_sys_tmp3034;
	wire signed [31:0] w_sys_tmp3039;
	wire signed [31:0] w_sys_tmp3040;
	wire signed [31:0] w_sys_tmp3045;
	wire signed [31:0] w_sys_tmp3046;
	wire signed [31:0] w_sys_tmp3051;
	wire signed [31:0] w_sys_tmp3052;
	wire signed [31:0] w_sys_tmp3069;
	wire signed [31:0] w_sys_tmp3070;
	wire signed [31:0] w_sys_tmp3075;
	wire signed [31:0] w_sys_tmp3076;
	wire signed [31:0] w_sys_tmp3081;
	wire signed [31:0] w_sys_tmp3082;
	wire signed [31:0] w_sys_tmp3087;
	wire signed [31:0] w_sys_tmp3088;
	wire signed [31:0] w_sys_tmp3093;
	wire signed [31:0] w_sys_tmp3094;
	wire signed [31:0] w_sys_tmp3099;
	wire signed [31:0] w_sys_tmp3100;
	wire signed [31:0] w_sys_tmp3105;
	wire signed [31:0] w_sys_tmp3106;
	wire signed [31:0] w_sys_tmp3111;
	wire signed [31:0] w_sys_tmp3112;
	wire signed [31:0] w_sys_tmp3117;
	wire signed [31:0] w_sys_tmp3118;
	wire signed [31:0] w_sys_tmp3123;
	wire signed [31:0] w_sys_tmp3124;
	wire signed [31:0] w_sys_tmp3129;
	wire signed [31:0] w_sys_tmp3130;
	wire signed [31:0] w_sys_tmp3135;
	wire signed [31:0] w_sys_tmp3136;
	wire signed [31:0] w_sys_tmp3141;
	wire signed [31:0] w_sys_tmp3142;
	wire signed [31:0] w_sys_tmp3147;
	wire signed [31:0] w_sys_tmp3148;
	wire signed [31:0] w_sys_tmp3153;
	wire signed [31:0] w_sys_tmp3154;
	wire signed [31:0] w_sys_tmp3159;
	wire signed [31:0] w_sys_tmp3160;
	wire signed [31:0] w_sys_tmp3165;
	wire signed [31:0] w_sys_tmp3166;
	wire signed [31:0] w_sys_tmp3171;
	wire signed [31:0] w_sys_tmp3172;
	wire signed [31:0] w_sys_tmp3177;
	wire signed [31:0] w_sys_tmp3178;
	wire signed [31:0] w_sys_tmp3183;
	wire signed [31:0] w_sys_tmp3184;
	wire signed [31:0] w_sys_tmp3189;
	wire signed [31:0] w_sys_tmp3190;
	wire signed [31:0] w_sys_tmp3195;
	wire signed [31:0] w_sys_tmp3196;
	wire signed [31:0] w_sys_tmp3201;
	wire signed [31:0] w_sys_tmp3202;
	wire signed [31:0] w_sys_tmp3207;
	wire signed [31:0] w_sys_tmp3208;
	wire signed [31:0] w_sys_tmp3213;
	wire signed [31:0] w_sys_tmp3214;
	wire signed [31:0] w_sys_tmp3219;
	wire signed [31:0] w_sys_tmp3220;
	wire signed [31:0] w_sys_tmp3225;
	wire signed [31:0] w_sys_tmp3226;
	wire signed [31:0] w_sys_tmp3231;
	wire signed [31:0] w_sys_tmp3232;
	wire signed [31:0] w_sys_tmp3237;
	wire signed [31:0] w_sys_tmp3238;
	wire signed [31:0] w_sys_tmp3243;
	wire signed [31:0] w_sys_tmp3244;
	wire signed [31:0] w_sys_tmp3249;
	wire signed [31:0] w_sys_tmp3250;
	wire signed [31:0] w_sys_tmp3255;
	wire signed [31:0] w_sys_tmp3256;
	wire signed [31:0] w_sys_tmp3273;
	wire signed [31:0] w_sys_tmp3274;
	wire signed [31:0] w_sys_tmp3279;
	wire signed [31:0] w_sys_tmp3280;
	wire signed [31:0] w_sys_tmp3285;
	wire signed [31:0] w_sys_tmp3286;
	wire signed [31:0] w_sys_tmp3291;
	wire signed [31:0] w_sys_tmp3292;
	wire signed [31:0] w_sys_tmp3297;
	wire signed [31:0] w_sys_tmp3298;
	wire signed [31:0] w_sys_tmp3303;
	wire signed [31:0] w_sys_tmp3304;
	wire signed [31:0] w_sys_tmp3309;
	wire signed [31:0] w_sys_tmp3310;
	wire signed [31:0] w_sys_tmp3315;
	wire signed [31:0] w_sys_tmp3316;
	wire signed [31:0] w_sys_tmp3321;
	wire signed [31:0] w_sys_tmp3322;
	wire signed [31:0] w_sys_tmp3327;
	wire signed [31:0] w_sys_tmp3328;
	wire signed [31:0] w_sys_tmp3333;
	wire signed [31:0] w_sys_tmp3334;
	wire signed [31:0] w_sys_tmp3339;
	wire signed [31:0] w_sys_tmp3340;
	wire signed [31:0] w_sys_tmp3345;
	wire signed [31:0] w_sys_tmp3346;
	wire signed [31:0] w_sys_tmp3351;
	wire signed [31:0] w_sys_tmp3352;
	wire signed [31:0] w_sys_tmp3357;
	wire signed [31:0] w_sys_tmp3358;
	wire signed [31:0] w_sys_tmp3363;
	wire signed [31:0] w_sys_tmp3364;
	wire signed [31:0] w_sys_tmp3369;
	wire signed [31:0] w_sys_tmp3370;
	wire signed [31:0] w_sys_tmp3375;
	wire signed [31:0] w_sys_tmp3376;
	wire signed [31:0] w_sys_tmp3381;
	wire signed [31:0] w_sys_tmp3382;
	wire signed [31:0] w_sys_tmp3387;
	wire signed [31:0] w_sys_tmp3388;
	wire signed [31:0] w_sys_tmp3393;
	wire signed [31:0] w_sys_tmp3394;
	wire signed [31:0] w_sys_tmp3399;
	wire signed [31:0] w_sys_tmp3400;
	wire signed [31:0] w_sys_tmp3405;
	wire signed [31:0] w_sys_tmp3406;
	wire signed [31:0] w_sys_tmp3411;
	wire signed [31:0] w_sys_tmp3412;
	wire signed [31:0] w_sys_tmp3417;
	wire signed [31:0] w_sys_tmp3418;
	wire signed [31:0] w_sys_tmp3423;
	wire signed [31:0] w_sys_tmp3424;
	wire signed [31:0] w_sys_tmp3429;
	wire signed [31:0] w_sys_tmp3430;
	wire signed [31:0] w_sys_tmp3435;
	wire signed [31:0] w_sys_tmp3436;
	wire signed [31:0] w_sys_tmp3441;
	wire signed [31:0] w_sys_tmp3442;
	wire signed [31:0] w_sys_tmp3447;
	wire signed [31:0] w_sys_tmp3448;
	wire signed [31:0] w_sys_tmp3453;
	wire signed [31:0] w_sys_tmp3454;
	wire signed [31:0] w_sys_tmp3459;
	wire signed [31:0] w_sys_tmp3460;
	wire signed [31:0] w_sys_tmp3461;
	wire signed [31:0] w_sys_tmp3462;
	wire               w_sys_tmp3463;
	wire               w_sys_tmp3464;
	wire signed [31:0] w_sys_tmp3465;
	wire signed [31:0] w_sys_tmp3466;
	wire signed [31:0] w_sys_tmp3467;
	wire               w_sys_tmp3468;
	wire               w_sys_tmp3469;
	wire signed [31:0] w_sys_tmp3470;
	wire signed [31:0] w_sys_tmp3473;
	wire signed [31:0] w_sys_tmp3474;
	wire signed [31:0] w_sys_tmp3475;
	wire        [31:0] w_sys_tmp3476;
	wire signed [31:0] w_sys_tmp3477;
	wire signed [31:0] w_sys_tmp3478;
	wire signed [31:0] w_sys_tmp3480;
	wire signed [31:0] w_sys_tmp3481;
	wire signed [31:0] w_sys_tmp3542;
	wire               w_sys_tmp3543;
	wire               w_sys_tmp3544;
	wire signed [31:0] w_sys_tmp3545;
	wire signed [31:0] w_sys_tmp3548;
	wire signed [31:0] w_sys_tmp3549;
	wire signed [31:0] w_sys_tmp3550;
	wire        [31:0] w_sys_tmp3551;
	wire signed [31:0] w_sys_tmp3552;
	wire signed [31:0] w_sys_tmp3553;
	wire signed [31:0] w_sys_tmp3554;
	wire signed [31:0] w_sys_tmp3555;
	wire signed [31:0] w_sys_tmp3557;
	wire signed [31:0] w_sys_tmp3558;
	wire signed [31:0] w_sys_tmp3631;
	wire               w_sys_tmp3632;
	wire               w_sys_tmp3633;
	wire signed [31:0] w_sys_tmp3634;
	wire signed [31:0] w_sys_tmp3637;
	wire signed [31:0] w_sys_tmp3638;
	wire signed [31:0] w_sys_tmp3639;
	wire        [31:0] w_sys_tmp3640;
	wire signed [31:0] w_sys_tmp3641;
	wire signed [31:0] w_sys_tmp3642;
	wire signed [31:0] w_sys_tmp3643;
	wire signed [31:0] w_sys_tmp3644;
	wire signed [31:0] w_sys_tmp3646;
	wire signed [31:0] w_sys_tmp3647;
	wire signed [31:0] w_sys_tmp3720;
	wire               w_sys_tmp3721;
	wire               w_sys_tmp3722;
	wire signed [31:0] w_sys_tmp3723;
	wire signed [31:0] w_sys_tmp3726;
	wire signed [31:0] w_sys_tmp3727;
	wire signed [31:0] w_sys_tmp3728;
	wire        [31:0] w_sys_tmp3729;
	wire signed [31:0] w_sys_tmp3730;
	wire signed [31:0] w_sys_tmp3731;
	wire signed [31:0] w_sys_tmp3732;
	wire signed [31:0] w_sys_tmp3733;
	wire signed [31:0] w_sys_tmp3735;
	wire signed [31:0] w_sys_tmp3736;
	wire signed [31:0] w_sys_tmp3809;
	wire               w_sys_tmp3810;
	wire               w_sys_tmp3811;
	wire signed [31:0] w_sys_tmp3812;
	wire signed [31:0] w_sys_tmp3813;
	wire signed [31:0] w_sys_tmp3814;
	wire               w_sys_tmp3815;
	wire               w_sys_tmp3816;
	wire signed [31:0] w_sys_tmp3817;
	wire signed [31:0] w_sys_tmp3820;
	wire signed [31:0] w_sys_tmp3821;
	wire signed [31:0] w_sys_tmp3822;
	wire        [31:0] w_sys_tmp3823;
	wire signed [31:0] w_sys_tmp3824;
	wire signed [31:0] w_sys_tmp3825;
	wire signed [31:0] w_sys_tmp3827;
	wire signed [31:0] w_sys_tmp3828;
	wire signed [31:0] w_sys_tmp3889;
	wire               w_sys_tmp3890;
	wire               w_sys_tmp3891;
	wire signed [31:0] w_sys_tmp3892;
	wire signed [31:0] w_sys_tmp3895;
	wire signed [31:0] w_sys_tmp3896;
	wire signed [31:0] w_sys_tmp3897;
	wire        [31:0] w_sys_tmp3898;
	wire signed [31:0] w_sys_tmp3899;
	wire signed [31:0] w_sys_tmp3900;
	wire signed [31:0] w_sys_tmp3901;
	wire signed [31:0] w_sys_tmp3902;
	wire signed [31:0] w_sys_tmp3904;
	wire signed [31:0] w_sys_tmp3905;
	wire signed [31:0] w_sys_tmp3978;
	wire               w_sys_tmp3979;
	wire               w_sys_tmp3980;
	wire signed [31:0] w_sys_tmp3981;
	wire signed [31:0] w_sys_tmp3984;
	wire signed [31:0] w_sys_tmp3985;
	wire signed [31:0] w_sys_tmp3986;
	wire        [31:0] w_sys_tmp3987;
	wire signed [31:0] w_sys_tmp3988;
	wire signed [31:0] w_sys_tmp3989;
	wire signed [31:0] w_sys_tmp3990;
	wire signed [31:0] w_sys_tmp3991;
	wire signed [31:0] w_sys_tmp3993;
	wire signed [31:0] w_sys_tmp3994;
	wire signed [31:0] w_sys_tmp4067;
	wire               w_sys_tmp4068;
	wire               w_sys_tmp4069;
	wire signed [31:0] w_sys_tmp4070;
	wire signed [31:0] w_sys_tmp4073;
	wire signed [31:0] w_sys_tmp4074;
	wire signed [31:0] w_sys_tmp4075;
	wire        [31:0] w_sys_tmp4076;
	wire signed [31:0] w_sys_tmp4077;
	wire signed [31:0] w_sys_tmp4078;
	wire signed [31:0] w_sys_tmp4079;
	wire signed [31:0] w_sys_tmp4080;
	wire signed [31:0] w_sys_tmp4082;
	wire signed [31:0] w_sys_tmp4083;
	wire signed [31:0] w_sys_tmp4156;
	wire               w_sys_tmp4157;
	wire               w_sys_tmp4158;
	wire signed [31:0] w_sys_tmp4159;
	wire signed [31:0] w_sys_tmp4160;
	wire signed [31:0] w_sys_tmp4161;
	wire               w_sys_tmp4162;
	wire               w_sys_tmp4163;
	wire signed [31:0] w_sys_tmp4164;
	wire signed [31:0] w_sys_tmp4167;
	wire signed [31:0] w_sys_tmp4168;
	wire signed [31:0] w_sys_tmp4169;
	wire        [31:0] w_sys_tmp4170;
	wire signed [31:0] w_sys_tmp4171;
	wire signed [31:0] w_sys_tmp4172;
	wire signed [31:0] w_sys_tmp4174;
	wire signed [31:0] w_sys_tmp4175;
	wire signed [31:0] w_sys_tmp4236;
	wire               w_sys_tmp4237;
	wire               w_sys_tmp4238;
	wire signed [31:0] w_sys_tmp4239;
	wire signed [31:0] w_sys_tmp4242;
	wire signed [31:0] w_sys_tmp4243;
	wire signed [31:0] w_sys_tmp4244;
	wire        [31:0] w_sys_tmp4245;
	wire signed [31:0] w_sys_tmp4246;
	wire signed [31:0] w_sys_tmp4247;
	wire signed [31:0] w_sys_tmp4248;
	wire signed [31:0] w_sys_tmp4249;
	wire signed [31:0] w_sys_tmp4251;
	wire signed [31:0] w_sys_tmp4252;
	wire signed [31:0] w_sys_tmp4325;
	wire               w_sys_tmp4326;
	wire               w_sys_tmp4327;
	wire signed [31:0] w_sys_tmp4328;
	wire signed [31:0] w_sys_tmp4331;
	wire signed [31:0] w_sys_tmp4332;
	wire signed [31:0] w_sys_tmp4333;
	wire        [31:0] w_sys_tmp4334;
	wire signed [31:0] w_sys_tmp4335;
	wire signed [31:0] w_sys_tmp4336;
	wire signed [31:0] w_sys_tmp4337;
	wire signed [31:0] w_sys_tmp4338;
	wire signed [31:0] w_sys_tmp4340;
	wire signed [31:0] w_sys_tmp4341;
	wire signed [31:0] w_sys_tmp4414;
	wire               w_sys_tmp4415;
	wire               w_sys_tmp4416;
	wire signed [31:0] w_sys_tmp4417;
	wire signed [31:0] w_sys_tmp4420;
	wire signed [31:0] w_sys_tmp4421;
	wire signed [31:0] w_sys_tmp4422;
	wire        [31:0] w_sys_tmp4423;
	wire signed [31:0] w_sys_tmp4424;
	wire signed [31:0] w_sys_tmp4425;
	wire signed [31:0] w_sys_tmp4426;
	wire signed [31:0] w_sys_tmp4427;
	wire signed [31:0] w_sys_tmp4429;
	wire signed [31:0] w_sys_tmp4430;
	wire signed [31:0] w_sys_tmp4503;
	wire               w_sys_tmp4504;
	wire               w_sys_tmp4505;
	wire signed [31:0] w_sys_tmp4506;
	wire signed [31:0] w_sys_tmp4507;
	wire signed [31:0] w_sys_tmp4508;
	wire               w_sys_tmp4509;
	wire               w_sys_tmp4510;
	wire signed [31:0] w_sys_tmp4511;
	wire signed [31:0] w_sys_tmp4514;
	wire signed [31:0] w_sys_tmp4515;
	wire signed [31:0] w_sys_tmp4516;
	wire        [31:0] w_sys_tmp4517;
	wire signed [31:0] w_sys_tmp4518;
	wire signed [31:0] w_sys_tmp4519;
	wire signed [31:0] w_sys_tmp4521;
	wire signed [31:0] w_sys_tmp4522;
	wire signed [31:0] w_sys_tmp4583;
	wire               w_sys_tmp4584;
	wire               w_sys_tmp4585;
	wire signed [31:0] w_sys_tmp4586;
	wire signed [31:0] w_sys_tmp4589;
	wire signed [31:0] w_sys_tmp4590;
	wire signed [31:0] w_sys_tmp4591;
	wire        [31:0] w_sys_tmp4592;
	wire signed [31:0] w_sys_tmp4593;
	wire signed [31:0] w_sys_tmp4594;
	wire signed [31:0] w_sys_tmp4595;
	wire signed [31:0] w_sys_tmp4596;
	wire signed [31:0] w_sys_tmp4598;
	wire signed [31:0] w_sys_tmp4599;
	wire signed [31:0] w_sys_tmp4672;
	wire               w_sys_tmp4673;
	wire               w_sys_tmp4674;
	wire signed [31:0] w_sys_tmp4675;
	wire signed [31:0] w_sys_tmp4678;
	wire signed [31:0] w_sys_tmp4679;
	wire signed [31:0] w_sys_tmp4680;
	wire        [31:0] w_sys_tmp4681;
	wire signed [31:0] w_sys_tmp4682;
	wire signed [31:0] w_sys_tmp4683;
	wire signed [31:0] w_sys_tmp4684;
	wire signed [31:0] w_sys_tmp4685;
	wire signed [31:0] w_sys_tmp4687;
	wire signed [31:0] w_sys_tmp4688;
	wire signed [31:0] w_sys_tmp4761;
	wire               w_sys_tmp4762;
	wire               w_sys_tmp4763;
	wire signed [31:0] w_sys_tmp4764;
	wire signed [31:0] w_sys_tmp4767;
	wire signed [31:0] w_sys_tmp4768;
	wire signed [31:0] w_sys_tmp4769;
	wire        [31:0] w_sys_tmp4770;
	wire signed [31:0] w_sys_tmp4771;
	wire signed [31:0] w_sys_tmp4772;
	wire signed [31:0] w_sys_tmp4773;
	wire signed [31:0] w_sys_tmp4774;
	wire signed [31:0] w_sys_tmp4776;
	wire signed [31:0] w_sys_tmp4777;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 5'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 9'h1);
	assign w_fld_u_0_addr_0 = 15'sh0;
	assign w_fld_u_0_datain_0 = 32'h0;
	assign w_fld_u_0_r_w_0 = 1'h0;
	assign w_fld_u_0_ce_0 = w_sys_ce;
	assign w_fld_u_0_ce_1 = w_sys_ce;
	assign w_sub09_u_addr = ( (|r_sys_processing_methodID) ? r_sub09_u_addr : 13'sh0 ) ;
	assign w_sub09_u_datain = ( (|r_sys_processing_methodID) ? r_sub09_u_datain : 32'h0 ) ;
	assign w_sub09_u_r_w = ( (|r_sys_processing_methodID) ? r_sub09_u_r_w : 1'h0 ) ;
	assign w_sub09_result_addr = ( (|r_sys_processing_methodID) ? r_sub09_result_addr : 13'sh0 ) ;
	assign w_sub09_result_datain = ( (|r_sys_processing_methodID) ? r_sub09_result_datain : 32'h0 ) ;
	assign w_sub09_result_r_w = ( (|r_sys_processing_methodID) ? r_sub09_result_r_w : 1'h0 ) ;
	assign w_sub08_u_addr = ( (|r_sys_processing_methodID) ? r_sub08_u_addr : 13'sh0 ) ;
	assign w_sub08_u_datain = ( (|r_sys_processing_methodID) ? r_sub08_u_datain : 32'h0 ) ;
	assign w_sub08_u_r_w = ( (|r_sys_processing_methodID) ? r_sub08_u_r_w : 1'h0 ) ;
	assign w_sub08_result_addr = ( (|r_sys_processing_methodID) ? r_sub08_result_addr : 13'sh0 ) ;
	assign w_sub08_result_datain = ( (|r_sys_processing_methodID) ? r_sub08_result_datain : 32'h0 ) ;
	assign w_sub08_result_r_w = ( (|r_sys_processing_methodID) ? r_sub08_result_r_w : 1'h0 ) ;
	assign w_sub12_u_addr = ( (|r_sys_processing_methodID) ? r_sub12_u_addr : 13'sh0 ) ;
	assign w_sub12_u_datain = ( (|r_sys_processing_methodID) ? r_sub12_u_datain : 32'h0 ) ;
	assign w_sub12_u_r_w = ( (|r_sys_processing_methodID) ? r_sub12_u_r_w : 1'h0 ) ;
	assign w_sub12_result_addr = ( (|r_sys_processing_methodID) ? r_sub12_result_addr : 13'sh0 ) ;
	assign w_sub12_result_datain = ( (|r_sys_processing_methodID) ? r_sub12_result_datain : 32'h0 ) ;
	assign w_sub12_result_r_w = ( (|r_sys_processing_methodID) ? r_sub12_result_r_w : 1'h0 ) ;
	assign w_sub03_u_addr = ( (|r_sys_processing_methodID) ? r_sub03_u_addr : 13'sh0 ) ;
	assign w_sub03_u_datain = ( (|r_sys_processing_methodID) ? r_sub03_u_datain : 32'h0 ) ;
	assign w_sub03_u_r_w = ( (|r_sys_processing_methodID) ? r_sub03_u_r_w : 1'h0 ) ;
	assign w_sub03_result_addr = ( (|r_sys_processing_methodID) ? r_sub03_result_addr : 13'sh0 ) ;
	assign w_sub03_result_datain = ( (|r_sys_processing_methodID) ? r_sub03_result_datain : 32'h0 ) ;
	assign w_sub03_result_r_w = ( (|r_sys_processing_methodID) ? r_sub03_result_r_w : 1'h0 ) ;
	assign w_sub02_u_addr = ( (|r_sys_processing_methodID) ? r_sub02_u_addr : 13'sh0 ) ;
	assign w_sub02_u_datain = ( (|r_sys_processing_methodID) ? r_sub02_u_datain : 32'h0 ) ;
	assign w_sub02_u_r_w = ( (|r_sys_processing_methodID) ? r_sub02_u_r_w : 1'h0 ) ;
	assign w_sub02_result_addr = ( (|r_sys_processing_methodID) ? r_sub02_result_addr : 13'sh0 ) ;
	assign w_sub02_result_datain = ( (|r_sys_processing_methodID) ? r_sub02_result_datain : 32'h0 ) ;
	assign w_sub02_result_r_w = ( (|r_sys_processing_methodID) ? r_sub02_result_r_w : 1'h0 ) ;
	assign w_sub11_u_addr = ( (|r_sys_processing_methodID) ? r_sub11_u_addr : 13'sh0 ) ;
	assign w_sub11_u_datain = ( (|r_sys_processing_methodID) ? r_sub11_u_datain : 32'h0 ) ;
	assign w_sub11_u_r_w = ( (|r_sys_processing_methodID) ? r_sub11_u_r_w : 1'h0 ) ;
	assign w_sub11_result_addr = ( (|r_sys_processing_methodID) ? r_sub11_result_addr : 13'sh0 ) ;
	assign w_sub11_result_datain = ( (|r_sys_processing_methodID) ? r_sub11_result_datain : 32'h0 ) ;
	assign w_sub11_result_r_w = ( (|r_sys_processing_methodID) ? r_sub11_result_r_w : 1'h0 ) ;
	assign w_sub14_u_addr = ( (|r_sys_processing_methodID) ? r_sub14_u_addr : 13'sh0 ) ;
	assign w_sub14_u_datain = ( (|r_sys_processing_methodID) ? r_sub14_u_datain : 32'h0 ) ;
	assign w_sub14_u_r_w = ( (|r_sys_processing_methodID) ? r_sub14_u_r_w : 1'h0 ) ;
	assign w_sub14_result_addr = ( (|r_sys_processing_methodID) ? r_sub14_result_addr : 13'sh0 ) ;
	assign w_sub14_result_datain = ( (|r_sys_processing_methodID) ? r_sub14_result_datain : 32'h0 ) ;
	assign w_sub14_result_r_w = ( (|r_sys_processing_methodID) ? r_sub14_result_r_w : 1'h0 ) ;
	assign w_sub01_u_addr = ( (|r_sys_processing_methodID) ? r_sub01_u_addr : 13'sh0 ) ;
	assign w_sub01_u_datain = ( (|r_sys_processing_methodID) ? r_sub01_u_datain : 32'h0 ) ;
	assign w_sub01_u_r_w = ( (|r_sys_processing_methodID) ? r_sub01_u_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 13'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub13_u_addr = ( (|r_sys_processing_methodID) ? r_sub13_u_addr : 13'sh0 ) ;
	assign w_sub13_u_datain = ( (|r_sys_processing_methodID) ? r_sub13_u_datain : 32'h0 ) ;
	assign w_sub13_u_r_w = ( (|r_sys_processing_methodID) ? r_sub13_u_r_w : 1'h0 ) ;
	assign w_sub13_result_addr = ( (|r_sys_processing_methodID) ? r_sub13_result_addr : 13'sh0 ) ;
	assign w_sub13_result_datain = ( (|r_sys_processing_methodID) ? r_sub13_result_datain : 32'h0 ) ;
	assign w_sub13_result_r_w = ( (|r_sys_processing_methodID) ? r_sub13_result_r_w : 1'h0 ) ;
	assign w_sub00_u_addr = ( (|r_sys_processing_methodID) ? r_sub00_u_addr : 13'sh0 ) ;
	assign w_sub00_u_datain = ( (|r_sys_processing_methodID) ? r_sub00_u_datain : 32'h0 ) ;
	assign w_sub00_u_r_w = ( (|r_sys_processing_methodID) ? r_sub00_u_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 13'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sub07_u_addr = ( (|r_sys_processing_methodID) ? r_sub07_u_addr : 13'sh0 ) ;
	assign w_sub07_u_datain = ( (|r_sys_processing_methodID) ? r_sub07_u_datain : 32'h0 ) ;
	assign w_sub07_u_r_w = ( (|r_sys_processing_methodID) ? r_sub07_u_r_w : 1'h0 ) ;
	assign w_sub07_result_addr = ( (|r_sys_processing_methodID) ? r_sub07_result_addr : 13'sh0 ) ;
	assign w_sub07_result_datain = ( (|r_sys_processing_methodID) ? r_sub07_result_datain : 32'h0 ) ;
	assign w_sub07_result_r_w = ( (|r_sys_processing_methodID) ? r_sub07_result_r_w : 1'h0 ) ;
	assign w_sub06_u_addr = ( (|r_sys_processing_methodID) ? r_sub06_u_addr : 13'sh0 ) ;
	assign w_sub06_u_datain = ( (|r_sys_processing_methodID) ? r_sub06_u_datain : 32'h0 ) ;
	assign w_sub06_u_r_w = ( (|r_sys_processing_methodID) ? r_sub06_u_r_w : 1'h0 ) ;
	assign w_sub06_result_addr = ( (|r_sys_processing_methodID) ? r_sub06_result_addr : 13'sh0 ) ;
	assign w_sub06_result_datain = ( (|r_sys_processing_methodID) ? r_sub06_result_datain : 32'h0 ) ;
	assign w_sub06_result_r_w = ( (|r_sys_processing_methodID) ? r_sub06_result_r_w : 1'h0 ) ;
	assign w_sub15_u_addr = ( (|r_sys_processing_methodID) ? r_sub15_u_addr : 13'sh0 ) ;
	assign w_sub15_u_datain = ( (|r_sys_processing_methodID) ? r_sub15_u_datain : 32'h0 ) ;
	assign w_sub15_u_r_w = ( (|r_sys_processing_methodID) ? r_sub15_u_r_w : 1'h0 ) ;
	assign w_sub15_result_addr = ( (|r_sys_processing_methodID) ? r_sub15_result_addr : 13'sh0 ) ;
	assign w_sub15_result_datain = ( (|r_sys_processing_methodID) ? r_sub15_result_datain : 32'h0 ) ;
	assign w_sub15_result_r_w = ( (|r_sys_processing_methodID) ? r_sub15_result_r_w : 1'h0 ) ;
	assign w_sub05_u_addr = ( (|r_sys_processing_methodID) ? r_sub05_u_addr : 13'sh0 ) ;
	assign w_sub05_u_datain = ( (|r_sys_processing_methodID) ? r_sub05_u_datain : 32'h0 ) ;
	assign w_sub05_u_r_w = ( (|r_sys_processing_methodID) ? r_sub05_u_r_w : 1'h0 ) ;
	assign w_sub05_result_addr = ( (|r_sys_processing_methodID) ? r_sub05_result_addr : 13'sh0 ) ;
	assign w_sub05_result_datain = ( (|r_sys_processing_methodID) ? r_sub05_result_datain : 32'h0 ) ;
	assign w_sub05_result_r_w = ( (|r_sys_processing_methodID) ? r_sub05_result_r_w : 1'h0 ) ;
	assign w_sub04_u_addr = ( (|r_sys_processing_methodID) ? r_sub04_u_addr : 13'sh0 ) ;
	assign w_sub04_u_datain = ( (|r_sys_processing_methodID) ? r_sub04_u_datain : 32'h0 ) ;
	assign w_sub04_u_r_w = ( (|r_sys_processing_methodID) ? r_sub04_u_r_w : 1'h0 ) ;
	assign w_sub04_result_addr = ( (|r_sys_processing_methodID) ? r_sub04_result_addr : 13'sh0 ) ;
	assign w_sub04_result_datain = ( (|r_sys_processing_methodID) ? r_sub04_result_datain : 32'h0 ) ;
	assign w_sub04_result_r_w = ( (|r_sys_processing_methodID) ? r_sub04_result_r_w : 1'h0 ) ;
	assign w_sub10_u_addr = ( (|r_sys_processing_methodID) ? r_sub10_u_addr : 13'sh0 ) ;
	assign w_sub10_u_datain = ( (|r_sys_processing_methodID) ? r_sub10_u_datain : 32'h0 ) ;
	assign w_sub10_u_r_w = ( (|r_sys_processing_methodID) ? r_sub10_u_r_w : 1'h0 ) ;
	assign w_sub10_result_addr = ( (|r_sys_processing_methodID) ? r_sub10_result_addr : 13'sh0 ) ;
	assign w_sub10_result_datain = ( (|r_sys_processing_methodID) ? r_sub10_result_datain : 32'h0 ) ;
	assign w_sub10_result_r_w = ( (|r_sys_processing_methodID) ? r_sub10_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh00000081;
	assign w_sys_tmp3 = ( !w_sys_tmp4 );
	assign w_sys_tmp4 = (r_run_my_21 < r_run_k_17);
	assign w_sys_tmp5 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp6 = ( !w_sys_tmp7 );
	assign w_sys_tmp7 = (r_run_mx_20 < r_run_j_18);
	assign w_sys_tmp10 = (w_sys_tmp11 + r_run_k_17);
	assign w_sys_tmp11 = (r_run_j_18 * w_sys_tmp12);
	assign w_sys_tmp12 = 32'sh00000081;
	assign w_sys_tmp13 = 32'h0;
	assign w_sys_tmp14 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp51 = ( !w_sys_tmp52 );
	assign w_sys_tmp52 = (r_run_nlast_22 < r_run_n_19);
	assign w_sys_tmp53 = (r_run_n_19 + w_sys_intOne);
	assign w_sys_tmp54 = ( !w_sys_tmp55 );
	assign w_sys_tmp55 = (r_run_my_21 < r_run_j_18);
	assign w_sys_tmp58 = (w_sys_tmp59 + r_run_j_18);
	assign w_sys_tmp59 = 32'sh00000081;
	assign w_sys_tmp60 = 32'h3f000000;
	assign w_sys_tmp62 = (w_sys_tmp63 + r_run_copy2_j_25);
	assign w_sys_tmp63 = 32'sh00004101;
	assign w_sys_tmp64 = 32'h0;
	assign w_sys_tmp66 = (w_sys_tmp67 + w_sys_intOne);
	assign w_sys_tmp67 = (r_run_copy1_j_24 * w_sys_tmp59);
	assign w_sys_tmp69 = 32'h3f800000;
	assign w_sys_tmp71 = (w_sys_tmp72 + r_run_my_21);
	assign w_sys_tmp72 = (r_run_copy0_j_23 * w_sys_tmp59);
	assign w_sys_tmp75 = (r_run_copy0_j_23 + w_sys_intOne);
	assign w_sys_tmp76 = (r_run_copy1_j_24 + w_sys_intOne);
	assign w_sys_tmp77 = (r_run_copy2_j_25 + w_sys_intOne);
	assign w_sys_tmp78 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp211 = ( !w_sys_tmp212 );
	assign w_sys_tmp212 = (w_sys_tmp213 < r_run_k_17);
	assign w_sys_tmp213 = 32'sh00000021;
	assign w_sys_tmp216 = (w_sys_tmp217 + r_run_k_17);
	assign w_sys_tmp217 = 32'sh00000081;
	assign w_sys_tmp218 = w_fld_u_0_dataout_1;
	assign w_sys_tmp222 = (w_sys_tmp223 + r_run_k_17);
	assign w_sys_tmp223 = 32'sh00000102;
	assign w_sys_tmp228 = (w_sys_tmp229 + r_run_k_17);
	assign w_sys_tmp229 = 32'sh00000183;
	assign w_sys_tmp234 = (w_sys_tmp235 + r_run_k_17);
	assign w_sys_tmp235 = 32'sh00000204;
	assign w_sys_tmp240 = (w_sys_tmp241 + r_run_k_17);
	assign w_sys_tmp241 = 32'sh00000285;
	assign w_sys_tmp246 = (w_sys_tmp247 + r_run_k_17);
	assign w_sys_tmp247 = 32'sh00000306;
	assign w_sys_tmp252 = (w_sys_tmp253 + r_run_k_17);
	assign w_sys_tmp253 = 32'sh00000387;
	assign w_sys_tmp258 = (w_sys_tmp259 + r_run_k_17);
	assign w_sys_tmp259 = 32'sh00000408;
	assign w_sys_tmp264 = (w_sys_tmp265 + r_run_k_17);
	assign w_sys_tmp265 = 32'sh00000489;
	assign w_sys_tmp270 = (w_sys_tmp271 + r_run_k_17);
	assign w_sys_tmp271 = 32'sh0000050a;
	assign w_sys_tmp276 = (w_sys_tmp277 + r_run_k_17);
	assign w_sys_tmp277 = 32'sh0000058b;
	assign w_sys_tmp282 = (w_sys_tmp283 + r_run_k_17);
	assign w_sys_tmp283 = 32'sh0000060c;
	assign w_sys_tmp288 = (w_sys_tmp289 + r_run_k_17);
	assign w_sys_tmp289 = 32'sh0000068d;
	assign w_sys_tmp294 = (w_sys_tmp295 + r_run_k_17);
	assign w_sys_tmp295 = 32'sh0000070e;
	assign w_sys_tmp300 = (w_sys_tmp301 + r_run_k_17);
	assign w_sys_tmp301 = 32'sh0000078f;
	assign w_sys_tmp306 = (w_sys_tmp307 + r_run_k_17);
	assign w_sys_tmp307 = 32'sh00000810;
	assign w_sys_tmp312 = (w_sys_tmp313 + r_run_k_17);
	assign w_sys_tmp313 = 32'sh00000891;
	assign w_sys_tmp318 = (w_sys_tmp319 + r_run_k_17);
	assign w_sys_tmp319 = 32'sh00000912;
	assign w_sys_tmp324 = (w_sys_tmp325 + r_run_k_17);
	assign w_sys_tmp325 = 32'sh00000993;
	assign w_sys_tmp330 = (w_sys_tmp331 + r_run_k_17);
	assign w_sys_tmp331 = 32'sh00000a14;
	assign w_sys_tmp336 = (w_sys_tmp337 + r_run_k_17);
	assign w_sys_tmp337 = 32'sh00000a95;
	assign w_sys_tmp342 = (w_sys_tmp343 + r_run_k_17);
	assign w_sys_tmp343 = 32'sh00000b16;
	assign w_sys_tmp348 = (w_sys_tmp349 + r_run_k_17);
	assign w_sys_tmp349 = 32'sh00000b97;
	assign w_sys_tmp354 = (w_sys_tmp355 + r_run_k_17);
	assign w_sys_tmp355 = 32'sh00000c18;
	assign w_sys_tmp360 = (w_sys_tmp361 + r_run_k_17);
	assign w_sys_tmp361 = 32'sh00000c99;
	assign w_sys_tmp366 = (w_sys_tmp367 + r_run_k_17);
	assign w_sys_tmp367 = 32'sh00000d1a;
	assign w_sys_tmp372 = (w_sys_tmp373 + r_run_k_17);
	assign w_sys_tmp373 = 32'sh00000d9b;
	assign w_sys_tmp378 = (w_sys_tmp379 + r_run_k_17);
	assign w_sys_tmp379 = 32'sh00000e1c;
	assign w_sys_tmp384 = (w_sys_tmp385 + r_run_k_17);
	assign w_sys_tmp385 = 32'sh00000e9d;
	assign w_sys_tmp390 = (w_sys_tmp391 + r_run_k_17);
	assign w_sys_tmp391 = 32'sh00000f1e;
	assign w_sys_tmp396 = (w_sys_tmp397 + r_run_k_17);
	assign w_sys_tmp397 = 32'sh00000f9f;
	assign w_sys_tmp402 = (w_sys_tmp403 + r_run_k_17);
	assign w_sys_tmp403 = 32'sh00001020;
	assign w_sys_tmp408 = (w_sys_tmp409 + r_run_k_17);
	assign w_sys_tmp409 = 32'sh000010a1;
	assign w_sys_tmp429 = (w_sys_tmp430 + r_run_k_17);
	assign w_sys_tmp430 = 32'sh00001122;
	assign w_sys_tmp435 = (w_sys_tmp436 + r_run_k_17);
	assign w_sys_tmp436 = 32'sh000011a3;
	assign w_sys_tmp441 = (w_sys_tmp442 + r_run_k_17);
	assign w_sys_tmp442 = 32'sh00001224;
	assign w_sys_tmp447 = (w_sys_tmp448 + r_run_k_17);
	assign w_sys_tmp448 = 32'sh000012a5;
	assign w_sys_tmp453 = (w_sys_tmp454 + r_run_k_17);
	assign w_sys_tmp454 = 32'sh00001326;
	assign w_sys_tmp459 = (w_sys_tmp460 + r_run_k_17);
	assign w_sys_tmp460 = 32'sh000013a7;
	assign w_sys_tmp465 = (w_sys_tmp466 + r_run_k_17);
	assign w_sys_tmp466 = 32'sh00001428;
	assign w_sys_tmp471 = (w_sys_tmp472 + r_run_k_17);
	assign w_sys_tmp472 = 32'sh000014a9;
	assign w_sys_tmp477 = (w_sys_tmp478 + r_run_k_17);
	assign w_sys_tmp478 = 32'sh0000152a;
	assign w_sys_tmp483 = (w_sys_tmp484 + r_run_k_17);
	assign w_sys_tmp484 = 32'sh000015ab;
	assign w_sys_tmp489 = (w_sys_tmp490 + r_run_k_17);
	assign w_sys_tmp490 = 32'sh0000162c;
	assign w_sys_tmp495 = (w_sys_tmp496 + r_run_k_17);
	assign w_sys_tmp496 = 32'sh000016ad;
	assign w_sys_tmp501 = (w_sys_tmp502 + r_run_k_17);
	assign w_sys_tmp502 = 32'sh0000172e;
	assign w_sys_tmp507 = (w_sys_tmp508 + r_run_k_17);
	assign w_sys_tmp508 = 32'sh000017af;
	assign w_sys_tmp513 = (w_sys_tmp514 + r_run_k_17);
	assign w_sys_tmp514 = 32'sh00001830;
	assign w_sys_tmp519 = (w_sys_tmp520 + r_run_k_17);
	assign w_sys_tmp520 = 32'sh000018b1;
	assign w_sys_tmp525 = (w_sys_tmp526 + r_run_k_17);
	assign w_sys_tmp526 = 32'sh00001932;
	assign w_sys_tmp531 = (w_sys_tmp532 + r_run_k_17);
	assign w_sys_tmp532 = 32'sh000019b3;
	assign w_sys_tmp537 = (w_sys_tmp538 + r_run_k_17);
	assign w_sys_tmp538 = 32'sh00001a34;
	assign w_sys_tmp543 = (w_sys_tmp544 + r_run_k_17);
	assign w_sys_tmp544 = 32'sh00001ab5;
	assign w_sys_tmp549 = (w_sys_tmp550 + r_run_k_17);
	assign w_sys_tmp550 = 32'sh00001b36;
	assign w_sys_tmp555 = (w_sys_tmp556 + r_run_k_17);
	assign w_sys_tmp556 = 32'sh00001bb7;
	assign w_sys_tmp561 = (w_sys_tmp562 + r_run_k_17);
	assign w_sys_tmp562 = 32'sh00001c38;
	assign w_sys_tmp567 = (w_sys_tmp568 + r_run_k_17);
	assign w_sys_tmp568 = 32'sh00001cb9;
	assign w_sys_tmp573 = (w_sys_tmp574 + r_run_k_17);
	assign w_sys_tmp574 = 32'sh00001d3a;
	assign w_sys_tmp579 = (w_sys_tmp580 + r_run_k_17);
	assign w_sys_tmp580 = 32'sh00001dbb;
	assign w_sys_tmp585 = (w_sys_tmp586 + r_run_k_17);
	assign w_sys_tmp586 = 32'sh00001e3c;
	assign w_sys_tmp591 = (w_sys_tmp592 + r_run_k_17);
	assign w_sys_tmp592 = 32'sh00001ebd;
	assign w_sys_tmp597 = (w_sys_tmp598 + r_run_k_17);
	assign w_sys_tmp598 = 32'sh00001f3e;
	assign w_sys_tmp603 = (w_sys_tmp604 + r_run_k_17);
	assign w_sys_tmp604 = 32'sh00001fbf;
	assign w_sys_tmp609 = (w_sys_tmp610 + r_run_k_17);
	assign w_sys_tmp610 = 32'sh00002040;
	assign w_sys_tmp615 = (w_sys_tmp616 + r_run_k_17);
	assign w_sys_tmp616 = 32'sh000020c1;
	assign w_sys_tmp633 = (w_sys_tmp634 + r_run_k_17);
	assign w_sys_tmp634 = 32'sh00002142;
	assign w_sys_tmp639 = (w_sys_tmp640 + r_run_k_17);
	assign w_sys_tmp640 = 32'sh000021c3;
	assign w_sys_tmp645 = (w_sys_tmp646 + r_run_k_17);
	assign w_sys_tmp646 = 32'sh00002244;
	assign w_sys_tmp651 = (w_sys_tmp652 + r_run_k_17);
	assign w_sys_tmp652 = 32'sh000022c5;
	assign w_sys_tmp657 = (w_sys_tmp658 + r_run_k_17);
	assign w_sys_tmp658 = 32'sh00002346;
	assign w_sys_tmp663 = (w_sys_tmp664 + r_run_k_17);
	assign w_sys_tmp664 = 32'sh000023c7;
	assign w_sys_tmp669 = (w_sys_tmp670 + r_run_k_17);
	assign w_sys_tmp670 = 32'sh00002448;
	assign w_sys_tmp675 = (w_sys_tmp676 + r_run_k_17);
	assign w_sys_tmp676 = 32'sh000024c9;
	assign w_sys_tmp681 = (w_sys_tmp682 + r_run_k_17);
	assign w_sys_tmp682 = 32'sh0000254a;
	assign w_sys_tmp687 = (w_sys_tmp688 + r_run_k_17);
	assign w_sys_tmp688 = 32'sh000025cb;
	assign w_sys_tmp693 = (w_sys_tmp694 + r_run_k_17);
	assign w_sys_tmp694 = 32'sh0000264c;
	assign w_sys_tmp699 = (w_sys_tmp700 + r_run_k_17);
	assign w_sys_tmp700 = 32'sh000026cd;
	assign w_sys_tmp705 = (w_sys_tmp706 + r_run_k_17);
	assign w_sys_tmp706 = 32'sh0000274e;
	assign w_sys_tmp711 = (w_sys_tmp712 + r_run_k_17);
	assign w_sys_tmp712 = 32'sh000027cf;
	assign w_sys_tmp717 = (w_sys_tmp718 + r_run_k_17);
	assign w_sys_tmp718 = 32'sh00002850;
	assign w_sys_tmp723 = (w_sys_tmp724 + r_run_k_17);
	assign w_sys_tmp724 = 32'sh000028d1;
	assign w_sys_tmp729 = (w_sys_tmp730 + r_run_k_17);
	assign w_sys_tmp730 = 32'sh00002952;
	assign w_sys_tmp735 = (w_sys_tmp736 + r_run_k_17);
	assign w_sys_tmp736 = 32'sh000029d3;
	assign w_sys_tmp741 = (w_sys_tmp742 + r_run_k_17);
	assign w_sys_tmp742 = 32'sh00002a54;
	assign w_sys_tmp747 = (w_sys_tmp748 + r_run_k_17);
	assign w_sys_tmp748 = 32'sh00002ad5;
	assign w_sys_tmp753 = (w_sys_tmp754 + r_run_k_17);
	assign w_sys_tmp754 = 32'sh00002b56;
	assign w_sys_tmp759 = (w_sys_tmp760 + r_run_k_17);
	assign w_sys_tmp760 = 32'sh00002bd7;
	assign w_sys_tmp765 = (w_sys_tmp766 + r_run_k_17);
	assign w_sys_tmp766 = 32'sh00002c58;
	assign w_sys_tmp771 = (w_sys_tmp772 + r_run_k_17);
	assign w_sys_tmp772 = 32'sh00002cd9;
	assign w_sys_tmp777 = (w_sys_tmp778 + r_run_k_17);
	assign w_sys_tmp778 = 32'sh00002d5a;
	assign w_sys_tmp783 = (w_sys_tmp784 + r_run_k_17);
	assign w_sys_tmp784 = 32'sh00002ddb;
	assign w_sys_tmp789 = (w_sys_tmp790 + r_run_k_17);
	assign w_sys_tmp790 = 32'sh00002e5c;
	assign w_sys_tmp795 = (w_sys_tmp796 + r_run_k_17);
	assign w_sys_tmp796 = 32'sh00002edd;
	assign w_sys_tmp801 = (w_sys_tmp802 + r_run_k_17);
	assign w_sys_tmp802 = 32'sh00002f5e;
	assign w_sys_tmp807 = (w_sys_tmp808 + r_run_k_17);
	assign w_sys_tmp808 = 32'sh00002fdf;
	assign w_sys_tmp813 = (w_sys_tmp814 + r_run_k_17);
	assign w_sys_tmp814 = 32'sh00003060;
	assign w_sys_tmp819 = (w_sys_tmp820 + r_run_k_17);
	assign w_sys_tmp820 = 32'sh000030e1;
	assign w_sys_tmp837 = (w_sys_tmp838 + r_run_k_17);
	assign w_sys_tmp838 = 32'sh00003162;
	assign w_sys_tmp843 = (w_sys_tmp844 + r_run_k_17);
	assign w_sys_tmp844 = 32'sh000031e3;
	assign w_sys_tmp849 = (w_sys_tmp850 + r_run_k_17);
	assign w_sys_tmp850 = 32'sh00003264;
	assign w_sys_tmp855 = (w_sys_tmp856 + r_run_k_17);
	assign w_sys_tmp856 = 32'sh000032e5;
	assign w_sys_tmp861 = (w_sys_tmp862 + r_run_k_17);
	assign w_sys_tmp862 = 32'sh00003366;
	assign w_sys_tmp867 = (w_sys_tmp868 + r_run_k_17);
	assign w_sys_tmp868 = 32'sh000033e7;
	assign w_sys_tmp873 = (w_sys_tmp874 + r_run_k_17);
	assign w_sys_tmp874 = 32'sh00003468;
	assign w_sys_tmp879 = (w_sys_tmp880 + r_run_k_17);
	assign w_sys_tmp880 = 32'sh000034e9;
	assign w_sys_tmp885 = (w_sys_tmp886 + r_run_k_17);
	assign w_sys_tmp886 = 32'sh0000356a;
	assign w_sys_tmp891 = (w_sys_tmp892 + r_run_k_17);
	assign w_sys_tmp892 = 32'sh000035eb;
	assign w_sys_tmp897 = (w_sys_tmp898 + r_run_k_17);
	assign w_sys_tmp898 = 32'sh0000366c;
	assign w_sys_tmp903 = (w_sys_tmp904 + r_run_k_17);
	assign w_sys_tmp904 = 32'sh000036ed;
	assign w_sys_tmp909 = (w_sys_tmp910 + r_run_k_17);
	assign w_sys_tmp910 = 32'sh0000376e;
	assign w_sys_tmp915 = (w_sys_tmp916 + r_run_k_17);
	assign w_sys_tmp916 = 32'sh000037ef;
	assign w_sys_tmp921 = (w_sys_tmp922 + r_run_k_17);
	assign w_sys_tmp922 = 32'sh00003870;
	assign w_sys_tmp927 = (w_sys_tmp928 + r_run_k_17);
	assign w_sys_tmp928 = 32'sh000038f1;
	assign w_sys_tmp933 = (w_sys_tmp934 + r_run_k_17);
	assign w_sys_tmp934 = 32'sh00003972;
	assign w_sys_tmp939 = (w_sys_tmp940 + r_run_k_17);
	assign w_sys_tmp940 = 32'sh000039f3;
	assign w_sys_tmp945 = (w_sys_tmp946 + r_run_k_17);
	assign w_sys_tmp946 = 32'sh00003a74;
	assign w_sys_tmp951 = (w_sys_tmp952 + r_run_k_17);
	assign w_sys_tmp952 = 32'sh00003af5;
	assign w_sys_tmp957 = (w_sys_tmp958 + r_run_k_17);
	assign w_sys_tmp958 = 32'sh00003b76;
	assign w_sys_tmp963 = (w_sys_tmp964 + r_run_k_17);
	assign w_sys_tmp964 = 32'sh00003bf7;
	assign w_sys_tmp969 = (w_sys_tmp970 + r_run_k_17);
	assign w_sys_tmp970 = 32'sh00003c78;
	assign w_sys_tmp975 = (w_sys_tmp976 + r_run_k_17);
	assign w_sys_tmp976 = 32'sh00003cf9;
	assign w_sys_tmp981 = (w_sys_tmp982 + r_run_k_17);
	assign w_sys_tmp982 = 32'sh00003d7a;
	assign w_sys_tmp987 = (w_sys_tmp988 + r_run_k_17);
	assign w_sys_tmp988 = 32'sh00003dfb;
	assign w_sys_tmp993 = (w_sys_tmp994 + r_run_k_17);
	assign w_sys_tmp994 = 32'sh00003e7c;
	assign w_sys_tmp999 = (w_sys_tmp1000 + r_run_k_17);
	assign w_sys_tmp1000 = 32'sh00003efd;
	assign w_sys_tmp1005 = (w_sys_tmp1006 + r_run_k_17);
	assign w_sys_tmp1006 = 32'sh00003f7e;
	assign w_sys_tmp1011 = (w_sys_tmp1012 + r_run_k_17);
	assign w_sys_tmp1012 = 32'sh00003fff;
	assign w_sys_tmp1017 = (w_sys_tmp1018 + r_run_k_17);
	assign w_sys_tmp1018 = 32'sh00004080;
	assign w_sys_tmp1023 = (w_sys_tmp1024 + r_run_k_17);
	assign w_sys_tmp1024 = 32'sh00004101;
	assign w_sys_tmp1025 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp1026 = 32'sh00000020;
	assign w_sys_tmp1027 = ( !w_sys_tmp1028 );
	assign w_sys_tmp1028 = (w_sys_tmp1029 < r_run_k_17);
	assign w_sys_tmp1029 = 32'sh00000041;
	assign w_sys_tmp1032 = (w_sys_tmp1033 + r_run_k_17);
	assign w_sys_tmp1033 = 32'sh00000081;
	assign w_sys_tmp1034 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1038 = (w_sys_tmp1039 + r_run_k_17);
	assign w_sys_tmp1039 = 32'sh00000102;
	assign w_sys_tmp1044 = (w_sys_tmp1045 + r_run_k_17);
	assign w_sys_tmp1045 = 32'sh00000183;
	assign w_sys_tmp1050 = (w_sys_tmp1051 + r_run_k_17);
	assign w_sys_tmp1051 = 32'sh00000204;
	assign w_sys_tmp1056 = (w_sys_tmp1057 + r_run_k_17);
	assign w_sys_tmp1057 = 32'sh00000285;
	assign w_sys_tmp1062 = (w_sys_tmp1063 + r_run_k_17);
	assign w_sys_tmp1063 = 32'sh00000306;
	assign w_sys_tmp1068 = (w_sys_tmp1069 + r_run_k_17);
	assign w_sys_tmp1069 = 32'sh00000387;
	assign w_sys_tmp1074 = (w_sys_tmp1075 + r_run_k_17);
	assign w_sys_tmp1075 = 32'sh00000408;
	assign w_sys_tmp1080 = (w_sys_tmp1081 + r_run_k_17);
	assign w_sys_tmp1081 = 32'sh00000489;
	assign w_sys_tmp1086 = (w_sys_tmp1087 + r_run_k_17);
	assign w_sys_tmp1087 = 32'sh0000050a;
	assign w_sys_tmp1092 = (w_sys_tmp1093 + r_run_k_17);
	assign w_sys_tmp1093 = 32'sh0000058b;
	assign w_sys_tmp1098 = (w_sys_tmp1099 + r_run_k_17);
	assign w_sys_tmp1099 = 32'sh0000060c;
	assign w_sys_tmp1104 = (w_sys_tmp1105 + r_run_k_17);
	assign w_sys_tmp1105 = 32'sh0000068d;
	assign w_sys_tmp1110 = (w_sys_tmp1111 + r_run_k_17);
	assign w_sys_tmp1111 = 32'sh0000070e;
	assign w_sys_tmp1116 = (w_sys_tmp1117 + r_run_k_17);
	assign w_sys_tmp1117 = 32'sh0000078f;
	assign w_sys_tmp1122 = (w_sys_tmp1123 + r_run_k_17);
	assign w_sys_tmp1123 = 32'sh00000810;
	assign w_sys_tmp1128 = (w_sys_tmp1129 + r_run_k_17);
	assign w_sys_tmp1129 = 32'sh00000891;
	assign w_sys_tmp1134 = (w_sys_tmp1135 + r_run_k_17);
	assign w_sys_tmp1135 = 32'sh00000912;
	assign w_sys_tmp1140 = (w_sys_tmp1141 + r_run_k_17);
	assign w_sys_tmp1141 = 32'sh00000993;
	assign w_sys_tmp1146 = (w_sys_tmp1147 + r_run_k_17);
	assign w_sys_tmp1147 = 32'sh00000a14;
	assign w_sys_tmp1152 = (w_sys_tmp1153 + r_run_k_17);
	assign w_sys_tmp1153 = 32'sh00000a95;
	assign w_sys_tmp1158 = (w_sys_tmp1159 + r_run_k_17);
	assign w_sys_tmp1159 = 32'sh00000b16;
	assign w_sys_tmp1164 = (w_sys_tmp1165 + r_run_k_17);
	assign w_sys_tmp1165 = 32'sh00000b97;
	assign w_sys_tmp1170 = (w_sys_tmp1171 + r_run_k_17);
	assign w_sys_tmp1171 = 32'sh00000c18;
	assign w_sys_tmp1176 = (w_sys_tmp1177 + r_run_k_17);
	assign w_sys_tmp1177 = 32'sh00000c99;
	assign w_sys_tmp1182 = (w_sys_tmp1183 + r_run_k_17);
	assign w_sys_tmp1183 = 32'sh00000d1a;
	assign w_sys_tmp1188 = (w_sys_tmp1189 + r_run_k_17);
	assign w_sys_tmp1189 = 32'sh00000d9b;
	assign w_sys_tmp1194 = (w_sys_tmp1195 + r_run_k_17);
	assign w_sys_tmp1195 = 32'sh00000e1c;
	assign w_sys_tmp1200 = (w_sys_tmp1201 + r_run_k_17);
	assign w_sys_tmp1201 = 32'sh00000e9d;
	assign w_sys_tmp1206 = (w_sys_tmp1207 + r_run_k_17);
	assign w_sys_tmp1207 = 32'sh00000f1e;
	assign w_sys_tmp1212 = (w_sys_tmp1213 + r_run_k_17);
	assign w_sys_tmp1213 = 32'sh00000f9f;
	assign w_sys_tmp1218 = (w_sys_tmp1219 + r_run_k_17);
	assign w_sys_tmp1219 = 32'sh00001020;
	assign w_sys_tmp1224 = (w_sys_tmp1225 + r_run_k_17);
	assign w_sys_tmp1225 = 32'sh000010a1;
	assign w_sys_tmp1245 = (w_sys_tmp1246 + r_run_k_17);
	assign w_sys_tmp1246 = 32'sh00001122;
	assign w_sys_tmp1251 = (w_sys_tmp1252 + r_run_k_17);
	assign w_sys_tmp1252 = 32'sh000011a3;
	assign w_sys_tmp1257 = (w_sys_tmp1258 + r_run_k_17);
	assign w_sys_tmp1258 = 32'sh00001224;
	assign w_sys_tmp1263 = (w_sys_tmp1264 + r_run_k_17);
	assign w_sys_tmp1264 = 32'sh000012a5;
	assign w_sys_tmp1269 = (w_sys_tmp1270 + r_run_k_17);
	assign w_sys_tmp1270 = 32'sh00001326;
	assign w_sys_tmp1275 = (w_sys_tmp1276 + r_run_k_17);
	assign w_sys_tmp1276 = 32'sh000013a7;
	assign w_sys_tmp1281 = (w_sys_tmp1282 + r_run_k_17);
	assign w_sys_tmp1282 = 32'sh00001428;
	assign w_sys_tmp1287 = (w_sys_tmp1288 + r_run_k_17);
	assign w_sys_tmp1288 = 32'sh000014a9;
	assign w_sys_tmp1293 = (w_sys_tmp1294 + r_run_k_17);
	assign w_sys_tmp1294 = 32'sh0000152a;
	assign w_sys_tmp1299 = (w_sys_tmp1300 + r_run_k_17);
	assign w_sys_tmp1300 = 32'sh000015ab;
	assign w_sys_tmp1305 = (w_sys_tmp1306 + r_run_k_17);
	assign w_sys_tmp1306 = 32'sh0000162c;
	assign w_sys_tmp1311 = (w_sys_tmp1312 + r_run_k_17);
	assign w_sys_tmp1312 = 32'sh000016ad;
	assign w_sys_tmp1317 = (w_sys_tmp1318 + r_run_k_17);
	assign w_sys_tmp1318 = 32'sh0000172e;
	assign w_sys_tmp1323 = (w_sys_tmp1324 + r_run_k_17);
	assign w_sys_tmp1324 = 32'sh000017af;
	assign w_sys_tmp1329 = (w_sys_tmp1330 + r_run_k_17);
	assign w_sys_tmp1330 = 32'sh00001830;
	assign w_sys_tmp1335 = (w_sys_tmp1336 + r_run_k_17);
	assign w_sys_tmp1336 = 32'sh000018b1;
	assign w_sys_tmp1341 = (w_sys_tmp1342 + r_run_k_17);
	assign w_sys_tmp1342 = 32'sh00001932;
	assign w_sys_tmp1347 = (w_sys_tmp1348 + r_run_k_17);
	assign w_sys_tmp1348 = 32'sh000019b3;
	assign w_sys_tmp1353 = (w_sys_tmp1354 + r_run_k_17);
	assign w_sys_tmp1354 = 32'sh00001a34;
	assign w_sys_tmp1359 = (w_sys_tmp1360 + r_run_k_17);
	assign w_sys_tmp1360 = 32'sh00001ab5;
	assign w_sys_tmp1365 = (w_sys_tmp1366 + r_run_k_17);
	assign w_sys_tmp1366 = 32'sh00001b36;
	assign w_sys_tmp1371 = (w_sys_tmp1372 + r_run_k_17);
	assign w_sys_tmp1372 = 32'sh00001bb7;
	assign w_sys_tmp1377 = (w_sys_tmp1378 + r_run_k_17);
	assign w_sys_tmp1378 = 32'sh00001c38;
	assign w_sys_tmp1383 = (w_sys_tmp1384 + r_run_k_17);
	assign w_sys_tmp1384 = 32'sh00001cb9;
	assign w_sys_tmp1389 = (w_sys_tmp1390 + r_run_k_17);
	assign w_sys_tmp1390 = 32'sh00001d3a;
	assign w_sys_tmp1395 = (w_sys_tmp1396 + r_run_k_17);
	assign w_sys_tmp1396 = 32'sh00001dbb;
	assign w_sys_tmp1401 = (w_sys_tmp1402 + r_run_k_17);
	assign w_sys_tmp1402 = 32'sh00001e3c;
	assign w_sys_tmp1407 = (w_sys_tmp1408 + r_run_k_17);
	assign w_sys_tmp1408 = 32'sh00001ebd;
	assign w_sys_tmp1413 = (w_sys_tmp1414 + r_run_k_17);
	assign w_sys_tmp1414 = 32'sh00001f3e;
	assign w_sys_tmp1419 = (w_sys_tmp1420 + r_run_k_17);
	assign w_sys_tmp1420 = 32'sh00001fbf;
	assign w_sys_tmp1425 = (w_sys_tmp1426 + r_run_k_17);
	assign w_sys_tmp1426 = 32'sh00002040;
	assign w_sys_tmp1431 = (w_sys_tmp1432 + r_run_k_17);
	assign w_sys_tmp1432 = 32'sh000020c1;
	assign w_sys_tmp1449 = (w_sys_tmp1450 + r_run_k_17);
	assign w_sys_tmp1450 = 32'sh00002142;
	assign w_sys_tmp1455 = (w_sys_tmp1456 + r_run_k_17);
	assign w_sys_tmp1456 = 32'sh000021c3;
	assign w_sys_tmp1461 = (w_sys_tmp1462 + r_run_k_17);
	assign w_sys_tmp1462 = 32'sh00002244;
	assign w_sys_tmp1467 = (w_sys_tmp1468 + r_run_k_17);
	assign w_sys_tmp1468 = 32'sh000022c5;
	assign w_sys_tmp1473 = (w_sys_tmp1474 + r_run_k_17);
	assign w_sys_tmp1474 = 32'sh00002346;
	assign w_sys_tmp1479 = (w_sys_tmp1480 + r_run_k_17);
	assign w_sys_tmp1480 = 32'sh000023c7;
	assign w_sys_tmp1485 = (w_sys_tmp1486 + r_run_k_17);
	assign w_sys_tmp1486 = 32'sh00002448;
	assign w_sys_tmp1491 = (w_sys_tmp1492 + r_run_k_17);
	assign w_sys_tmp1492 = 32'sh000024c9;
	assign w_sys_tmp1497 = (w_sys_tmp1498 + r_run_k_17);
	assign w_sys_tmp1498 = 32'sh0000254a;
	assign w_sys_tmp1503 = (w_sys_tmp1504 + r_run_k_17);
	assign w_sys_tmp1504 = 32'sh000025cb;
	assign w_sys_tmp1509 = (w_sys_tmp1510 + r_run_k_17);
	assign w_sys_tmp1510 = 32'sh0000264c;
	assign w_sys_tmp1515 = (w_sys_tmp1516 + r_run_k_17);
	assign w_sys_tmp1516 = 32'sh000026cd;
	assign w_sys_tmp1521 = (w_sys_tmp1522 + r_run_k_17);
	assign w_sys_tmp1522 = 32'sh0000274e;
	assign w_sys_tmp1527 = (w_sys_tmp1528 + r_run_k_17);
	assign w_sys_tmp1528 = 32'sh000027cf;
	assign w_sys_tmp1533 = (w_sys_tmp1534 + r_run_k_17);
	assign w_sys_tmp1534 = 32'sh00002850;
	assign w_sys_tmp1539 = (w_sys_tmp1540 + r_run_k_17);
	assign w_sys_tmp1540 = 32'sh000028d1;
	assign w_sys_tmp1545 = (w_sys_tmp1546 + r_run_k_17);
	assign w_sys_tmp1546 = 32'sh00002952;
	assign w_sys_tmp1551 = (w_sys_tmp1552 + r_run_k_17);
	assign w_sys_tmp1552 = 32'sh000029d3;
	assign w_sys_tmp1557 = (w_sys_tmp1558 + r_run_k_17);
	assign w_sys_tmp1558 = 32'sh00002a54;
	assign w_sys_tmp1563 = (w_sys_tmp1564 + r_run_k_17);
	assign w_sys_tmp1564 = 32'sh00002ad5;
	assign w_sys_tmp1569 = (w_sys_tmp1570 + r_run_k_17);
	assign w_sys_tmp1570 = 32'sh00002b56;
	assign w_sys_tmp1575 = (w_sys_tmp1576 + r_run_k_17);
	assign w_sys_tmp1576 = 32'sh00002bd7;
	assign w_sys_tmp1581 = (w_sys_tmp1582 + r_run_k_17);
	assign w_sys_tmp1582 = 32'sh00002c58;
	assign w_sys_tmp1587 = (w_sys_tmp1588 + r_run_k_17);
	assign w_sys_tmp1588 = 32'sh00002cd9;
	assign w_sys_tmp1593 = (w_sys_tmp1594 + r_run_k_17);
	assign w_sys_tmp1594 = 32'sh00002d5a;
	assign w_sys_tmp1599 = (w_sys_tmp1600 + r_run_k_17);
	assign w_sys_tmp1600 = 32'sh00002ddb;
	assign w_sys_tmp1605 = (w_sys_tmp1606 + r_run_k_17);
	assign w_sys_tmp1606 = 32'sh00002e5c;
	assign w_sys_tmp1611 = (w_sys_tmp1612 + r_run_k_17);
	assign w_sys_tmp1612 = 32'sh00002edd;
	assign w_sys_tmp1617 = (w_sys_tmp1618 + r_run_k_17);
	assign w_sys_tmp1618 = 32'sh00002f5e;
	assign w_sys_tmp1623 = (w_sys_tmp1624 + r_run_k_17);
	assign w_sys_tmp1624 = 32'sh00002fdf;
	assign w_sys_tmp1629 = (w_sys_tmp1630 + r_run_k_17);
	assign w_sys_tmp1630 = 32'sh00003060;
	assign w_sys_tmp1635 = (w_sys_tmp1636 + r_run_k_17);
	assign w_sys_tmp1636 = 32'sh000030e1;
	assign w_sys_tmp1653 = (w_sys_tmp1654 + r_run_k_17);
	assign w_sys_tmp1654 = 32'sh00003162;
	assign w_sys_tmp1659 = (w_sys_tmp1660 + r_run_k_17);
	assign w_sys_tmp1660 = 32'sh000031e3;
	assign w_sys_tmp1665 = (w_sys_tmp1666 + r_run_k_17);
	assign w_sys_tmp1666 = 32'sh00003264;
	assign w_sys_tmp1671 = (w_sys_tmp1672 + r_run_k_17);
	assign w_sys_tmp1672 = 32'sh000032e5;
	assign w_sys_tmp1677 = (w_sys_tmp1678 + r_run_k_17);
	assign w_sys_tmp1678 = 32'sh00003366;
	assign w_sys_tmp1683 = (w_sys_tmp1684 + r_run_k_17);
	assign w_sys_tmp1684 = 32'sh000033e7;
	assign w_sys_tmp1689 = (w_sys_tmp1690 + r_run_k_17);
	assign w_sys_tmp1690 = 32'sh00003468;
	assign w_sys_tmp1695 = (w_sys_tmp1696 + r_run_k_17);
	assign w_sys_tmp1696 = 32'sh000034e9;
	assign w_sys_tmp1701 = (w_sys_tmp1702 + r_run_k_17);
	assign w_sys_tmp1702 = 32'sh0000356a;
	assign w_sys_tmp1707 = (w_sys_tmp1708 + r_run_k_17);
	assign w_sys_tmp1708 = 32'sh000035eb;
	assign w_sys_tmp1713 = (w_sys_tmp1714 + r_run_k_17);
	assign w_sys_tmp1714 = 32'sh0000366c;
	assign w_sys_tmp1719 = (w_sys_tmp1720 + r_run_k_17);
	assign w_sys_tmp1720 = 32'sh000036ed;
	assign w_sys_tmp1725 = (w_sys_tmp1726 + r_run_k_17);
	assign w_sys_tmp1726 = 32'sh0000376e;
	assign w_sys_tmp1731 = (w_sys_tmp1732 + r_run_k_17);
	assign w_sys_tmp1732 = 32'sh000037ef;
	assign w_sys_tmp1737 = (w_sys_tmp1738 + r_run_k_17);
	assign w_sys_tmp1738 = 32'sh00003870;
	assign w_sys_tmp1743 = (w_sys_tmp1744 + r_run_k_17);
	assign w_sys_tmp1744 = 32'sh000038f1;
	assign w_sys_tmp1749 = (w_sys_tmp1750 + r_run_k_17);
	assign w_sys_tmp1750 = 32'sh00003972;
	assign w_sys_tmp1755 = (w_sys_tmp1756 + r_run_k_17);
	assign w_sys_tmp1756 = 32'sh000039f3;
	assign w_sys_tmp1761 = (w_sys_tmp1762 + r_run_k_17);
	assign w_sys_tmp1762 = 32'sh00003a74;
	assign w_sys_tmp1767 = (w_sys_tmp1768 + r_run_k_17);
	assign w_sys_tmp1768 = 32'sh00003af5;
	assign w_sys_tmp1773 = (w_sys_tmp1774 + r_run_k_17);
	assign w_sys_tmp1774 = 32'sh00003b76;
	assign w_sys_tmp1779 = (w_sys_tmp1780 + r_run_k_17);
	assign w_sys_tmp1780 = 32'sh00003bf7;
	assign w_sys_tmp1785 = (w_sys_tmp1786 + r_run_k_17);
	assign w_sys_tmp1786 = 32'sh00003c78;
	assign w_sys_tmp1791 = (w_sys_tmp1792 + r_run_k_17);
	assign w_sys_tmp1792 = 32'sh00003cf9;
	assign w_sys_tmp1797 = (w_sys_tmp1798 + r_run_k_17);
	assign w_sys_tmp1798 = 32'sh00003d7a;
	assign w_sys_tmp1803 = (w_sys_tmp1804 + r_run_k_17);
	assign w_sys_tmp1804 = 32'sh00003dfb;
	assign w_sys_tmp1809 = (w_sys_tmp1810 + r_run_k_17);
	assign w_sys_tmp1810 = 32'sh00003e7c;
	assign w_sys_tmp1815 = (w_sys_tmp1816 + r_run_k_17);
	assign w_sys_tmp1816 = 32'sh00003efd;
	assign w_sys_tmp1821 = (w_sys_tmp1822 + r_run_k_17);
	assign w_sys_tmp1822 = 32'sh00003f7e;
	assign w_sys_tmp1827 = (w_sys_tmp1828 + r_run_k_17);
	assign w_sys_tmp1828 = 32'sh00003fff;
	assign w_sys_tmp1833 = (w_sys_tmp1834 + r_run_k_17);
	assign w_sys_tmp1834 = 32'sh00004080;
	assign w_sys_tmp1839 = (w_sys_tmp1840 + r_run_k_17);
	assign w_sys_tmp1840 = 32'sh00004101;
	assign w_sys_tmp1842 = (w_sys_tmp1843 + r_run_k_17);
	assign w_sys_tmp1843 = 32'sh000000a1;
	assign w_sys_tmp1848 = (w_sys_tmp1849 + r_run_k_17);
	assign w_sys_tmp1849 = 32'sh00000122;
	assign w_sys_tmp1854 = (w_sys_tmp1855 + r_run_k_17);
	assign w_sys_tmp1855 = 32'sh000001a3;
	assign w_sys_tmp1860 = (w_sys_tmp1861 + r_run_k_17);
	assign w_sys_tmp1861 = 32'sh00000224;
	assign w_sys_tmp1866 = (w_sys_tmp1867 + r_run_k_17);
	assign w_sys_tmp1867 = 32'sh000002a5;
	assign w_sys_tmp1872 = (w_sys_tmp1873 + r_run_k_17);
	assign w_sys_tmp1873 = 32'sh00000326;
	assign w_sys_tmp1878 = (w_sys_tmp1879 + r_run_k_17);
	assign w_sys_tmp1879 = 32'sh000003a7;
	assign w_sys_tmp1884 = (w_sys_tmp1885 + r_run_k_17);
	assign w_sys_tmp1885 = 32'sh00000428;
	assign w_sys_tmp1890 = (w_sys_tmp1891 + r_run_k_17);
	assign w_sys_tmp1891 = 32'sh000004a9;
	assign w_sys_tmp1896 = (w_sys_tmp1897 + r_run_k_17);
	assign w_sys_tmp1897 = 32'sh0000052a;
	assign w_sys_tmp1902 = (w_sys_tmp1903 + r_run_k_17);
	assign w_sys_tmp1903 = 32'sh000005ab;
	assign w_sys_tmp1908 = (w_sys_tmp1909 + r_run_k_17);
	assign w_sys_tmp1909 = 32'sh0000062c;
	assign w_sys_tmp1914 = (w_sys_tmp1915 + r_run_k_17);
	assign w_sys_tmp1915 = 32'sh000006ad;
	assign w_sys_tmp1920 = (w_sys_tmp1921 + r_run_k_17);
	assign w_sys_tmp1921 = 32'sh0000072e;
	assign w_sys_tmp1926 = (w_sys_tmp1927 + r_run_k_17);
	assign w_sys_tmp1927 = 32'sh000007af;
	assign w_sys_tmp1932 = (w_sys_tmp1933 + r_run_k_17);
	assign w_sys_tmp1933 = 32'sh00000830;
	assign w_sys_tmp1938 = (w_sys_tmp1939 + r_run_k_17);
	assign w_sys_tmp1939 = 32'sh000008b1;
	assign w_sys_tmp1944 = (w_sys_tmp1945 + r_run_k_17);
	assign w_sys_tmp1945 = 32'sh00000932;
	assign w_sys_tmp1950 = (w_sys_tmp1951 + r_run_k_17);
	assign w_sys_tmp1951 = 32'sh000009b3;
	assign w_sys_tmp1956 = (w_sys_tmp1957 + r_run_k_17);
	assign w_sys_tmp1957 = 32'sh00000a34;
	assign w_sys_tmp1962 = (w_sys_tmp1963 + r_run_k_17);
	assign w_sys_tmp1963 = 32'sh00000ab5;
	assign w_sys_tmp1968 = (w_sys_tmp1969 + r_run_k_17);
	assign w_sys_tmp1969 = 32'sh00000b36;
	assign w_sys_tmp1974 = (w_sys_tmp1975 + r_run_k_17);
	assign w_sys_tmp1975 = 32'sh00000bb7;
	assign w_sys_tmp1980 = (w_sys_tmp1981 + r_run_k_17);
	assign w_sys_tmp1981 = 32'sh00000c38;
	assign w_sys_tmp1986 = (w_sys_tmp1987 + r_run_k_17);
	assign w_sys_tmp1987 = 32'sh00000cb9;
	assign w_sys_tmp1992 = (w_sys_tmp1993 + r_run_k_17);
	assign w_sys_tmp1993 = 32'sh00000d3a;
	assign w_sys_tmp1998 = (w_sys_tmp1999 + r_run_k_17);
	assign w_sys_tmp1999 = 32'sh00000dbb;
	assign w_sys_tmp2004 = (w_sys_tmp2005 + r_run_k_17);
	assign w_sys_tmp2005 = 32'sh00000e3c;
	assign w_sys_tmp2010 = (w_sys_tmp2011 + r_run_k_17);
	assign w_sys_tmp2011 = 32'sh00000ebd;
	assign w_sys_tmp2016 = (w_sys_tmp2017 + r_run_k_17);
	assign w_sys_tmp2017 = 32'sh00000f3e;
	assign w_sys_tmp2022 = (w_sys_tmp2023 + r_run_k_17);
	assign w_sys_tmp2023 = 32'sh00000fbf;
	assign w_sys_tmp2028 = (w_sys_tmp2029 + r_run_k_17);
	assign w_sys_tmp2029 = 32'sh00001040;
	assign w_sys_tmp2034 = (w_sys_tmp2035 + r_run_k_17);
	assign w_sys_tmp2035 = 32'sh000010c1;
	assign w_sys_tmp2055 = (w_sys_tmp2056 + r_run_k_17);
	assign w_sys_tmp2056 = 32'sh00001142;
	assign w_sys_tmp2061 = (w_sys_tmp2062 + r_run_k_17);
	assign w_sys_tmp2062 = 32'sh000011c3;
	assign w_sys_tmp2067 = (w_sys_tmp2068 + r_run_k_17);
	assign w_sys_tmp2068 = 32'sh00001244;
	assign w_sys_tmp2073 = (w_sys_tmp2074 + r_run_k_17);
	assign w_sys_tmp2074 = 32'sh000012c5;
	assign w_sys_tmp2079 = (w_sys_tmp2080 + r_run_k_17);
	assign w_sys_tmp2080 = 32'sh00001346;
	assign w_sys_tmp2085 = (w_sys_tmp2086 + r_run_k_17);
	assign w_sys_tmp2086 = 32'sh000013c7;
	assign w_sys_tmp2091 = (w_sys_tmp2092 + r_run_k_17);
	assign w_sys_tmp2092 = 32'sh00001448;
	assign w_sys_tmp2097 = (w_sys_tmp2098 + r_run_k_17);
	assign w_sys_tmp2098 = 32'sh000014c9;
	assign w_sys_tmp2103 = (w_sys_tmp2104 + r_run_k_17);
	assign w_sys_tmp2104 = 32'sh0000154a;
	assign w_sys_tmp2109 = (w_sys_tmp2110 + r_run_k_17);
	assign w_sys_tmp2110 = 32'sh000015cb;
	assign w_sys_tmp2115 = (w_sys_tmp2116 + r_run_k_17);
	assign w_sys_tmp2116 = 32'sh0000164c;
	assign w_sys_tmp2121 = (w_sys_tmp2122 + r_run_k_17);
	assign w_sys_tmp2122 = 32'sh000016cd;
	assign w_sys_tmp2127 = (w_sys_tmp2128 + r_run_k_17);
	assign w_sys_tmp2128 = 32'sh0000174e;
	assign w_sys_tmp2133 = (w_sys_tmp2134 + r_run_k_17);
	assign w_sys_tmp2134 = 32'sh000017cf;
	assign w_sys_tmp2139 = (w_sys_tmp2140 + r_run_k_17);
	assign w_sys_tmp2140 = 32'sh00001850;
	assign w_sys_tmp2145 = (w_sys_tmp2146 + r_run_k_17);
	assign w_sys_tmp2146 = 32'sh000018d1;
	assign w_sys_tmp2151 = (w_sys_tmp2152 + r_run_k_17);
	assign w_sys_tmp2152 = 32'sh00001952;
	assign w_sys_tmp2157 = (w_sys_tmp2158 + r_run_k_17);
	assign w_sys_tmp2158 = 32'sh000019d3;
	assign w_sys_tmp2163 = (w_sys_tmp2164 + r_run_k_17);
	assign w_sys_tmp2164 = 32'sh00001a54;
	assign w_sys_tmp2169 = (w_sys_tmp2170 + r_run_k_17);
	assign w_sys_tmp2170 = 32'sh00001ad5;
	assign w_sys_tmp2175 = (w_sys_tmp2176 + r_run_k_17);
	assign w_sys_tmp2176 = 32'sh00001b56;
	assign w_sys_tmp2181 = (w_sys_tmp2182 + r_run_k_17);
	assign w_sys_tmp2182 = 32'sh00001bd7;
	assign w_sys_tmp2187 = (w_sys_tmp2188 + r_run_k_17);
	assign w_sys_tmp2188 = 32'sh00001c58;
	assign w_sys_tmp2193 = (w_sys_tmp2194 + r_run_k_17);
	assign w_sys_tmp2194 = 32'sh00001cd9;
	assign w_sys_tmp2199 = (w_sys_tmp2200 + r_run_k_17);
	assign w_sys_tmp2200 = 32'sh00001d5a;
	assign w_sys_tmp2205 = (w_sys_tmp2206 + r_run_k_17);
	assign w_sys_tmp2206 = 32'sh00001ddb;
	assign w_sys_tmp2211 = (w_sys_tmp2212 + r_run_k_17);
	assign w_sys_tmp2212 = 32'sh00001e5c;
	assign w_sys_tmp2217 = (w_sys_tmp2218 + r_run_k_17);
	assign w_sys_tmp2218 = 32'sh00001edd;
	assign w_sys_tmp2223 = (w_sys_tmp2224 + r_run_k_17);
	assign w_sys_tmp2224 = 32'sh00001f5e;
	assign w_sys_tmp2229 = (w_sys_tmp2230 + r_run_k_17);
	assign w_sys_tmp2230 = 32'sh00001fdf;
	assign w_sys_tmp2235 = (w_sys_tmp2236 + r_run_k_17);
	assign w_sys_tmp2236 = 32'sh00002060;
	assign w_sys_tmp2241 = (w_sys_tmp2242 + r_run_k_17);
	assign w_sys_tmp2242 = 32'sh000020e1;
	assign w_sys_tmp2259 = (w_sys_tmp2260 + r_run_k_17);
	assign w_sys_tmp2260 = 32'sh00002162;
	assign w_sys_tmp2265 = (w_sys_tmp2266 + r_run_k_17);
	assign w_sys_tmp2266 = 32'sh000021e3;
	assign w_sys_tmp2271 = (w_sys_tmp2272 + r_run_k_17);
	assign w_sys_tmp2272 = 32'sh00002264;
	assign w_sys_tmp2277 = (w_sys_tmp2278 + r_run_k_17);
	assign w_sys_tmp2278 = 32'sh000022e5;
	assign w_sys_tmp2283 = (w_sys_tmp2284 + r_run_k_17);
	assign w_sys_tmp2284 = 32'sh00002366;
	assign w_sys_tmp2289 = (w_sys_tmp2290 + r_run_k_17);
	assign w_sys_tmp2290 = 32'sh000023e7;
	assign w_sys_tmp2295 = (w_sys_tmp2296 + r_run_k_17);
	assign w_sys_tmp2296 = 32'sh00002468;
	assign w_sys_tmp2301 = (w_sys_tmp2302 + r_run_k_17);
	assign w_sys_tmp2302 = 32'sh000024e9;
	assign w_sys_tmp2307 = (w_sys_tmp2308 + r_run_k_17);
	assign w_sys_tmp2308 = 32'sh0000256a;
	assign w_sys_tmp2313 = (w_sys_tmp2314 + r_run_k_17);
	assign w_sys_tmp2314 = 32'sh000025eb;
	assign w_sys_tmp2319 = (w_sys_tmp2320 + r_run_k_17);
	assign w_sys_tmp2320 = 32'sh0000266c;
	assign w_sys_tmp2325 = (w_sys_tmp2326 + r_run_k_17);
	assign w_sys_tmp2326 = 32'sh000026ed;
	assign w_sys_tmp2331 = (w_sys_tmp2332 + r_run_k_17);
	assign w_sys_tmp2332 = 32'sh0000276e;
	assign w_sys_tmp2337 = (w_sys_tmp2338 + r_run_k_17);
	assign w_sys_tmp2338 = 32'sh000027ef;
	assign w_sys_tmp2343 = (w_sys_tmp2344 + r_run_k_17);
	assign w_sys_tmp2344 = 32'sh00002870;
	assign w_sys_tmp2349 = (w_sys_tmp2350 + r_run_k_17);
	assign w_sys_tmp2350 = 32'sh000028f1;
	assign w_sys_tmp2355 = (w_sys_tmp2356 + r_run_k_17);
	assign w_sys_tmp2356 = 32'sh00002972;
	assign w_sys_tmp2361 = (w_sys_tmp2362 + r_run_k_17);
	assign w_sys_tmp2362 = 32'sh000029f3;
	assign w_sys_tmp2367 = (w_sys_tmp2368 + r_run_k_17);
	assign w_sys_tmp2368 = 32'sh00002a74;
	assign w_sys_tmp2373 = (w_sys_tmp2374 + r_run_k_17);
	assign w_sys_tmp2374 = 32'sh00002af5;
	assign w_sys_tmp2379 = (w_sys_tmp2380 + r_run_k_17);
	assign w_sys_tmp2380 = 32'sh00002b76;
	assign w_sys_tmp2385 = (w_sys_tmp2386 + r_run_k_17);
	assign w_sys_tmp2386 = 32'sh00002bf7;
	assign w_sys_tmp2391 = (w_sys_tmp2392 + r_run_k_17);
	assign w_sys_tmp2392 = 32'sh00002c78;
	assign w_sys_tmp2397 = (w_sys_tmp2398 + r_run_k_17);
	assign w_sys_tmp2398 = 32'sh00002cf9;
	assign w_sys_tmp2403 = (w_sys_tmp2404 + r_run_k_17);
	assign w_sys_tmp2404 = 32'sh00002d7a;
	assign w_sys_tmp2409 = (w_sys_tmp2410 + r_run_k_17);
	assign w_sys_tmp2410 = 32'sh00002dfb;
	assign w_sys_tmp2415 = (w_sys_tmp2416 + r_run_k_17);
	assign w_sys_tmp2416 = 32'sh00002e7c;
	assign w_sys_tmp2421 = (w_sys_tmp2422 + r_run_k_17);
	assign w_sys_tmp2422 = 32'sh00002efd;
	assign w_sys_tmp2427 = (w_sys_tmp2428 + r_run_k_17);
	assign w_sys_tmp2428 = 32'sh00002f7e;
	assign w_sys_tmp2433 = (w_sys_tmp2434 + r_run_k_17);
	assign w_sys_tmp2434 = 32'sh00002fff;
	assign w_sys_tmp2439 = (w_sys_tmp2440 + r_run_k_17);
	assign w_sys_tmp2440 = 32'sh00003080;
	assign w_sys_tmp2445 = (w_sys_tmp2446 + r_run_k_17);
	assign w_sys_tmp2446 = 32'sh00003101;
	assign w_sys_tmp2463 = (w_sys_tmp2464 + r_run_k_17);
	assign w_sys_tmp2464 = 32'sh00003182;
	assign w_sys_tmp2469 = (w_sys_tmp2470 + r_run_k_17);
	assign w_sys_tmp2470 = 32'sh00003203;
	assign w_sys_tmp2475 = (w_sys_tmp2476 + r_run_k_17);
	assign w_sys_tmp2476 = 32'sh00003284;
	assign w_sys_tmp2481 = (w_sys_tmp2482 + r_run_k_17);
	assign w_sys_tmp2482 = 32'sh00003305;
	assign w_sys_tmp2487 = (w_sys_tmp2488 + r_run_k_17);
	assign w_sys_tmp2488 = 32'sh00003386;
	assign w_sys_tmp2493 = (w_sys_tmp2494 + r_run_k_17);
	assign w_sys_tmp2494 = 32'sh00003407;
	assign w_sys_tmp2499 = (w_sys_tmp2500 + r_run_k_17);
	assign w_sys_tmp2500 = 32'sh00003488;
	assign w_sys_tmp2505 = (w_sys_tmp2506 + r_run_k_17);
	assign w_sys_tmp2506 = 32'sh00003509;
	assign w_sys_tmp2511 = (w_sys_tmp2512 + r_run_k_17);
	assign w_sys_tmp2512 = 32'sh0000358a;
	assign w_sys_tmp2517 = (w_sys_tmp2518 + r_run_k_17);
	assign w_sys_tmp2518 = 32'sh0000360b;
	assign w_sys_tmp2523 = (w_sys_tmp2524 + r_run_k_17);
	assign w_sys_tmp2524 = 32'sh0000368c;
	assign w_sys_tmp2529 = (w_sys_tmp2530 + r_run_k_17);
	assign w_sys_tmp2530 = 32'sh0000370d;
	assign w_sys_tmp2535 = (w_sys_tmp2536 + r_run_k_17);
	assign w_sys_tmp2536 = 32'sh0000378e;
	assign w_sys_tmp2541 = (w_sys_tmp2542 + r_run_k_17);
	assign w_sys_tmp2542 = 32'sh0000380f;
	assign w_sys_tmp2547 = (w_sys_tmp2548 + r_run_k_17);
	assign w_sys_tmp2548 = 32'sh00003890;
	assign w_sys_tmp2553 = (w_sys_tmp2554 + r_run_k_17);
	assign w_sys_tmp2554 = 32'sh00003911;
	assign w_sys_tmp2559 = (w_sys_tmp2560 + r_run_k_17);
	assign w_sys_tmp2560 = 32'sh00003992;
	assign w_sys_tmp2565 = (w_sys_tmp2566 + r_run_k_17);
	assign w_sys_tmp2566 = 32'sh00003a13;
	assign w_sys_tmp2571 = (w_sys_tmp2572 + r_run_k_17);
	assign w_sys_tmp2572 = 32'sh00003a94;
	assign w_sys_tmp2577 = (w_sys_tmp2578 + r_run_k_17);
	assign w_sys_tmp2578 = 32'sh00003b15;
	assign w_sys_tmp2583 = (w_sys_tmp2584 + r_run_k_17);
	assign w_sys_tmp2584 = 32'sh00003b96;
	assign w_sys_tmp2589 = (w_sys_tmp2590 + r_run_k_17);
	assign w_sys_tmp2590 = 32'sh00003c17;
	assign w_sys_tmp2595 = (w_sys_tmp2596 + r_run_k_17);
	assign w_sys_tmp2596 = 32'sh00003c98;
	assign w_sys_tmp2601 = (w_sys_tmp2602 + r_run_k_17);
	assign w_sys_tmp2602 = 32'sh00003d19;
	assign w_sys_tmp2607 = (w_sys_tmp2608 + r_run_k_17);
	assign w_sys_tmp2608 = 32'sh00003d9a;
	assign w_sys_tmp2613 = (w_sys_tmp2614 + r_run_k_17);
	assign w_sys_tmp2614 = 32'sh00003e1b;
	assign w_sys_tmp2619 = (w_sys_tmp2620 + r_run_k_17);
	assign w_sys_tmp2620 = 32'sh00003e9c;
	assign w_sys_tmp2625 = (w_sys_tmp2626 + r_run_k_17);
	assign w_sys_tmp2626 = 32'sh00003f1d;
	assign w_sys_tmp2631 = (w_sys_tmp2632 + r_run_k_17);
	assign w_sys_tmp2632 = 32'sh00003f9e;
	assign w_sys_tmp2637 = (w_sys_tmp2638 + r_run_k_17);
	assign w_sys_tmp2638 = 32'sh0000401f;
	assign w_sys_tmp2643 = (w_sys_tmp2644 + r_run_k_17);
	assign w_sys_tmp2644 = 32'sh000040a0;
	assign w_sys_tmp2649 = (w_sys_tmp2650 + r_run_k_17);
	assign w_sys_tmp2650 = 32'sh00004121;
	assign w_sys_tmp2652 = (w_sys_tmp2653 + r_run_k_17);
	assign w_sys_tmp2653 = 32'sh000000c1;
	assign w_sys_tmp2658 = (w_sys_tmp2659 + r_run_k_17);
	assign w_sys_tmp2659 = 32'sh00000142;
	assign w_sys_tmp2664 = (w_sys_tmp2665 + r_run_k_17);
	assign w_sys_tmp2665 = 32'sh000001c3;
	assign w_sys_tmp2670 = (w_sys_tmp2671 + r_run_k_17);
	assign w_sys_tmp2671 = 32'sh00000244;
	assign w_sys_tmp2676 = (w_sys_tmp2677 + r_run_k_17);
	assign w_sys_tmp2677 = 32'sh000002c5;
	assign w_sys_tmp2682 = (w_sys_tmp2683 + r_run_k_17);
	assign w_sys_tmp2683 = 32'sh00000346;
	assign w_sys_tmp2688 = (w_sys_tmp2689 + r_run_k_17);
	assign w_sys_tmp2689 = 32'sh000003c7;
	assign w_sys_tmp2694 = (w_sys_tmp2695 + r_run_k_17);
	assign w_sys_tmp2695 = 32'sh00000448;
	assign w_sys_tmp2700 = (w_sys_tmp2701 + r_run_k_17);
	assign w_sys_tmp2701 = 32'sh000004c9;
	assign w_sys_tmp2706 = (w_sys_tmp2707 + r_run_k_17);
	assign w_sys_tmp2707 = 32'sh0000054a;
	assign w_sys_tmp2712 = (w_sys_tmp2713 + r_run_k_17);
	assign w_sys_tmp2713 = 32'sh000005cb;
	assign w_sys_tmp2718 = (w_sys_tmp2719 + r_run_k_17);
	assign w_sys_tmp2719 = 32'sh0000064c;
	assign w_sys_tmp2724 = (w_sys_tmp2725 + r_run_k_17);
	assign w_sys_tmp2725 = 32'sh000006cd;
	assign w_sys_tmp2730 = (w_sys_tmp2731 + r_run_k_17);
	assign w_sys_tmp2731 = 32'sh0000074e;
	assign w_sys_tmp2736 = (w_sys_tmp2737 + r_run_k_17);
	assign w_sys_tmp2737 = 32'sh000007cf;
	assign w_sys_tmp2742 = (w_sys_tmp2743 + r_run_k_17);
	assign w_sys_tmp2743 = 32'sh00000850;
	assign w_sys_tmp2748 = (w_sys_tmp2749 + r_run_k_17);
	assign w_sys_tmp2749 = 32'sh000008d1;
	assign w_sys_tmp2754 = (w_sys_tmp2755 + r_run_k_17);
	assign w_sys_tmp2755 = 32'sh00000952;
	assign w_sys_tmp2760 = (w_sys_tmp2761 + r_run_k_17);
	assign w_sys_tmp2761 = 32'sh000009d3;
	assign w_sys_tmp2766 = (w_sys_tmp2767 + r_run_k_17);
	assign w_sys_tmp2767 = 32'sh00000a54;
	assign w_sys_tmp2772 = (w_sys_tmp2773 + r_run_k_17);
	assign w_sys_tmp2773 = 32'sh00000ad5;
	assign w_sys_tmp2778 = (w_sys_tmp2779 + r_run_k_17);
	assign w_sys_tmp2779 = 32'sh00000b56;
	assign w_sys_tmp2784 = (w_sys_tmp2785 + r_run_k_17);
	assign w_sys_tmp2785 = 32'sh00000bd7;
	assign w_sys_tmp2790 = (w_sys_tmp2791 + r_run_k_17);
	assign w_sys_tmp2791 = 32'sh00000c58;
	assign w_sys_tmp2796 = (w_sys_tmp2797 + r_run_k_17);
	assign w_sys_tmp2797 = 32'sh00000cd9;
	assign w_sys_tmp2802 = (w_sys_tmp2803 + r_run_k_17);
	assign w_sys_tmp2803 = 32'sh00000d5a;
	assign w_sys_tmp2808 = (w_sys_tmp2809 + r_run_k_17);
	assign w_sys_tmp2809 = 32'sh00000ddb;
	assign w_sys_tmp2814 = (w_sys_tmp2815 + r_run_k_17);
	assign w_sys_tmp2815 = 32'sh00000e5c;
	assign w_sys_tmp2820 = (w_sys_tmp2821 + r_run_k_17);
	assign w_sys_tmp2821 = 32'sh00000edd;
	assign w_sys_tmp2826 = (w_sys_tmp2827 + r_run_k_17);
	assign w_sys_tmp2827 = 32'sh00000f5e;
	assign w_sys_tmp2832 = (w_sys_tmp2833 + r_run_k_17);
	assign w_sys_tmp2833 = 32'sh00000fdf;
	assign w_sys_tmp2838 = (w_sys_tmp2839 + r_run_k_17);
	assign w_sys_tmp2839 = 32'sh00001060;
	assign w_sys_tmp2844 = (w_sys_tmp2845 + r_run_k_17);
	assign w_sys_tmp2845 = 32'sh000010e1;
	assign w_sys_tmp2865 = (w_sys_tmp2866 + r_run_k_17);
	assign w_sys_tmp2866 = 32'sh00001162;
	assign w_sys_tmp2871 = (w_sys_tmp2872 + r_run_k_17);
	assign w_sys_tmp2872 = 32'sh000011e3;
	assign w_sys_tmp2877 = (w_sys_tmp2878 + r_run_k_17);
	assign w_sys_tmp2878 = 32'sh00001264;
	assign w_sys_tmp2883 = (w_sys_tmp2884 + r_run_k_17);
	assign w_sys_tmp2884 = 32'sh000012e5;
	assign w_sys_tmp2889 = (w_sys_tmp2890 + r_run_k_17);
	assign w_sys_tmp2890 = 32'sh00001366;
	assign w_sys_tmp2895 = (w_sys_tmp2896 + r_run_k_17);
	assign w_sys_tmp2896 = 32'sh000013e7;
	assign w_sys_tmp2901 = (w_sys_tmp2902 + r_run_k_17);
	assign w_sys_tmp2902 = 32'sh00001468;
	assign w_sys_tmp2907 = (w_sys_tmp2908 + r_run_k_17);
	assign w_sys_tmp2908 = 32'sh000014e9;
	assign w_sys_tmp2913 = (w_sys_tmp2914 + r_run_k_17);
	assign w_sys_tmp2914 = 32'sh0000156a;
	assign w_sys_tmp2919 = (w_sys_tmp2920 + r_run_k_17);
	assign w_sys_tmp2920 = 32'sh000015eb;
	assign w_sys_tmp2925 = (w_sys_tmp2926 + r_run_k_17);
	assign w_sys_tmp2926 = 32'sh0000166c;
	assign w_sys_tmp2931 = (w_sys_tmp2932 + r_run_k_17);
	assign w_sys_tmp2932 = 32'sh000016ed;
	assign w_sys_tmp2937 = (w_sys_tmp2938 + r_run_k_17);
	assign w_sys_tmp2938 = 32'sh0000176e;
	assign w_sys_tmp2943 = (w_sys_tmp2944 + r_run_k_17);
	assign w_sys_tmp2944 = 32'sh000017ef;
	assign w_sys_tmp2949 = (w_sys_tmp2950 + r_run_k_17);
	assign w_sys_tmp2950 = 32'sh00001870;
	assign w_sys_tmp2955 = (w_sys_tmp2956 + r_run_k_17);
	assign w_sys_tmp2956 = 32'sh000018f1;
	assign w_sys_tmp2961 = (w_sys_tmp2962 + r_run_k_17);
	assign w_sys_tmp2962 = 32'sh00001972;
	assign w_sys_tmp2967 = (w_sys_tmp2968 + r_run_k_17);
	assign w_sys_tmp2968 = 32'sh000019f3;
	assign w_sys_tmp2973 = (w_sys_tmp2974 + r_run_k_17);
	assign w_sys_tmp2974 = 32'sh00001a74;
	assign w_sys_tmp2979 = (w_sys_tmp2980 + r_run_k_17);
	assign w_sys_tmp2980 = 32'sh00001af5;
	assign w_sys_tmp2985 = (w_sys_tmp2986 + r_run_k_17);
	assign w_sys_tmp2986 = 32'sh00001b76;
	assign w_sys_tmp2991 = (w_sys_tmp2992 + r_run_k_17);
	assign w_sys_tmp2992 = 32'sh00001bf7;
	assign w_sys_tmp2997 = (w_sys_tmp2998 + r_run_k_17);
	assign w_sys_tmp2998 = 32'sh00001c78;
	assign w_sys_tmp3003 = (w_sys_tmp3004 + r_run_k_17);
	assign w_sys_tmp3004 = 32'sh00001cf9;
	assign w_sys_tmp3009 = (w_sys_tmp3010 + r_run_k_17);
	assign w_sys_tmp3010 = 32'sh00001d7a;
	assign w_sys_tmp3015 = (w_sys_tmp3016 + r_run_k_17);
	assign w_sys_tmp3016 = 32'sh00001dfb;
	assign w_sys_tmp3021 = (w_sys_tmp3022 + r_run_k_17);
	assign w_sys_tmp3022 = 32'sh00001e7c;
	assign w_sys_tmp3027 = (w_sys_tmp3028 + r_run_k_17);
	assign w_sys_tmp3028 = 32'sh00001efd;
	assign w_sys_tmp3033 = (w_sys_tmp3034 + r_run_k_17);
	assign w_sys_tmp3034 = 32'sh00001f7e;
	assign w_sys_tmp3039 = (w_sys_tmp3040 + r_run_k_17);
	assign w_sys_tmp3040 = 32'sh00001fff;
	assign w_sys_tmp3045 = (w_sys_tmp3046 + r_run_k_17);
	assign w_sys_tmp3046 = 32'sh00002080;
	assign w_sys_tmp3051 = (w_sys_tmp3052 + r_run_k_17);
	assign w_sys_tmp3052 = 32'sh00002101;
	assign w_sys_tmp3069 = (w_sys_tmp3070 + r_run_k_17);
	assign w_sys_tmp3070 = 32'sh00002182;
	assign w_sys_tmp3075 = (w_sys_tmp3076 + r_run_k_17);
	assign w_sys_tmp3076 = 32'sh00002203;
	assign w_sys_tmp3081 = (w_sys_tmp3082 + r_run_k_17);
	assign w_sys_tmp3082 = 32'sh00002284;
	assign w_sys_tmp3087 = (w_sys_tmp3088 + r_run_k_17);
	assign w_sys_tmp3088 = 32'sh00002305;
	assign w_sys_tmp3093 = (w_sys_tmp3094 + r_run_k_17);
	assign w_sys_tmp3094 = 32'sh00002386;
	assign w_sys_tmp3099 = (w_sys_tmp3100 + r_run_k_17);
	assign w_sys_tmp3100 = 32'sh00002407;
	assign w_sys_tmp3105 = (w_sys_tmp3106 + r_run_k_17);
	assign w_sys_tmp3106 = 32'sh00002488;
	assign w_sys_tmp3111 = (w_sys_tmp3112 + r_run_k_17);
	assign w_sys_tmp3112 = 32'sh00002509;
	assign w_sys_tmp3117 = (w_sys_tmp3118 + r_run_k_17);
	assign w_sys_tmp3118 = 32'sh0000258a;
	assign w_sys_tmp3123 = (w_sys_tmp3124 + r_run_k_17);
	assign w_sys_tmp3124 = 32'sh0000260b;
	assign w_sys_tmp3129 = (w_sys_tmp3130 + r_run_k_17);
	assign w_sys_tmp3130 = 32'sh0000268c;
	assign w_sys_tmp3135 = (w_sys_tmp3136 + r_run_k_17);
	assign w_sys_tmp3136 = 32'sh0000270d;
	assign w_sys_tmp3141 = (w_sys_tmp3142 + r_run_k_17);
	assign w_sys_tmp3142 = 32'sh0000278e;
	assign w_sys_tmp3147 = (w_sys_tmp3148 + r_run_k_17);
	assign w_sys_tmp3148 = 32'sh0000280f;
	assign w_sys_tmp3153 = (w_sys_tmp3154 + r_run_k_17);
	assign w_sys_tmp3154 = 32'sh00002890;
	assign w_sys_tmp3159 = (w_sys_tmp3160 + r_run_k_17);
	assign w_sys_tmp3160 = 32'sh00002911;
	assign w_sys_tmp3165 = (w_sys_tmp3166 + r_run_k_17);
	assign w_sys_tmp3166 = 32'sh00002992;
	assign w_sys_tmp3171 = (w_sys_tmp3172 + r_run_k_17);
	assign w_sys_tmp3172 = 32'sh00002a13;
	assign w_sys_tmp3177 = (w_sys_tmp3178 + r_run_k_17);
	assign w_sys_tmp3178 = 32'sh00002a94;
	assign w_sys_tmp3183 = (w_sys_tmp3184 + r_run_k_17);
	assign w_sys_tmp3184 = 32'sh00002b15;
	assign w_sys_tmp3189 = (w_sys_tmp3190 + r_run_k_17);
	assign w_sys_tmp3190 = 32'sh00002b96;
	assign w_sys_tmp3195 = (w_sys_tmp3196 + r_run_k_17);
	assign w_sys_tmp3196 = 32'sh00002c17;
	assign w_sys_tmp3201 = (w_sys_tmp3202 + r_run_k_17);
	assign w_sys_tmp3202 = 32'sh00002c98;
	assign w_sys_tmp3207 = (w_sys_tmp3208 + r_run_k_17);
	assign w_sys_tmp3208 = 32'sh00002d19;
	assign w_sys_tmp3213 = (w_sys_tmp3214 + r_run_k_17);
	assign w_sys_tmp3214 = 32'sh00002d9a;
	assign w_sys_tmp3219 = (w_sys_tmp3220 + r_run_k_17);
	assign w_sys_tmp3220 = 32'sh00002e1b;
	assign w_sys_tmp3225 = (w_sys_tmp3226 + r_run_k_17);
	assign w_sys_tmp3226 = 32'sh00002e9c;
	assign w_sys_tmp3231 = (w_sys_tmp3232 + r_run_k_17);
	assign w_sys_tmp3232 = 32'sh00002f1d;
	assign w_sys_tmp3237 = (w_sys_tmp3238 + r_run_k_17);
	assign w_sys_tmp3238 = 32'sh00002f9e;
	assign w_sys_tmp3243 = (w_sys_tmp3244 + r_run_k_17);
	assign w_sys_tmp3244 = 32'sh0000301f;
	assign w_sys_tmp3249 = (w_sys_tmp3250 + r_run_k_17);
	assign w_sys_tmp3250 = 32'sh000030a0;
	assign w_sys_tmp3255 = (w_sys_tmp3256 + r_run_k_17);
	assign w_sys_tmp3256 = 32'sh00003121;
	assign w_sys_tmp3273 = (w_sys_tmp3274 + r_run_k_17);
	assign w_sys_tmp3274 = 32'sh000031a2;
	assign w_sys_tmp3279 = (w_sys_tmp3280 + r_run_k_17);
	assign w_sys_tmp3280 = 32'sh00003223;
	assign w_sys_tmp3285 = (w_sys_tmp3286 + r_run_k_17);
	assign w_sys_tmp3286 = 32'sh000032a4;
	assign w_sys_tmp3291 = (w_sys_tmp3292 + r_run_k_17);
	assign w_sys_tmp3292 = 32'sh00003325;
	assign w_sys_tmp3297 = (w_sys_tmp3298 + r_run_k_17);
	assign w_sys_tmp3298 = 32'sh000033a6;
	assign w_sys_tmp3303 = (w_sys_tmp3304 + r_run_k_17);
	assign w_sys_tmp3304 = 32'sh00003427;
	assign w_sys_tmp3309 = (w_sys_tmp3310 + r_run_k_17);
	assign w_sys_tmp3310 = 32'sh000034a8;
	assign w_sys_tmp3315 = (w_sys_tmp3316 + r_run_k_17);
	assign w_sys_tmp3316 = 32'sh00003529;
	assign w_sys_tmp3321 = (w_sys_tmp3322 + r_run_k_17);
	assign w_sys_tmp3322 = 32'sh000035aa;
	assign w_sys_tmp3327 = (w_sys_tmp3328 + r_run_k_17);
	assign w_sys_tmp3328 = 32'sh0000362b;
	assign w_sys_tmp3333 = (w_sys_tmp3334 + r_run_k_17);
	assign w_sys_tmp3334 = 32'sh000036ac;
	assign w_sys_tmp3339 = (w_sys_tmp3340 + r_run_k_17);
	assign w_sys_tmp3340 = 32'sh0000372d;
	assign w_sys_tmp3345 = (w_sys_tmp3346 + r_run_k_17);
	assign w_sys_tmp3346 = 32'sh000037ae;
	assign w_sys_tmp3351 = (w_sys_tmp3352 + r_run_k_17);
	assign w_sys_tmp3352 = 32'sh0000382f;
	assign w_sys_tmp3357 = (w_sys_tmp3358 + r_run_k_17);
	assign w_sys_tmp3358 = 32'sh000038b0;
	assign w_sys_tmp3363 = (w_sys_tmp3364 + r_run_k_17);
	assign w_sys_tmp3364 = 32'sh00003931;
	assign w_sys_tmp3369 = (w_sys_tmp3370 + r_run_k_17);
	assign w_sys_tmp3370 = 32'sh000039b2;
	assign w_sys_tmp3375 = (w_sys_tmp3376 + r_run_k_17);
	assign w_sys_tmp3376 = 32'sh00003a33;
	assign w_sys_tmp3381 = (w_sys_tmp3382 + r_run_k_17);
	assign w_sys_tmp3382 = 32'sh00003ab4;
	assign w_sys_tmp3387 = (w_sys_tmp3388 + r_run_k_17);
	assign w_sys_tmp3388 = 32'sh00003b35;
	assign w_sys_tmp3393 = (w_sys_tmp3394 + r_run_k_17);
	assign w_sys_tmp3394 = 32'sh00003bb6;
	assign w_sys_tmp3399 = (w_sys_tmp3400 + r_run_k_17);
	assign w_sys_tmp3400 = 32'sh00003c37;
	assign w_sys_tmp3405 = (w_sys_tmp3406 + r_run_k_17);
	assign w_sys_tmp3406 = 32'sh00003cb8;
	assign w_sys_tmp3411 = (w_sys_tmp3412 + r_run_k_17);
	assign w_sys_tmp3412 = 32'sh00003d39;
	assign w_sys_tmp3417 = (w_sys_tmp3418 + r_run_k_17);
	assign w_sys_tmp3418 = 32'sh00003dba;
	assign w_sys_tmp3423 = (w_sys_tmp3424 + r_run_k_17);
	assign w_sys_tmp3424 = 32'sh00003e3b;
	assign w_sys_tmp3429 = (w_sys_tmp3430 + r_run_k_17);
	assign w_sys_tmp3430 = 32'sh00003ebc;
	assign w_sys_tmp3435 = (w_sys_tmp3436 + r_run_k_17);
	assign w_sys_tmp3436 = 32'sh00003f3d;
	assign w_sys_tmp3441 = (w_sys_tmp3442 + r_run_k_17);
	assign w_sys_tmp3442 = 32'sh00003fbe;
	assign w_sys_tmp3447 = (w_sys_tmp3448 + r_run_k_17);
	assign w_sys_tmp3448 = 32'sh0000403f;
	assign w_sys_tmp3453 = (w_sys_tmp3454 + r_run_k_17);
	assign w_sys_tmp3454 = 32'sh000040c0;
	assign w_sys_tmp3459 = (w_sys_tmp3460 + r_run_k_17);
	assign w_sys_tmp3460 = 32'sh00004141;
	assign w_sys_tmp3461 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp3462 = 32'sh00000002;
	assign w_sys_tmp3463 = ( !w_sys_tmp3464 );
	assign w_sys_tmp3464 = (w_sys_tmp3465 < r_run_k_17);
	assign w_sys_tmp3465 = 32'sh00000020;
	assign w_sys_tmp3466 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp3467 = 32'sh00000002;
	assign w_sys_tmp3468 = ( !w_sys_tmp3469 );
	assign w_sys_tmp3469 = (w_sys_tmp3470 < r_run_j_18);
	assign w_sys_tmp3470 = 32'sh00000020;
	assign w_sys_tmp3473 = (w_sys_tmp3474 + r_run_k_17);
	assign w_sys_tmp3474 = (r_run_j_18 * w_sys_tmp3475);
	assign w_sys_tmp3475 = 32'sh00000081;
	assign w_sys_tmp3476 = w_sub00_result_dataout;
	assign w_sys_tmp3477 = (w_sys_tmp3478 + r_run_k_17);
	assign w_sys_tmp3478 = (r_run_copy0_j_26 * w_sys_tmp3475);
	assign w_sys_tmp3480 = (r_run_copy0_j_26 + w_sys_intOne);
	assign w_sys_tmp3481 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp3542 = 32'sh00000021;
	assign w_sys_tmp3543 = ( !w_sys_tmp3544 );
	assign w_sys_tmp3544 = (w_sys_tmp3545 < r_run_j_18);
	assign w_sys_tmp3545 = 32'sh00000040;
	assign w_sys_tmp3548 = (w_sys_tmp3549 + r_run_k_17);
	assign w_sys_tmp3549 = (r_run_j_18 * w_sys_tmp3550);
	assign w_sys_tmp3550 = 32'sh00000081;
	assign w_sys_tmp3551 = w_sub01_result_dataout;
	assign w_sys_tmp3552 = (w_sys_tmp3553 + r_run_k_17);
	assign w_sys_tmp3553 = (w_sys_tmp3554 * w_sys_tmp3550);
	assign w_sys_tmp3554 = (r_run_copy0_j_27 - w_sys_tmp3555);
	assign w_sys_tmp3555 = 32'sh0000001f;
	assign w_sys_tmp3557 = (r_run_copy0_j_27 + w_sys_intOne);
	assign w_sys_tmp3558 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp3631 = 32'sh00000041;
	assign w_sys_tmp3632 = ( !w_sys_tmp3633 );
	assign w_sys_tmp3633 = (w_sys_tmp3634 < r_run_j_18);
	assign w_sys_tmp3634 = 32'sh00000060;
	assign w_sys_tmp3637 = (w_sys_tmp3638 + r_run_k_17);
	assign w_sys_tmp3638 = (r_run_j_18 * w_sys_tmp3639);
	assign w_sys_tmp3639 = 32'sh00000081;
	assign w_sys_tmp3640 = w_sub02_result_dataout;
	assign w_sys_tmp3641 = (w_sys_tmp3642 + r_run_k_17);
	assign w_sys_tmp3642 = (w_sys_tmp3643 * w_sys_tmp3639);
	assign w_sys_tmp3643 = (r_run_copy0_j_28 - w_sys_tmp3644);
	assign w_sys_tmp3644 = 32'sh0000003f;
	assign w_sys_tmp3646 = (r_run_copy0_j_28 + w_sys_intOne);
	assign w_sys_tmp3647 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp3720 = 32'sh00000061;
	assign w_sys_tmp3721 = ( !w_sys_tmp3722 );
	assign w_sys_tmp3722 = (w_sys_tmp3723 < r_run_j_18);
	assign w_sys_tmp3723 = 32'sh00000080;
	assign w_sys_tmp3726 = (w_sys_tmp3727 + r_run_k_17);
	assign w_sys_tmp3727 = (r_run_j_18 * w_sys_tmp3728);
	assign w_sys_tmp3728 = 32'sh00000081;
	assign w_sys_tmp3729 = w_sub03_result_dataout;
	assign w_sys_tmp3730 = (w_sys_tmp3731 + r_run_k_17);
	assign w_sys_tmp3731 = (w_sys_tmp3732 * w_sys_tmp3728);
	assign w_sys_tmp3732 = (r_run_copy0_j_29 - w_sys_tmp3733);
	assign w_sys_tmp3733 = 32'sh0000005f;
	assign w_sys_tmp3735 = (r_run_copy0_j_29 + w_sys_intOne);
	assign w_sys_tmp3736 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp3809 = 32'sh00000021;
	assign w_sys_tmp3810 = ( !w_sys_tmp3811 );
	assign w_sys_tmp3811 = (w_sys_tmp3812 < r_run_k_17);
	assign w_sys_tmp3812 = 32'sh00000040;
	assign w_sys_tmp3813 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp3814 = 32'sh00000002;
	assign w_sys_tmp3815 = ( !w_sys_tmp3816 );
	assign w_sys_tmp3816 = (w_sys_tmp3817 < r_run_j_18);
	assign w_sys_tmp3817 = 32'sh00000020;
	assign w_sys_tmp3820 = (w_sys_tmp3821 + r_run_k_17);
	assign w_sys_tmp3821 = (r_run_j_18 * w_sys_tmp3822);
	assign w_sys_tmp3822 = 32'sh00000081;
	assign w_sys_tmp3823 = w_sub04_result_dataout;
	assign w_sys_tmp3824 = (w_sys_tmp3825 + r_run_k_17);
	assign w_sys_tmp3825 = (r_run_copy0_j_30 * w_sys_tmp3822);
	assign w_sys_tmp3827 = (r_run_copy0_j_30 + w_sys_intOne);
	assign w_sys_tmp3828 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp3889 = 32'sh00000021;
	assign w_sys_tmp3890 = ( !w_sys_tmp3891 );
	assign w_sys_tmp3891 = (w_sys_tmp3892 < r_run_j_18);
	assign w_sys_tmp3892 = 32'sh00000040;
	assign w_sys_tmp3895 = (w_sys_tmp3896 + r_run_k_17);
	assign w_sys_tmp3896 = (r_run_j_18 * w_sys_tmp3897);
	assign w_sys_tmp3897 = 32'sh00000081;
	assign w_sys_tmp3898 = w_sub05_result_dataout;
	assign w_sys_tmp3899 = (w_sys_tmp3900 + r_run_k_17);
	assign w_sys_tmp3900 = (w_sys_tmp3901 * w_sys_tmp3897);
	assign w_sys_tmp3901 = (r_run_copy0_j_31 - w_sys_tmp3902);
	assign w_sys_tmp3902 = 32'sh0000001f;
	assign w_sys_tmp3904 = (r_run_copy0_j_31 + w_sys_intOne);
	assign w_sys_tmp3905 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp3978 = 32'sh00000041;
	assign w_sys_tmp3979 = ( !w_sys_tmp3980 );
	assign w_sys_tmp3980 = (w_sys_tmp3981 < r_run_j_18);
	assign w_sys_tmp3981 = 32'sh00000060;
	assign w_sys_tmp3984 = (w_sys_tmp3985 + r_run_k_17);
	assign w_sys_tmp3985 = (r_run_j_18 * w_sys_tmp3986);
	assign w_sys_tmp3986 = 32'sh00000081;
	assign w_sys_tmp3987 = w_sub06_result_dataout;
	assign w_sys_tmp3988 = (w_sys_tmp3989 + r_run_k_17);
	assign w_sys_tmp3989 = (w_sys_tmp3990 * w_sys_tmp3986);
	assign w_sys_tmp3990 = (r_run_copy0_j_32 - w_sys_tmp3991);
	assign w_sys_tmp3991 = 32'sh0000003f;
	assign w_sys_tmp3993 = (r_run_copy0_j_32 + w_sys_intOne);
	assign w_sys_tmp3994 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp4067 = 32'sh00000061;
	assign w_sys_tmp4068 = ( !w_sys_tmp4069 );
	assign w_sys_tmp4069 = (w_sys_tmp4070 < r_run_j_18);
	assign w_sys_tmp4070 = 32'sh00000080;
	assign w_sys_tmp4073 = (w_sys_tmp4074 + r_run_k_17);
	assign w_sys_tmp4074 = (r_run_j_18 * w_sys_tmp4075);
	assign w_sys_tmp4075 = 32'sh00000081;
	assign w_sys_tmp4076 = w_sub07_result_dataout;
	assign w_sys_tmp4077 = (w_sys_tmp4078 + r_run_k_17);
	assign w_sys_tmp4078 = (w_sys_tmp4079 * w_sys_tmp4075);
	assign w_sys_tmp4079 = (r_run_copy0_j_33 - w_sys_tmp4080);
	assign w_sys_tmp4080 = 32'sh0000005f;
	assign w_sys_tmp4082 = (r_run_copy0_j_33 + w_sys_intOne);
	assign w_sys_tmp4083 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp4156 = 32'sh00000041;
	assign w_sys_tmp4157 = ( !w_sys_tmp4158 );
	assign w_sys_tmp4158 = (w_sys_tmp4159 < r_run_k_17);
	assign w_sys_tmp4159 = 32'sh00000060;
	assign w_sys_tmp4160 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp4161 = 32'sh00000002;
	assign w_sys_tmp4162 = ( !w_sys_tmp4163 );
	assign w_sys_tmp4163 = (w_sys_tmp4164 < r_run_j_18);
	assign w_sys_tmp4164 = 32'sh00000020;
	assign w_sys_tmp4167 = (w_sys_tmp4168 + r_run_k_17);
	assign w_sys_tmp4168 = (r_run_j_18 * w_sys_tmp4169);
	assign w_sys_tmp4169 = 32'sh00000081;
	assign w_sys_tmp4170 = w_sub08_result_dataout;
	assign w_sys_tmp4171 = (w_sys_tmp4172 + r_run_k_17);
	assign w_sys_tmp4172 = (r_run_copy0_j_34 * w_sys_tmp4169);
	assign w_sys_tmp4174 = (r_run_copy0_j_34 + w_sys_intOne);
	assign w_sys_tmp4175 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp4236 = 32'sh00000021;
	assign w_sys_tmp4237 = ( !w_sys_tmp4238 );
	assign w_sys_tmp4238 = (w_sys_tmp4239 < r_run_j_18);
	assign w_sys_tmp4239 = 32'sh00000040;
	assign w_sys_tmp4242 = (w_sys_tmp4243 + r_run_k_17);
	assign w_sys_tmp4243 = (r_run_j_18 * w_sys_tmp4244);
	assign w_sys_tmp4244 = 32'sh00000081;
	assign w_sys_tmp4245 = w_sub09_result_dataout;
	assign w_sys_tmp4246 = (w_sys_tmp4247 + r_run_k_17);
	assign w_sys_tmp4247 = (w_sys_tmp4248 * w_sys_tmp4244);
	assign w_sys_tmp4248 = (r_run_copy0_j_35 - w_sys_tmp4249);
	assign w_sys_tmp4249 = 32'sh0000001f;
	assign w_sys_tmp4251 = (r_run_copy0_j_35 + w_sys_intOne);
	assign w_sys_tmp4252 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp4325 = 32'sh00000041;
	assign w_sys_tmp4326 = ( !w_sys_tmp4327 );
	assign w_sys_tmp4327 = (w_sys_tmp4328 < r_run_j_18);
	assign w_sys_tmp4328 = 32'sh00000060;
	assign w_sys_tmp4331 = (w_sys_tmp4332 + r_run_k_17);
	assign w_sys_tmp4332 = (r_run_j_18 * w_sys_tmp4333);
	assign w_sys_tmp4333 = 32'sh00000081;
	assign w_sys_tmp4334 = w_sub10_result_dataout;
	assign w_sys_tmp4335 = (w_sys_tmp4336 + r_run_k_17);
	assign w_sys_tmp4336 = (w_sys_tmp4337 * w_sys_tmp4333);
	assign w_sys_tmp4337 = (r_run_copy0_j_36 - w_sys_tmp4338);
	assign w_sys_tmp4338 = 32'sh0000003f;
	assign w_sys_tmp4340 = (r_run_copy0_j_36 + w_sys_intOne);
	assign w_sys_tmp4341 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp4414 = 32'sh00000061;
	assign w_sys_tmp4415 = ( !w_sys_tmp4416 );
	assign w_sys_tmp4416 = (w_sys_tmp4417 < r_run_j_18);
	assign w_sys_tmp4417 = 32'sh00000080;
	assign w_sys_tmp4420 = (w_sys_tmp4421 + r_run_k_17);
	assign w_sys_tmp4421 = (r_run_j_18 * w_sys_tmp4422);
	assign w_sys_tmp4422 = 32'sh00000081;
	assign w_sys_tmp4423 = w_sub11_result_dataout;
	assign w_sys_tmp4424 = (w_sys_tmp4425 + r_run_k_17);
	assign w_sys_tmp4425 = (w_sys_tmp4426 * w_sys_tmp4422);
	assign w_sys_tmp4426 = (r_run_copy0_j_37 - w_sys_tmp4427);
	assign w_sys_tmp4427 = 32'sh0000005f;
	assign w_sys_tmp4429 = (r_run_copy0_j_37 + w_sys_intOne);
	assign w_sys_tmp4430 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp4503 = 32'sh00000061;
	assign w_sys_tmp4504 = ( !w_sys_tmp4505 );
	assign w_sys_tmp4505 = (w_sys_tmp4506 < r_run_k_17);
	assign w_sys_tmp4506 = 32'sh00000080;
	assign w_sys_tmp4507 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp4508 = 32'sh00000002;
	assign w_sys_tmp4509 = ( !w_sys_tmp4510 );
	assign w_sys_tmp4510 = (w_sys_tmp4511 < r_run_j_18);
	assign w_sys_tmp4511 = 32'sh00000020;
	assign w_sys_tmp4514 = (w_sys_tmp4515 + r_run_k_17);
	assign w_sys_tmp4515 = (r_run_j_18 * w_sys_tmp4516);
	assign w_sys_tmp4516 = 32'sh00000081;
	assign w_sys_tmp4517 = w_sub12_result_dataout;
	assign w_sys_tmp4518 = (w_sys_tmp4519 + r_run_k_17);
	assign w_sys_tmp4519 = (r_run_copy0_j_38 * w_sys_tmp4516);
	assign w_sys_tmp4521 = (r_run_copy0_j_38 + w_sys_intOne);
	assign w_sys_tmp4522 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp4583 = 32'sh00000021;
	assign w_sys_tmp4584 = ( !w_sys_tmp4585 );
	assign w_sys_tmp4585 = (w_sys_tmp4586 < r_run_j_18);
	assign w_sys_tmp4586 = 32'sh00000040;
	assign w_sys_tmp4589 = (w_sys_tmp4590 + r_run_k_17);
	assign w_sys_tmp4590 = (r_run_j_18 * w_sys_tmp4591);
	assign w_sys_tmp4591 = 32'sh00000081;
	assign w_sys_tmp4592 = w_sub13_result_dataout;
	assign w_sys_tmp4593 = (w_sys_tmp4594 + r_run_k_17);
	assign w_sys_tmp4594 = (w_sys_tmp4595 * w_sys_tmp4591);
	assign w_sys_tmp4595 = (r_run_copy0_j_39 - w_sys_tmp4596);
	assign w_sys_tmp4596 = 32'sh0000001f;
	assign w_sys_tmp4598 = (r_run_copy0_j_39 + w_sys_intOne);
	assign w_sys_tmp4599 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp4672 = 32'sh00000041;
	assign w_sys_tmp4673 = ( !w_sys_tmp4674 );
	assign w_sys_tmp4674 = (w_sys_tmp4675 < r_run_j_18);
	assign w_sys_tmp4675 = 32'sh00000060;
	assign w_sys_tmp4678 = (w_sys_tmp4679 + r_run_k_17);
	assign w_sys_tmp4679 = (r_run_j_18 * w_sys_tmp4680);
	assign w_sys_tmp4680 = 32'sh00000081;
	assign w_sys_tmp4681 = w_sub14_result_dataout;
	assign w_sys_tmp4682 = (w_sys_tmp4683 + r_run_k_17);
	assign w_sys_tmp4683 = (w_sys_tmp4684 * w_sys_tmp4680);
	assign w_sys_tmp4684 = (r_run_copy0_j_40 - w_sys_tmp4685);
	assign w_sys_tmp4685 = 32'sh0000003f;
	assign w_sys_tmp4687 = (r_run_copy0_j_40 + w_sys_intOne);
	assign w_sys_tmp4688 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp4761 = 32'sh00000061;
	assign w_sys_tmp4762 = ( !w_sys_tmp4763 );
	assign w_sys_tmp4763 = (w_sys_tmp4764 < r_run_j_18);
	assign w_sys_tmp4764 = 32'sh00000080;
	assign w_sys_tmp4767 = (w_sys_tmp4768 + r_run_k_17);
	assign w_sys_tmp4768 = (r_run_j_18 * w_sys_tmp4769);
	assign w_sys_tmp4769 = 32'sh00000081;
	assign w_sys_tmp4770 = w_sub15_result_dataout;
	assign w_sys_tmp4771 = (w_sys_tmp4772 + r_run_k_17);
	assign w_sys_tmp4772 = (w_sys_tmp4773 * w_sys_tmp4769);
	assign w_sys_tmp4773 = (r_run_copy0_j_41 - w_sys_tmp4774);
	assign w_sys_tmp4774 = 32'sh0000005f;
	assign w_sys_tmp4776 = (r_run_copy0_j_41 + w_sys_intOne);
	assign w_sys_tmp4777 = (r_run_j_18 + w_sys_intOne);


	sub09
		sub09_inst(
			.i_fld_result_1_addr_0 (w_sub09_result_addr),
			.i_fld_result_1_datain_0 (w_sub09_result_datain),
			.o_fld_result_1_dataout_0 (w_sub09_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub09_result_r_w),
			.i_fld_u_0_addr_0 (w_sub09_u_addr),
			.i_fld_u_0_datain_0 (w_sub09_u_datain),
			.o_fld_u_0_dataout_0 (w_sub09_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub09_u_r_w),
			.o_run_busy (w_sub09_run_busy),
			.i_run_req (r_sub09_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub08
		sub08_inst(
			.i_fld_result_1_addr_0 (w_sub08_result_addr),
			.i_fld_result_1_datain_0 (w_sub08_result_datain),
			.o_fld_result_1_dataout_0 (w_sub08_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub08_result_r_w),
			.i_fld_u_0_addr_0 (w_sub08_u_addr),
			.i_fld_u_0_datain_0 (w_sub08_u_datain),
			.o_fld_u_0_dataout_0 (w_sub08_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub08_u_r_w),
			.o_run_busy (w_sub08_run_busy),
			.i_run_req (r_sub08_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub12
		sub12_inst(
			.i_fld_result_1_addr_0 (w_sub12_result_addr),
			.i_fld_result_1_datain_0 (w_sub12_result_datain),
			.o_fld_result_1_dataout_0 (w_sub12_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub12_result_r_w),
			.i_fld_u_0_addr_0 (w_sub12_u_addr),
			.i_fld_u_0_datain_0 (w_sub12_u_datain),
			.o_fld_u_0_dataout_0 (w_sub12_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub12_u_r_w),
			.o_run_busy (w_sub12_run_busy),
			.i_run_req (r_sub12_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub03
		sub03_inst(
			.i_fld_result_1_addr_0 (w_sub03_result_addr),
			.i_fld_result_1_datain_0 (w_sub03_result_datain),
			.o_fld_result_1_dataout_0 (w_sub03_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub03_result_r_w),
			.i_fld_u_0_addr_0 (w_sub03_u_addr),
			.i_fld_u_0_datain_0 (w_sub03_u_datain),
			.o_fld_u_0_dataout_0 (w_sub03_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub03_u_r_w),
			.o_run_busy (w_sub03_run_busy),
			.i_run_req (r_sub03_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub02
		sub02_inst(
			.i_fld_result_1_addr_0 (w_sub02_result_addr),
			.i_fld_result_1_datain_0 (w_sub02_result_datain),
			.o_fld_result_1_dataout_0 (w_sub02_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub02_result_r_w),
			.i_fld_u_0_addr_0 (w_sub02_u_addr),
			.i_fld_u_0_datain_0 (w_sub02_u_datain),
			.o_fld_u_0_dataout_0 (w_sub02_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub02_u_r_w),
			.o_run_busy (w_sub02_run_busy),
			.i_run_req (r_sub02_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub11
		sub11_inst(
			.i_fld_result_1_addr_0 (w_sub11_result_addr),
			.i_fld_result_1_datain_0 (w_sub11_result_datain),
			.o_fld_result_1_dataout_0 (w_sub11_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub11_result_r_w),
			.i_fld_u_0_addr_0 (w_sub11_u_addr),
			.i_fld_u_0_datain_0 (w_sub11_u_datain),
			.o_fld_u_0_dataout_0 (w_sub11_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub11_u_r_w),
			.o_run_busy (w_sub11_run_busy),
			.i_run_req (r_sub11_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub14
		sub14_inst(
			.i_fld_result_1_addr_0 (w_sub14_result_addr),
			.i_fld_result_1_datain_0 (w_sub14_result_datain),
			.o_fld_result_1_dataout_0 (w_sub14_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub14_result_r_w),
			.i_fld_u_0_addr_0 (w_sub14_u_addr),
			.i_fld_u_0_datain_0 (w_sub14_u_datain),
			.o_fld_u_0_dataout_0 (w_sub14_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub14_u_r_w),
			.o_run_busy (w_sub14_run_busy),
			.i_run_req (r_sub14_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub01
		sub01_inst(
			.i_fld_result_1_addr_0 (w_sub01_result_addr),
			.i_fld_result_1_datain_0 (w_sub01_result_datain),
			.o_fld_result_1_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub01_result_r_w),
			.i_fld_u_0_addr_0 (w_sub01_u_addr),
			.i_fld_u_0_datain_0 (w_sub01_u_datain),
			.o_fld_u_0_dataout_0 (w_sub01_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub01_u_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub13
		sub13_inst(
			.i_fld_result_1_addr_0 (w_sub13_result_addr),
			.i_fld_result_1_datain_0 (w_sub13_result_datain),
			.o_fld_result_1_dataout_0 (w_sub13_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub13_result_r_w),
			.i_fld_u_0_addr_0 (w_sub13_u_addr),
			.i_fld_u_0_datain_0 (w_sub13_u_datain),
			.o_fld_u_0_dataout_0 (w_sub13_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub13_u_r_w),
			.o_run_busy (w_sub13_run_busy),
			.i_run_req (r_sub13_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub00
		sub00_inst(
			.i_fld_result_1_addr_0 (w_sub00_result_addr),
			.i_fld_result_1_datain_0 (w_sub00_result_datain),
			.o_fld_result_1_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub00_result_r_w),
			.i_fld_u_0_addr_0 (w_sub00_u_addr),
			.i_fld_u_0_datain_0 (w_sub00_u_datain),
			.o_fld_u_0_dataout_0 (w_sub00_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub00_u_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub07
		sub07_inst(
			.i_fld_result_1_addr_0 (w_sub07_result_addr),
			.i_fld_result_1_datain_0 (w_sub07_result_datain),
			.o_fld_result_1_dataout_0 (w_sub07_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub07_result_r_w),
			.i_fld_u_0_addr_0 (w_sub07_u_addr),
			.i_fld_u_0_datain_0 (w_sub07_u_datain),
			.o_fld_u_0_dataout_0 (w_sub07_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub07_u_r_w),
			.o_run_busy (w_sub07_run_busy),
			.i_run_req (r_sub07_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub06
		sub06_inst(
			.i_fld_result_1_addr_0 (w_sub06_result_addr),
			.i_fld_result_1_datain_0 (w_sub06_result_datain),
			.o_fld_result_1_dataout_0 (w_sub06_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub06_result_r_w),
			.i_fld_u_0_addr_0 (w_sub06_u_addr),
			.i_fld_u_0_datain_0 (w_sub06_u_datain),
			.o_fld_u_0_dataout_0 (w_sub06_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub06_u_r_w),
			.o_run_busy (w_sub06_run_busy),
			.i_run_req (r_sub06_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub15
		sub15_inst(
			.i_fld_result_1_addr_0 (w_sub15_result_addr),
			.i_fld_result_1_datain_0 (w_sub15_result_datain),
			.o_fld_result_1_dataout_0 (w_sub15_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub15_result_r_w),
			.i_fld_u_0_addr_0 (w_sub15_u_addr),
			.i_fld_u_0_datain_0 (w_sub15_u_datain),
			.o_fld_u_0_dataout_0 (w_sub15_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub15_u_r_w),
			.o_run_busy (w_sub15_run_busy),
			.i_run_req (r_sub15_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub05
		sub05_inst(
			.i_fld_result_1_addr_0 (w_sub05_result_addr),
			.i_fld_result_1_datain_0 (w_sub05_result_datain),
			.o_fld_result_1_dataout_0 (w_sub05_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub05_result_r_w),
			.i_fld_u_0_addr_0 (w_sub05_u_addr),
			.i_fld_u_0_datain_0 (w_sub05_u_datain),
			.o_fld_u_0_dataout_0 (w_sub05_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub05_u_r_w),
			.o_run_busy (w_sub05_run_busy),
			.i_run_req (r_sub05_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub04
		sub04_inst(
			.i_fld_result_1_addr_0 (w_sub04_result_addr),
			.i_fld_result_1_datain_0 (w_sub04_result_datain),
			.o_fld_result_1_dataout_0 (w_sub04_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub04_result_r_w),
			.i_fld_u_0_addr_0 (w_sub04_u_addr),
			.i_fld_u_0_datain_0 (w_sub04_u_datain),
			.o_fld_u_0_dataout_0 (w_sub04_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub04_u_r_w),
			.o_run_busy (w_sub04_run_busy),
			.i_run_req (r_sub04_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub10
		sub10_inst(
			.i_fld_result_1_addr_0 (w_sub10_result_addr),
			.i_fld_result_1_datain_0 (w_sub10_result_datain),
			.o_fld_result_1_dataout_0 (w_sub10_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub10_result_r_w),
			.i_fld_u_0_addr_0 (w_sub10_u_addr),
			.i_fld_u_0_datain_0 (w_sub10_u_datain),
			.o_fld_u_0_dataout_0 (w_sub10_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub10_u_r_w),
			.o_run_busy (w_sub10_run_busy),
			.i_run_req (r_sub10_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_u_0(
			.clk (clock),
			.ce_0 (w_fld_u_0_ce_0),
			.addr_0 (w_fld_u_0_addr_0),
			.datain_0 (w_fld_u_0_datain_0),
			.dataout_0 (w_fld_u_0_dataout_0),
			.r_w_0 (w_fld_u_0_r_w_0),
			.ce_1 (w_fld_u_0_ce_1),
			.addr_1 (r_fld_u_0_addr_1),
			.datain_1 (r_fld_u_0_datain_1),
			.dataout_1 (w_fld_u_0_dataout_1),
			.r_w_1 (r_fld_u_0_r_w_1)
		);

	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						8'h9d: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 8'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h0: begin
							r_sys_run_phase <= 8'h2;
						end

						8'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h4;

									end
								end

							endcase
						end

						8'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h5;

									end
								end

							endcase
						end

						8'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3) ? 8'h9 : 8'hf);

									end
								end

							endcase
						end

						8'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h5;

									end
								end

							endcase
						end

						8'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'ha;

									end
								end

							endcase
						end

						8'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6) ? 8'hd : 8'h6);

									end
								end

							endcase
						end

						8'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_run_phase <= 8'ha;

									end
								end

							endcase
						end

						8'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h10;

									end
								end

							endcase
						end

						8'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp51) ? 8'h14 : 8'h9d);

									end
								end

							endcase
						end

						8'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h10;

									end
								end

							endcase
						end

						8'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h15;

									end
								end

							endcase
						end

						8'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp54) ? 8'h18 : 8'h1a);

									end
								end

							endcase
						end

						8'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sys_run_phase <= 8'h15;

									end
								end

							endcase
						end

						8'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h1b;

									end
								end

							endcase
						end

						8'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp211) ? 8'h1e : 8'h20);

									end
								end

							endcase
						end

						8'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h88)) begin
										r_sys_run_phase <= 8'h1b;

									end
								end

							endcase
						end

						8'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h21;

									end
								end

							endcase
						end

						8'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1027) ? 8'h24 : 8'h25);

									end
								end

							endcase
						end

						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h196)) begin
										r_sys_run_phase <= 8'h21;

									end
								end

							endcase
						end

						8'h25: begin

							case(r_sys_run_stage) 
								5'h10: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_phase <= 8'h27;

									end
								end

							endcase
						end

						8'h27: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_phase <= 8'h29;

									end
								end

							endcase
						end

						8'h29: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h2a;

									end
								end

							endcase
						end

						8'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3463) ? 8'h2e : 8'h46);

									end
								end

							endcase
						end

						8'h2b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h2a;

									end
								end

							endcase
						end

						8'h2e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h2f;

									end
								end

							endcase
						end

						8'h2f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3468) ? 8'h32 : 8'h34);

									end
								end

							endcase
						end

						8'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_phase <= 8'h2f;

									end
								end

							endcase
						end

						8'h34: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h35;

									end
								end

							endcase
						end

						8'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3543) ? 8'h38 : 8'h3a);

									end
								end

							endcase
						end

						8'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_phase <= 8'h35;

									end
								end

							endcase
						end

						8'h3a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h3b;

									end
								end

							endcase
						end

						8'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3632) ? 8'h3e : 8'h40);

									end
								end

							endcase
						end

						8'h3e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_phase <= 8'h3b;

									end
								end

							endcase
						end

						8'h40: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h41;

									end
								end

							endcase
						end

						8'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3721) ? 8'h44 : 8'h2b);

									end
								end

							endcase
						end

						8'h44: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_phase <= 8'h41;

									end
								end

							endcase
						end

						8'h46: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h47;

									end
								end

							endcase
						end

						8'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3810) ? 8'h4b : 8'h63);

									end
								end

							endcase
						end

						8'h48: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h47;

									end
								end

							endcase
						end

						8'h4b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h4c;

									end
								end

							endcase
						end

						8'h4c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3815) ? 8'h4f : 8'h51);

									end
								end

							endcase
						end

						8'h4f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_phase <= 8'h4c;

									end
								end

							endcase
						end

						8'h51: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h52;

									end
								end

							endcase
						end

						8'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3890) ? 8'h55 : 8'h57);

									end
								end

							endcase
						end

						8'h55: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_phase <= 8'h52;

									end
								end

							endcase
						end

						8'h57: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h58;

									end
								end

							endcase
						end

						8'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3979) ? 8'h5b : 8'h5d);

									end
								end

							endcase
						end

						8'h5b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_phase <= 8'h58;

									end
								end

							endcase
						end

						8'h5d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h5e;

									end
								end

							endcase
						end

						8'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4068) ? 8'h61 : 8'h48);

									end
								end

							endcase
						end

						8'h61: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_phase <= 8'h5e;

									end
								end

							endcase
						end

						8'h63: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h64;

									end
								end

							endcase
						end

						8'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4157) ? 8'h68 : 8'h80);

									end
								end

							endcase
						end

						8'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h64;

									end
								end

							endcase
						end

						8'h68: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h69;

									end
								end

							endcase
						end

						8'h69: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4162) ? 8'h6c : 8'h6e);

									end
								end

							endcase
						end

						8'h6c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_phase <= 8'h69;

									end
								end

							endcase
						end

						8'h6e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h6f;

									end
								end

							endcase
						end

						8'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4237) ? 8'h72 : 8'h74);

									end
								end

							endcase
						end

						8'h72: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_phase <= 8'h6f;

									end
								end

							endcase
						end

						8'h74: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h75;

									end
								end

							endcase
						end

						8'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4326) ? 8'h78 : 8'h7a);

									end
								end

							endcase
						end

						8'h78: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_phase <= 8'h75;

									end
								end

							endcase
						end

						8'h7a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h7b;

									end
								end

							endcase
						end

						8'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4415) ? 8'h7e : 8'h65);

									end
								end

							endcase
						end

						8'h7e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_phase <= 8'h7b;

									end
								end

							endcase
						end

						8'h80: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h81;

									end
								end

							endcase
						end

						8'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4504) ? 8'h85 : 8'h11);

									end
								end

							endcase
						end

						8'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h81;

									end
								end

							endcase
						end

						8'h85: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h86;

									end
								end

							endcase
						end

						8'h86: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4509) ? 8'h89 : 8'h8b);

									end
								end

							endcase
						end

						8'h89: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_phase <= 8'h86;

									end
								end

							endcase
						end

						8'h8b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h8c;

									end
								end

							endcase
						end

						8'h8c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4584) ? 8'h8f : 8'h91);

									end
								end

							endcase
						end

						8'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_phase <= 8'h8c;

									end
								end

							endcase
						end

						8'h91: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h92;

									end
								end

							endcase
						end

						8'h92: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4673) ? 8'h95 : 8'h97);

									end
								end

							endcase
						end

						8'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_phase <= 8'h92;

									end
								end

							endcase
						end

						8'h97: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 8'h98;

									end
								end

							endcase
						end

						8'h98: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4762) ? 8'h9b : 8'h82);

									end
								end

							endcase
						end

						8'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_phase <= 8'h98;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sys_run_phase <= 8'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 5'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h88)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h196)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h29: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h2b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h2e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h2f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h34: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h3a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h3e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h40: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h44: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h46: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h48: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h4c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h4f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h51: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h55: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h57: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h5b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h5d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h61: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h63: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h68: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h69: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h6c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h6e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h72: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h74: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h78: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h7a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h7e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h80: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h85: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h86: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h89: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h8b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h8c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h91: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h92: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h97: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h98: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						8'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 9'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h5)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						8'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1a)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						8'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h88)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h87)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						8'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h196)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h195)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						8'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub00_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub01_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub02_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub03_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub04_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub05_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub06_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub07_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub08_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub09_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub10_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub11_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub12_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub13_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub14_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub15_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

							endcase
						end

						8'h29: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h2b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h2e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h2f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						8'h34: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						8'h3a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h3e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						8'h40: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h44: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						8'h46: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h48: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h4c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h4f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						8'h51: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h55: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						8'h57: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h5b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						8'h5d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h61: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						8'h63: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h68: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h69: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h6c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						8'h6e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h72: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						8'h74: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h78: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						8'h7a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h7e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						8'h80: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h85: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h86: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h89: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						8'h8b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h8c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						8'h91: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h92: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						8'h97: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h98: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						8'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						8'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						8'h9d: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp10[14:0] );

									end
								end

							endcase
						end

						8'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2) || (r_sys_run_step==9'h6) || (r_sys_run_step==9'ha) || (r_sys_run_step==9'he) || (r_sys_run_step==9'h12) || (r_sys_run_step==9'h16) || (r_sys_run_step==9'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp66[14:0] );

									end
									else
									if((r_sys_run_step==9'h3) || (r_sys_run_step==9'h7) || (r_sys_run_step==9'hb) || (r_sys_run_step==9'hf) || (r_sys_run_step==9'h13) || (r_sys_run_step==9'h17) || (r_sys_run_step==9'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp71[14:0] );

									end
									else
									if((r_sys_run_step==9'h1) || (r_sys_run_step==9'h5) || (r_sys_run_step==9'h9) || (r_sys_run_step==9'hd) || (r_sys_run_step==9'h11) || (r_sys_run_step==9'h15) || (r_sys_run_step==9'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp62[14:0] );

									end
									else
									if((r_sys_run_step==9'h0) || (r_sys_run_step==9'h4) || (r_sys_run_step==9'h8) || (r_sys_run_step==9'hc) || (r_sys_run_step==9'h10) || (r_sys_run_step==9'h14) || (r_sys_run_step==9'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp58[14:0] );

									end
								end

							endcase
						end

						8'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp336[14:0] );

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp435[14:0] );

									end
									else
									if((r_sys_run_step==9'h58)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp747[14:0] );

									end
									else
									if((r_sys_run_step==9'h56)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp735[14:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp360[14:0] );

									end
									else
									if((r_sys_run_step==9'h6a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp855[14:0] );

									end
									else
									if((r_sys_run_step==9'h5d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp777[14:0] );

									end
									else
									if((r_sys_run_step==9'h57)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp741[14:0] );

									end
									else
									if((r_sys_run_step==9'h5a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp759[14:0] );

									end
									else
									if((r_sys_run_step==9'h63) || (r_sys_run_step==9'h65)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp813[14:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp318[14:0] );

									end
									else
									if((r_sys_run_step==9'h48)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp651[14:0] );

									end
									else
									if((r_sys_run_step==9'h86)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1023[14:0] );

									end
									else
									if((r_sys_run_step==9'h83)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1005[14:0] );

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp585[14:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp348[14:0] );

									end
									else
									if((r_sys_run_step==9'h59)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp753[14:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp342[14:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp306[14:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp282[14:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp246[14:0] );

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp579[14:0] );

									end
									else
									if((r_sys_run_step==9'h5f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp789[14:0] );

									end
									else
									if((r_sys_run_step==9'h72)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp903[14:0] );

									end
									else
									if((r_sys_run_step==9'h6b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp861[14:0] );

									end
									else
									if((r_sys_run_step==9'h81)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp993[14:0] );

									end
									else
									if((r_sys_run_step==9'h2a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp471[14:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp390[14:0] );

									end
									else
									if((r_sys_run_step==9'h78)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp939[14:0] );

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp573[14:0] );

									end
									else
									if((r_sys_run_step==9'h3f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp597[14:0] );

									end
									else
									if((r_sys_run_step==9'h7c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp963[14:0] );

									end
									else
									if((r_sys_run_step==9'h7e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp975[14:0] );

									end
									else
									if((r_sys_run_step==9'h6f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp885[14:0] );

									end
									else
									if((r_sys_run_step==9'h68)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp843[14:0] );

									end
									else
									if((r_sys_run_step==9'h76)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp927[14:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp288[14:0] );

									end
									else
									if((r_sys_run_step==9'h36)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp543[14:0] );

									end
									else
									if((r_sys_run_step==9'h29)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp465[14:0] );

									end
									else
									if((r_sys_run_step==9'h33)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp525[14:0] );

									end
									else
									if((r_sys_run_step==9'h4f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp693[14:0] );

									end
									else
									if((r_sys_run_step==9'h20) || (r_sys_run_step==9'h22)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp408[14:0] );

									end
									else
									if((r_sys_run_step==9'h42) || (r_sys_run_step==9'h44)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp615[14:0] );

									end
									else
									if((r_sys_run_step==9'h84)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1011[14:0] );

									end
									else
									if((r_sys_run_step==9'h2d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp489[14:0] );

									end
									else
									if((r_sys_run_step==9'h53)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp717[14:0] );

									end
									else
									if((r_sys_run_step==9'h6d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp873[14:0] );

									end
									else
									if((r_sys_run_step==9'h82)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp999[14:0] );

									end
									else
									if((r_sys_run_step==9'h40)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp603[14:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp300[14:0] );

									end
									else
									if((r_sys_run_step==9'h85)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1017[14:0] );

									end
									else
									if((r_sys_run_step==9'h7f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp981[14:0] );

									end
									else
									if((r_sys_run_step==9'h69)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp849[14:0] );

									end
									else
									if((r_sys_run_step==9'h2e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp495[14:0] );

									end
									else
									if((r_sys_run_step==9'h50)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp699[14:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp396[14:0] );

									end
									else
									if((r_sys_run_step==9'h41) || (r_sys_run_step==9'h43)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp609[14:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp264[14:0] );

									end
									else
									if((r_sys_run_step==9'h5e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp783[14:0] );

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp441[14:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp324[14:0] );

									end
									else
									if((r_sys_run_step==9'h71)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp897[14:0] );

									end
									else
									if((r_sys_run_step==9'h70)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp891[14:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp258[14:0] );

									end
									else
									if((r_sys_run_step==9'h4a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp663[14:0] );

									end
									else
									if((r_sys_run_step==9'h32)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp519[14:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp240[14:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp276[14:0] );

									end
									else
									if((r_sys_run_step==9'h49)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp657[14:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp222[14:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp228[14:0] );

									end
									else
									if((r_sys_run_step==9'h62)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp807[14:0] );

									end
									else
									if((r_sys_run_step==9'h27)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp453[14:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp234[14:0] );

									end
									else
									if((r_sys_run_step==9'h35)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp537[14:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp216[14:0] );

									end
									else
									if((r_sys_run_step==9'h37)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp549[14:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp270[14:0] );

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp675[14:0] );

									end
									else
									if((r_sys_run_step==9'h55)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp729[14:0] );

									end
									else
									if((r_sys_run_step==9'h61)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp801[14:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp384[14:0] );

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp645[14:0] );

									end
									else
									if((r_sys_run_step==9'h74)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp915[14:0] );

									end
									else
									if((r_sys_run_step==9'h64) || (r_sys_run_step==9'h66)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp819[14:0] );

									end
									else
									if((r_sys_run_step==9'h2c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp483[14:0] );

									end
									else
									if((r_sys_run_step==9'h28)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp459[14:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp378[14:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp366[14:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp294[14:0] );

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp687[14:0] );

									end
									else
									if((r_sys_run_step==9'h2b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp477[14:0] );

									end
									else
									if((r_sys_run_step==9'h7a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp951[14:0] );

									end
									else
									if((r_sys_run_step==9'h73)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp909[14:0] );

									end
									else
									if((r_sys_run_step==9'h4d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp681[14:0] );

									end
									else
									if((r_sys_run_step==9'h67)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp837[14:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp330[14:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp354[14:0] );

									end
									else
									if((r_sys_run_step==9'h7d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp969[14:0] );

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp669[14:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp252[14:0] );

									end
									else
									if((r_sys_run_step==9'h60)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp795[14:0] );

									end
									else
									if((r_sys_run_step==9'h79)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp945[14:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp372[14:0] );

									end
									else
									if((r_sys_run_step==9'h1f) || (r_sys_run_step==9'h21)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp402[14:0] );

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp711[14:0] );

									end
									else
									if((r_sys_run_step==9'h30)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp507[14:0] );

									end
									else
									if((r_sys_run_step==9'h31)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp513[14:0] );

									end
									else
									if((r_sys_run_step==9'h6e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp879[14:0] );

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp501[14:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp312[14:0] );

									end
									else
									if((r_sys_run_step==9'h5b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp765[14:0] );

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp723[14:0] );

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp561[14:0] );

									end
									else
									if((r_sys_run_step==9'h77)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp933[14:0] );

									end
									else
									if((r_sys_run_step==9'h51)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp705[14:0] );

									end
									else
									if((r_sys_run_step==9'h75)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp921[14:0] );

									end
									else
									if((r_sys_run_step==9'h6c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp867[14:0] );

									end
									else
									if((r_sys_run_step==9'h7b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp957[14:0] );

									end
									else
									if((r_sys_run_step==9'h38)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp555[14:0] );

									end
									else
									if((r_sys_run_step==9'h34)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp531[14:0] );

									end
									else
									if((r_sys_run_step==9'h3a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp567[14:0] );

									end
									else
									if((r_sys_run_step==9'h45)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp633[14:0] );

									end
									else
									if((r_sys_run_step==9'h3e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp591[14:0] );

									end
									else
									if((r_sys_run_step==9'h80)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp987[14:0] );

									end
									else
									if((r_sys_run_step==9'h26)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp447[14:0] );

									end
									else
									if((r_sys_run_step==9'h46)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp639[14:0] );

									end
									else
									if((r_sys_run_step==9'h23)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp429[14:0] );

									end
									else
									if((r_sys_run_step==9'h5c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp771[14:0] );

									end
								end

							endcase
						end

						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h145)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2985[14:0] );

									end
									else
									if((r_sys_run_step==9'h30)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1323[14:0] );

									end
									else
									if((r_sys_run_step==9'ha5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2022[14:0] );

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1401[14:0] );

									end
									else
									if((r_sys_run_step==9'h8b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1866[14:0] );

									end
									else
									if((r_sys_run_step==9'hd9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2337[14:0] );

									end
									else
									if((r_sys_run_step==9'h161)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3153[14:0] );

									end
									else
									if((r_sys_run_step==9'h116)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2700[14:0] );

									end
									else
									if((r_sys_run_step==9'h117)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2706[14:0] );

									end
									else
									if((r_sys_run_step==9'h92)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1908[14:0] );

									end
									else
									if((r_sys_run_step==9'haa)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2055[14:0] );

									end
									else
									if((r_sys_run_step==9'hf9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2529[14:0] );

									end
									else
									if((r_sys_run_step==9'h144)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2979[14:0] );

									end
									else
									if((r_sys_run_step==9'h72)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1719[14:0] );

									end
									else
									if((r_sys_run_step==9'h2d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1305[14:0] );

									end
									else
									if((r_sys_run_step==9'hc8) || (r_sys_run_step==9'hca)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2235[14:0] );

									end
									else
									if((r_sys_run_step==9'h127)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2802[14:0] );

									end
									else
									if((r_sys_run_step==9'hdd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2361[14:0] );

									end
									else
									if((r_sys_run_step==9'h108)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2619[14:0] );

									end
									else
									if((r_sys_run_step==9'hbb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2157[14:0] );

									end
									else
									if((r_sys_run_step==9'h10d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2649[14:0] );

									end
									else
									if((r_sys_run_step==9'h150) || (r_sys_run_step==9'h152)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3051[14:0] );

									end
									else
									if((r_sys_run_step==9'h28)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1275[14:0] );

									end
									else
									if((r_sys_run_step==9'h7d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1785[14:0] );

									end
									else
									if((r_sys_run_step==9'h75)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1737[14:0] );

									end
									else
									if((r_sys_run_step==9'h15b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3117[14:0] );

									end
									else
									if((r_sys_run_step==9'h14b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3021[14:0] );

									end
									else
									if((r_sys_run_step==9'h110)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2664[14:0] );

									end
									else
									if((r_sys_run_step==9'hdb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2349[14:0] );

									end
									else
									if((r_sys_run_step==9'hd7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2325[14:0] );

									end
									else
									if((r_sys_run_step==9'h7a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1767[14:0] );

									end
									else
									if((r_sys_run_step==9'h113)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2682[14:0] );

									end
									else
									if((r_sys_run_step==9'h180)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3339[14:0] );

									end
									else
									if((r_sys_run_step==9'h15e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3135[14:0] );

									end
									else
									if((r_sys_run_step==9'h11f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2754[14:0] );

									end
									else
									if((r_sys_run_step==9'h36)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1359[14:0] );

									end
									else
									if((r_sys_run_step==9'h120)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2760[14:0] );

									end
									else
									if((r_sys_run_step==9'h7b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1773[14:0] );

									end
									else
									if((r_sys_run_step==9'h11a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2724[14:0] );

									end
									else
									if((r_sys_run_step==9'hac)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2067[14:0] );

									end
									else
									if((r_sys_run_step==9'h138)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2907[14:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1182[14:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1188[14:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1152[14:0] );

									end
									else
									if((r_sys_run_step==9'he7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2421[14:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1080[14:0] );

									end
									else
									if((r_sys_run_step==9'h148)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3003[14:0] );

									end
									else
									if((r_sys_run_step==9'h8f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1890[14:0] );

									end
									else
									if((r_sys_run_step==9'hda)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2343[14:0] );

									end
									else
									if((r_sys_run_step==9'h90)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1896[14:0] );

									end
									else
									if((r_sys_run_step==9'h45)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1449[14:0] );

									end
									else
									if((r_sys_run_step==9'h191)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3441[14:0] );

									end
									else
									if((r_sys_run_step==9'h134)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2883[14:0] );

									end
									else
									if((r_sys_run_step==9'h142)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2967[14:0] );

									end
									else
									if((r_sys_run_step==9'h74)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1731[14:0] );

									end
									else
									if((r_sys_run_step==9'hc7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2229[14:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1128[14:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1086[14:0] );

									end
									else
									if((r_sys_run_step==9'h91)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1902[14:0] );

									end
									else
									if((r_sys_run_step==9'h67)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1653[14:0] );

									end
									else
									if((r_sys_run_step==9'h170)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3243[14:0] );

									end
									else
									if((r_sys_run_step==9'h50)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1515[14:0] );

									end
									else
									if((r_sys_run_step==9'h27)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1269[14:0] );

									end
									else
									if((r_sys_run_step==9'h68)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1659[14:0] );

									end
									else
									if((r_sys_run_step==9'h141)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2961[14:0] );

									end
									else
									if((r_sys_run_step==9'h12a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2820[14:0] );

									end
									else
									if((r_sys_run_step==9'h51)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1521[14:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1056[14:0] );

									end
									else
									if((r_sys_run_step==9'h7e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1791[14:0] );

									end
									else
									if((r_sys_run_step==9'h123)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2778[14:0] );

									end
									else
									if((r_sys_run_step==9'ha6) || (r_sys_run_step==9'ha8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2028[14:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1074[14:0] );

									end
									else
									if((r_sys_run_step==9'he2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2391[14:0] );

									end
									else
									if((r_sys_run_step==9'h64) || (r_sys_run_step==9'h66)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1635[14:0] );

									end
									else
									if((r_sys_run_step==9'ha3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2010[14:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1062[14:0] );

									end
									else
									if((r_sys_run_step==9'h12d) || (r_sys_run_step==9'h12f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2838[14:0] );

									end
									else
									if((r_sys_run_step==9'h11b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2730[14:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1176[14:0] );

									end
									else
									if((r_sys_run_step==9'h155)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3081[14:0] );

									end
									else
									if((r_sys_run_step==9'h98)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1944[14:0] );

									end
									else
									if((r_sys_run_step==9'h6e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1695[14:0] );

									end
									else
									if((r_sys_run_step==9'h158)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3099[14:0] );

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1389[14:0] );

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1257[14:0] );

									end
									else
									if((r_sys_run_step==9'hb8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2139[14:0] );

									end
									else
									if((r_sys_run_step==9'h11e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2748[14:0] );

									end
									else
									if((r_sys_run_step==9'h5d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1593[14:0] );

									end
									else
									if((r_sys_run_step==9'haf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2085[14:0] );

									end
									else
									if((r_sys_run_step==9'hd0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2283[14:0] );

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1395[14:0] );

									end
									else
									if((r_sys_run_step==9'hba)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2151[14:0] );

									end
									else
									if((r_sys_run_step==9'hcc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2259[14:0] );

									end
									else
									if((r_sys_run_step==9'h189)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3393[14:0] );

									end
									else
									if((r_sys_run_step==9'h115)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2694[14:0] );

									end
									else
									if((r_sys_run_step==9'hb1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2097[14:0] );

									end
									else
									if((r_sys_run_step==9'h6c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1683[14:0] );

									end
									else
									if((r_sys_run_step==9'h149)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3009[14:0] );

									end
									else
									if((r_sys_run_step==9'h2b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1293[14:0] );

									end
									else
									if((r_sys_run_step==9'h48)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1467[14:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1200[14:0] );

									end
									else
									if((r_sys_run_step==9'h10c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2643[14:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1170[14:0] );

									end
									else
									if((r_sys_run_step==9'hb3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2109[14:0] );

									end
									else
									if((r_sys_run_step==9'h85)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1833[14:0] );

									end
									else
									if((r_sys_run_step==9'h16a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3207[14:0] );

									end
									else
									if((r_sys_run_step==9'he0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2379[14:0] );

									end
									else
									if((r_sys_run_step==9'h69)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1665[14:0] );

									end
									else
									if((r_sys_run_step==9'h12c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2832[14:0] );

									end
									else
									if((r_sys_run_step==9'h128)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2808[14:0] );

									end
									else
									if((r_sys_run_step==9'h9d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1974[14:0] );

									end
									else
									if((r_sys_run_step==9'he9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2433[14:0] );

									end
									else
									if((r_sys_run_step==9'h193)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3453[14:0] );

									end
									else
									if((r_sys_run_step==9'h122)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2772[14:0] );

									end
									else
									if((r_sys_run_step==9'h124)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2784[14:0] );

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1539[14:0] );

									end
									else
									if((r_sys_run_step==9'h9e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1980[14:0] );

									end
									else
									if((r_sys_run_step==9'h125)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2790[14:0] );

									end
									else
									if((r_sys_run_step==9'h153)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3069[14:0] );

									end
									else
									if((r_sys_run_step==9'hc4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2211[14:0] );

									end
									else
									if((r_sys_run_step==9'hc5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2217[14:0] );

									end
									else
									if((r_sys_run_step==9'h167)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3189[14:0] );

									end
									else
									if((r_sys_run_step==9'h12e) || (r_sys_run_step==9'h130)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2844[14:0] );

									end
									else
									if((r_sys_run_step==9'h106)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2607[14:0] );

									end
									else
									if((r_sys_run_step==9'hf3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2493[14:0] );

									end
									else
									if((r_sys_run_step==9'h140)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2955[14:0] );

									end
									else
									if((r_sys_run_step==9'h8e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1884[14:0] );

									end
									else
									if((r_sys_run_step==9'hc2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2199[14:0] );

									end
									else
									if((r_sys_run_step==9'h121)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2766[14:0] );

									end
									else
									if((r_sys_run_step==9'h111)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2670[14:0] );

									end
									else
									if((r_sys_run_step==9'hce)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2271[14:0] );

									end
									else
									if((r_sys_run_step==9'hd3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2301[14:0] );

									end
									else
									if((r_sys_run_step==9'h162)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3159[14:0] );

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1317[14:0] );

									end
									else
									if((r_sys_run_step==9'h7c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1779[14:0] );

									end
									else
									if((r_sys_run_step==9'h77)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1749[14:0] );

									end
									else
									if((r_sys_run_step==9'h96)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1932[14:0] );

									end
									else
									if((r_sys_run_step==9'h17d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3321[14:0] );

									end
									else
									if((r_sys_run_step==9'h13b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2925[14:0] );

									end
									else
									if((r_sys_run_step==9'h17e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3327[14:0] );

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1503[14:0] );

									end
									else
									if((r_sys_run_step==9'h3f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1413[14:0] );

									end
									else
									if((r_sys_run_step==9'h135)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2889[14:0] );

									end
									else
									if((r_sys_run_step==9'h4f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1509[14:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1158[14:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1212[14:0] );

									end
									else
									if((r_sys_run_step==9'h86)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1839[14:0] );

									end
									else
									if((r_sys_run_step==9'hb6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2127[14:0] );

									end
									else
									if((r_sys_run_step==9'h79)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1761[14:0] );

									end
									else
									if((r_sys_run_step==9'h184)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3363[14:0] );

									end
									else
									if((r_sys_run_step==9'h131)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2865[14:0] );

									end
									else
									if((r_sys_run_step==9'ha0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1992[14:0] );

									end
									else
									if((r_sys_run_step==9'he8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2427[14:0] );

									end
									else
									if((r_sys_run_step==9'h59)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1569[14:0] );

									end
									else
									if((r_sys_run_step==9'h15c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3123[14:0] );

									end
									else
									if((r_sys_run_step==9'h164)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3171[14:0] );

									end
									else
									if((r_sys_run_step==9'h119)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2718[14:0] );

									end
									else
									if((r_sys_run_step==9'h6b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1677[14:0] );

									end
									else
									if((r_sys_run_step==9'h13f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2949[14:0] );

									end
									else
									if((r_sys_run_step==9'h97)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1938[14:0] );

									end
									else
									if((r_sys_run_step==9'ha1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1998[14:0] );

									end
									else
									if((r_sys_run_step==9'ha2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2004[14:0] );

									end
									else
									if((r_sys_run_step==9'h14f) || (r_sys_run_step==9'h151)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3045[14:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1146[14:0] );

									end
									else
									if((r_sys_run_step==9'h15a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3111[14:0] );

									end
									else
									if((r_sys_run_step==9'hef)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2469[14:0] );

									end
									else
									if((r_sys_run_step==9'h3e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1407[14:0] );

									end
									else
									if((r_sys_run_step==9'h9f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1986[14:0] );

									end
									else
									if((r_sys_run_step==9'h137)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2901[14:0] );

									end
									else
									if((r_sys_run_step==9'h16d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3225[14:0] );

									end
									else
									if((r_sys_run_step==9'he1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2385[14:0] );

									end
									else
									if((r_sys_run_step==9'hab)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2061[14:0] );

									end
									else
									if((r_sys_run_step==9'hf5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2505[14:0] );

									end
									else
									if((r_sys_run_step==9'h118)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2712[14:0] );

									end
									else
									if((r_sys_run_step==9'hdf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2373[14:0] );

									end
									else
									if((r_sys_run_step==9'h56)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1551[14:0] );

									end
									else
									if((r_sys_run_step==9'h2a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1287[14:0] );

									end
									else
									if((r_sys_run_step==9'he6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2415[14:0] );

									end
									else
									if((r_sys_run_step==9'h34)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1347[14:0] );

									end
									else
									if((r_sys_run_step==9'h13a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2919[14:0] );

									end
									else
									if((r_sys_run_step==9'h9b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1962[14:0] );

									end
									else
									if((r_sys_run_step==9'hf2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2487[14:0] );

									end
									else
									if((r_sys_run_step==9'hdc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2355[14:0] );

									end
									else
									if((r_sys_run_step==9'h5c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1587[14:0] );

									end
									else
									if((r_sys_run_step==9'he3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2397[14:0] );

									end
									else
									if((r_sys_run_step==9'h103)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2589[14:0] );

									end
									else
									if((r_sys_run_step==9'h1f) || (r_sys_run_step==9'h21)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1218[14:0] );

									end
									else
									if((r_sys_run_step==9'h18d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3417[14:0] );

									end
									else
									if((r_sys_run_step==9'h14d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3033[14:0] );

									end
									else
									if((r_sys_run_step==9'h11c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2736[14:0] );

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1527[14:0] );

									end
									else
									if((r_sys_run_step==9'hbd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2169[14:0] );

									end
									else
									if((r_sys_run_step==9'h6f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1701[14:0] );

									end
									else
									if((r_sys_run_step==9'h31)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1329[14:0] );

									end
									else
									if((r_sys_run_step==9'h10e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2652[14:0] );

									end
									else
									if((r_sys_run_step==9'h160)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3147[14:0] );

									end
									else
									if((r_sys_run_step==9'h95)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1926[14:0] );

									end
									else
									if((r_sys_run_step==9'h26)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1263[14:0] );

									end
									else
									if((r_sys_run_step==9'h70)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1707[14:0] );

									end
									else
									if((r_sys_run_step==9'h146)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2991[14:0] );

									end
									else
									if((r_sys_run_step==9'hd4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2307[14:0] );

									end
									else
									if((r_sys_run_step==9'h35)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1353[14:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1068[14:0] );

									end
									else
									if((r_sys_run_step==9'hd5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2313[14:0] );

									end
									else
									if((r_sys_run_step==9'heb) || (r_sys_run_step==9'hed)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2445[14:0] );

									end
									else
									if((r_sys_run_step==9'h15d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3129[14:0] );

									end
									else
									if((r_sys_run_step==9'hf6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2511[14:0] );

									end
									else
									if((r_sys_run_step==9'h3a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1383[14:0] );

									end
									else
									if((r_sys_run_step==9'h101)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2577[14:0] );

									end
									else
									if((r_sys_run_step==9'hc3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2205[14:0] );

									end
									else
									if((r_sys_run_step==9'h55)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1545[14:0] );

									end
									else
									if((r_sys_run_step==9'h182)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3351[14:0] );

									end
									else
									if((r_sys_run_step==9'h89)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1854[14:0] );

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1377[14:0] );

									end
									else
									if((r_sys_run_step==9'hf4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2499[14:0] );

									end
									else
									if((r_sys_run_step==9'h62)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1623[14:0] );

									end
									else
									if((r_sys_run_step==9'h10b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2637[14:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1032[14:0] );

									end
									else
									if((r_sys_run_step==9'h165)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3177[14:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1116[14:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1194[14:0] );

									end
									else
									if((r_sys_run_step==9'h73)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1725[14:0] );

									end
									else
									if((r_sys_run_step==9'hae)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2079[14:0] );

									end
									else
									if((r_sys_run_step==9'hee)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2463[14:0] );

									end
									else
									if((r_sys_run_step==9'h175)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3273[14:0] );

									end
									else
									if((r_sys_run_step==9'h88)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1848[14:0] );

									end
									else
									if((r_sys_run_step==9'h9c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1968[14:0] );

									end
									else
									if((r_sys_run_step==9'h99)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1950[14:0] );

									end
									else
									if((r_sys_run_step==9'h41) || (r_sys_run_step==9'h43)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1425[14:0] );

									end
									else
									if((r_sys_run_step==9'hfa)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2535[14:0] );

									end
									else
									if((r_sys_run_step==9'h84)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1827[14:0] );

									end
									else
									if((r_sys_run_step==9'h29)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1281[14:0] );

									end
									else
									if((r_sys_run_step==9'hf1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2481[14:0] );

									end
									else
									if((r_sys_run_step==9'h94)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1920[14:0] );

									end
									else
									if((r_sys_run_step==9'h105)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2601[14:0] );

									end
									else
									if((r_sys_run_step==9'he4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2403[14:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1206[14:0] );

									end
									else
									if((r_sys_run_step==9'h17f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3333[14:0] );

									end
									else
									if((r_sys_run_step==9'h159)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3105[14:0] );

									end
									else
									if((r_sys_run_step==9'h6a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1671[14:0] );

									end
									else
									if((r_sys_run_step==9'hd6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2319[14:0] );

									end
									else
									if((r_sys_run_step==9'h76)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1743[14:0] );

									end
									else
									if((r_sys_run_step==9'h7f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1797[14:0] );

									end
									else
									if((r_sys_run_step==9'h42) || (r_sys_run_step==9'h44)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1431[14:0] );

									end
									else
									if((r_sys_run_step==9'h5e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1599[14:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1098[14:0] );

									end
									else
									if((r_sys_run_step==9'h132)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2871[14:0] );

									end
									else
									if((r_sys_run_step==9'h17b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3309[14:0] );

									end
									else
									if((r_sys_run_step==9'h168)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3195[14:0] );

									end
									else
									if((r_sys_run_step==9'h80)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1803[14:0] );

									end
									else
									if((r_sys_run_step==9'hb2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2103[14:0] );

									end
									else
									if((r_sys_run_step==9'hb5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2121[14:0] );

									end
									else
									if((r_sys_run_step==9'hc0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2187[14:0] );

									end
									else
									if((r_sys_run_step==9'h49)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1473[14:0] );

									end
									else
									if((r_sys_run_step==9'h8c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1872[14:0] );

									end
									else
									if((r_sys_run_step==9'h136)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2895[14:0] );

									end
									else
									if((r_sys_run_step==9'h156)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3087[14:0] );

									end
									else
									if((r_sys_run_step==9'h154)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3075[14:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1134[14:0] );

									end
									else
									if((r_sys_run_step==9'h8d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1878[14:0] );

									end
									else
									if((r_sys_run_step==9'h18b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3405[14:0] );

									end
									else
									if((r_sys_run_step==9'h181)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3345[14:0] );

									end
									else
									if((r_sys_run_step==9'h13d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2937[14:0] );

									end
									else
									if((r_sys_run_step==9'h57)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1557[14:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1122[14:0] );

									end
									else
									if((r_sys_run_step==9'h163)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3165[14:0] );

									end
									else
									if((r_sys_run_step==9'h15f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3141[14:0] );

									end
									else
									if((r_sys_run_step==9'hbc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2163[14:0] );

									end
									else
									if((r_sys_run_step==9'hf8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2523[14:0] );

									end
									else
									if((r_sys_run_step==9'h133)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2877[14:0] );

									end
									else
									if((r_sys_run_step==9'h112)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2676[14:0] );

									end
									else
									if((r_sys_run_step==9'h188)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3387[14:0] );

									end
									else
									if((r_sys_run_step==9'hc9) || (r_sys_run_step==9'hcb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2241[14:0] );

									end
									else
									if((r_sys_run_step==9'hf7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2517[14:0] );

									end
									else
									if((r_sys_run_step==9'hd1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2289[14:0] );

									end
									else
									if((r_sys_run_step==9'h58)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1563[14:0] );

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1461[14:0] );

									end
									else
									if((r_sys_run_step==9'h183)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3357[14:0] );

									end
									else
									if((r_sys_run_step==9'h171) || (r_sys_run_step==9'h173)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3249[14:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1044[14:0] );

									end
									else
									if((r_sys_run_step==9'h14a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3015[14:0] );

									end
									else
									if((r_sys_run_step==9'h190)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3435[14:0] );

									end
									else
									if((r_sys_run_step==9'h13e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2943[14:0] );

									end
									else
									if((r_sys_run_step==9'hfd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2553[14:0] );

									end
									else
									if((r_sys_run_step==9'hb9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2145[14:0] );

									end
									else
									if((r_sys_run_step==9'h139)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2913[14:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1164[14:0] );

									end
									else
									if((r_sys_run_step==9'h187)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3381[14:0] );

									end
									else
									if((r_sys_run_step==9'h20) || (r_sys_run_step==9'h22)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1224[14:0] );

									end
									else
									if((r_sys_run_step==9'h185)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3369[14:0] );

									end
									else
									if((r_sys_run_step==9'h169)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3201[14:0] );

									end
									else
									if((r_sys_run_step==9'h16f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3237[14:0] );

									end
									else
									if((r_sys_run_step==9'h172) || (r_sys_run_step==9'h174)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3255[14:0] );

									end
									else
									if((r_sys_run_step==9'h104)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2595[14:0] );

									end
									else
									if((r_sys_run_step==9'hf0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2475[14:0] );

									end
									else
									if((r_sys_run_step==9'hcf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2277[14:0] );

									end
									else
									if((r_sys_run_step==9'hc6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2223[14:0] );

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1485[14:0] );

									end
									else
									if((r_sys_run_step==9'ha7) || (r_sys_run_step==9'ha9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2034[14:0] );

									end
									else
									if((r_sys_run_step==9'h71)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1713[14:0] );

									end
									else
									if((r_sys_run_step==9'h60)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1611[14:0] );

									end
									else
									if((r_sys_run_step==9'hb0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2091[14:0] );

									end
									else
									if((r_sys_run_step==9'h107)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2613[14:0] );

									end
									else
									if((r_sys_run_step==9'hfe)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2559[14:0] );

									end
									else
									if((r_sys_run_step==9'h87)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1842[14:0] );

									end
									else
									if((r_sys_run_step==9'h18a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3399[14:0] );

									end
									else
									if((r_sys_run_step==9'h38)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1371[14:0] );

									end
									else
									if((r_sys_run_step==9'hcd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2265[14:0] );

									end
									else
									if((r_sys_run_step==9'hb7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2133[14:0] );

									end
									else
									if((r_sys_run_step==9'h16c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3219[14:0] );

									end
									else
									if((r_sys_run_step==9'h114)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2688[14:0] );

									end
									else
									if((r_sys_run_step==9'h78)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1755[14:0] );

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1491[14:0] );

									end
									else
									if((r_sys_run_step==9'hff)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2565[14:0] );

									end
									else
									if((r_sys_run_step==9'h2e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1311[14:0] );

									end
									else
									if((r_sys_run_step==9'h16e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3231[14:0] );

									end
									else
									if((r_sys_run_step==9'h5f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1605[14:0] );

									end
									else
									if((r_sys_run_step==9'h93)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1914[14:0] );

									end
									else
									if((r_sys_run_step==9'h11d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2742[14:0] );

									end
									else
									if((r_sys_run_step==9'h176)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3279[14:0] );

									end
									else
									if((r_sys_run_step==9'h14e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3039[14:0] );

									end
									else
									if((r_sys_run_step==9'h177)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3285[14:0] );

									end
									else
									if((r_sys_run_step==9'h109)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2625[14:0] );

									end
									else
									if((r_sys_run_step==9'h126)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2796[14:0] );

									end
									else
									if((r_sys_run_step==9'hbf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2181[14:0] );

									end
									else
									if((r_sys_run_step==9'hea) || (r_sys_run_step==9'hec)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2439[14:0] );

									end
									else
									if((r_sys_run_step==9'h192)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3447[14:0] );

									end
									else
									if((r_sys_run_step==9'h129)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2814[14:0] );

									end
									else
									if((r_sys_run_step==9'he5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2409[14:0] );

									end
									else
									if((r_sys_run_step==9'hde)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2367[14:0] );

									end
									else
									if((r_sys_run_step==9'hd8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2331[14:0] );

									end
									else
									if((r_sys_run_step==9'hbe)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2175[14:0] );

									end
									else
									if((r_sys_run_step==9'h14c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3027[14:0] );

									end
									else
									if((r_sys_run_step==9'h37)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1365[14:0] );

									end
									else
									if((r_sys_run_step==9'h8a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1860[14:0] );

									end
									else
									if((r_sys_run_step==9'hb4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2115[14:0] );

									end
									else
									if((r_sys_run_step==9'ha4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2016[14:0] );

									end
									else
									if((r_sys_run_step==9'hc1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2193[14:0] );

									end
									else
									if((r_sys_run_step==9'h4a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1479[14:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1140[14:0] );

									end
									else
									if((r_sys_run_step==9'hfc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2547[14:0] );

									end
									else
									if((r_sys_run_step==9'hfb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2541[14:0] );

									end
									else
									if((r_sys_run_step==9'h102)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2583[14:0] );

									end
									else
									if((r_sys_run_step==9'h6d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1689[14:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1104[14:0] );

									end
									else
									if((r_sys_run_step==9'h100)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2571[14:0] );

									end
									else
									if((r_sys_run_step==9'h40)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1419[14:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1110[14:0] );

									end
									else
									if((r_sys_run_step==9'h12b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2826[14:0] );

									end
									else
									if((r_sys_run_step==9'h61)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1617[14:0] );

									end
									else
									if((r_sys_run_step==9'h23)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1245[14:0] );

									end
									else
									if((r_sys_run_step==9'h81)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1809[14:0] );

									end
									else
									if((r_sys_run_step==9'h143)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2973[14:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1092[14:0] );

									end
									else
									if((r_sys_run_step==9'h82)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1815[14:0] );

									end
									else
									if((r_sys_run_step==9'h194)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3459[14:0] );

									end
									else
									if((r_sys_run_step==9'h10a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2631[14:0] );

									end
									else
									if((r_sys_run_step==9'h166)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3183[14:0] );

									end
									else
									if((r_sys_run_step==9'h83)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1821[14:0] );

									end
									else
									if((r_sys_run_step==9'h16b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3213[14:0] );

									end
									else
									if((r_sys_run_step==9'h33)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1341[14:0] );

									end
									else
									if((r_sys_run_step==9'h186)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3375[14:0] );

									end
									else
									if((r_sys_run_step==9'had)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2073[14:0] );

									end
									else
									if((r_sys_run_step==9'h46)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1455[14:0] );

									end
									else
									if((r_sys_run_step==9'h9a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1956[14:0] );

									end
									else
									if((r_sys_run_step==9'h53)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1533[14:0] );

									end
									else
									if((r_sys_run_step==9'h18c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3411[14:0] );

									end
									else
									if((r_sys_run_step==9'h17c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3315[14:0] );

									end
									else
									if((r_sys_run_step==9'h2c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1299[14:0] );

									end
									else
									if((r_sys_run_step==9'h13c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2931[14:0] );

									end
									else
									if((r_sys_run_step==9'h63) || (r_sys_run_step==9'h65)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1629[14:0] );

									end
									else
									if((r_sys_run_step==9'h18e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3423[14:0] );

									end
									else
									if((r_sys_run_step==9'h4d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1497[14:0] );

									end
									else
									if((r_sys_run_step==9'h178)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3291[14:0] );

									end
									else
									if((r_sys_run_step==9'h18f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3429[14:0] );

									end
									else
									if((r_sys_run_step==9'h17a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3303[14:0] );

									end
									else
									if((r_sys_run_step==9'hd2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2295[14:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1050[14:0] );

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1251[14:0] );

									end
									else
									if((r_sys_run_step==9'h179)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3297[14:0] );

									end
									else
									if((r_sys_run_step==9'h157)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3093[14:0] );

									end
									else
									if((r_sys_run_step==9'h147)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2997[14:0] );

									end
									else
									if((r_sys_run_step==9'h5b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1581[14:0] );

									end
									else
									if((r_sys_run_step==9'h32)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1335[14:0] );

									end
									else
									if((r_sys_run_step==9'h10f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2658[14:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1038[14:0] );

									end
									else
									if((r_sys_run_step==9'h5a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1575[14:0] );

									end
								end

							endcase
						end

						8'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3473[14:0] );

									end
								end

							endcase
						end

						8'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3548[14:0] );

									end
								end

							endcase
						end

						8'h3e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3637[14:0] );

									end
								end

							endcase
						end

						8'h44: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3726[14:0] );

									end
								end

							endcase
						end

						8'h4f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3820[14:0] );

									end
								end

							endcase
						end

						8'h55: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3895[14:0] );

									end
								end

							endcase
						end

						8'h5b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3984[14:0] );

									end
								end

							endcase
						end

						8'h61: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4073[14:0] );

									end
								end

							endcase
						end

						8'h6c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4167[14:0] );

									end
								end

							endcase
						end

						8'h72: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4242[14:0] );

									end
								end

							endcase
						end

						8'h78: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4331[14:0] );

									end
								end

							endcase
						end

						8'h7e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4420[14:0] );

									end
								end

							endcase
						end

						8'h89: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4514[14:0] );

									end
								end

							endcase
						end

						8'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4589[14:0] );

									end
								end

							endcase
						end

						8'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4678[14:0] );

									end
								end

							endcase
						end

						8'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4767[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp13;

									end
								end

							endcase
						end

						8'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1) || (r_sys_run_step==9'h3) || (r_sys_run_step==9'h5) || (r_sys_run_step==9'h7) || (r_sys_run_step==9'h9) || (r_sys_run_step==9'hb) || (r_sys_run_step==9'hd) || (r_sys_run_step==9'hf) || (r_sys_run_step==9'h11) || (r_sys_run_step==9'h13) || (r_sys_run_step==9'h15) || (r_sys_run_step==9'h17) || (r_sys_run_step==9'h19) || (r_sys_run_step==9'h1b)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp64;

									end
									else
									if((r_sys_run_step==9'h0) || (r_sys_run_step==9'h4) || (r_sys_run_step==9'h8) || (r_sys_run_step==9'hc) || (r_sys_run_step==9'h10) || (r_sys_run_step==9'h14) || (r_sys_run_step==9'h18)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp60;

									end
									else
									if((r_sys_run_step==9'h2) || (r_sys_run_step==9'h6) || (r_sys_run_step==9'ha) || (r_sys_run_step==9'he) || (r_sys_run_step==9'h12) || (r_sys_run_step==9'h16) || (r_sys_run_step==9'h1a)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp69;

									end
								end

							endcase
						end

						8'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp3476;

									end
								end

							endcase
						end

						8'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp3551;

									end
								end

							endcase
						end

						8'h3e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp3640;

									end
								end

							endcase
						end

						8'h44: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp3729;

									end
								end

							endcase
						end

						8'h4f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp3823;

									end
								end

							endcase
						end

						8'h55: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp3898;

									end
								end

							endcase
						end

						8'h5b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp3987;

									end
								end

							endcase
						end

						8'h61: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp4076;

									end
								end

							endcase
						end

						8'h6c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp4170;

									end
								end

							endcase
						end

						8'h72: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp4245;

									end
								end

							endcase
						end

						8'h78: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp4334;

									end
								end

							endcase
						end

						8'h7e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp4423;

									end
								end

							endcase
						end

						8'h89: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp4517;

									end
								end

							endcase
						end

						8'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp4592;

									end
								end

							endcase
						end

						8'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp4681;

									end
								end

							endcase
						end

						8'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp4770;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1b)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h86)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h194)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h3e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h44: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h4f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h55: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h5b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h61: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h6c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h72: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h78: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h7e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h89: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h9d: begin
							r_fld_u_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_17 <= w_sys_intOne;

									end
								end

							endcase
						end

						8'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_17 <= w_sys_tmp5;

									end
								end

							endcase
						end

						8'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_17 <= w_sys_intOne;

									end
								end

							endcase
						end

						8'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h88)) begin
										r_run_k_17 <= w_sys_tmp1025;

									end
								end

							endcase
						end

						8'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_17 <= w_sys_tmp1026;

									end
								end

							endcase
						end

						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h196)) begin
										r_run_k_17 <= w_sys_tmp3461;

									end
								end

							endcase
						end

						8'h29: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_17 <= w_sys_tmp3462;

									end
								end

							endcase
						end

						8'h2b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_17 <= w_sys_tmp3466;

									end
								end

							endcase
						end

						8'h46: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_17 <= w_sys_tmp3809;

									end
								end

							endcase
						end

						8'h48: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_17 <= w_sys_tmp3813;

									end
								end

							endcase
						end

						8'h63: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_17 <= w_sys_tmp4156;

									end
								end

							endcase
						end

						8'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_17 <= w_sys_tmp4160;

									end
								end

							endcase
						end

						8'h80: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_17 <= w_sys_tmp4503;

									end
								end

							endcase
						end

						8'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_17 <= w_sys_tmp4507;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_j_18 <= w_sys_intOne;

									end
								end

							endcase
						end

						8'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_run_j_18 <= w_sys_tmp14;

									end
								end

							endcase
						end

						8'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_j_18 <= w_sys_intOne;

									end
								end

							endcase
						end

						8'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0) || (r_sys_run_step==9'h4) || (r_sys_run_step==9'h8) || (r_sys_run_step==9'hc) || (r_sys_run_step==9'h10) || (r_sys_run_step==9'h14) || (r_sys_run_step==9'h18)) begin
										r_run_j_18 <= w_sys_tmp78;

									end
								end

							endcase
						end

						8'h2e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_j_18 <= w_sys_tmp3467;

									end
								end

							endcase
						end

						8'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_run_j_18 <= w_sys_tmp3481;

									end
								end

							endcase
						end

						8'h34: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_j_18 <= w_sys_tmp3542;

									end
								end

							endcase
						end

						8'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_run_j_18 <= w_sys_tmp3558;

									end
								end

							endcase
						end

						8'h3a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_j_18 <= w_sys_tmp3631;

									end
								end

							endcase
						end

						8'h3e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_run_j_18 <= w_sys_tmp3647;

									end
								end

							endcase
						end

						8'h40: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_j_18 <= w_sys_tmp3720;

									end
								end

							endcase
						end

						8'h44: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_run_j_18 <= w_sys_tmp3736;

									end
								end

							endcase
						end

						8'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_j_18 <= w_sys_tmp3814;

									end
								end

							endcase
						end

						8'h4f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_run_j_18 <= w_sys_tmp3828;

									end
								end

							endcase
						end

						8'h51: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_j_18 <= w_sys_tmp3889;

									end
								end

							endcase
						end

						8'h55: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_run_j_18 <= w_sys_tmp3905;

									end
								end

							endcase
						end

						8'h57: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_j_18 <= w_sys_tmp3978;

									end
								end

							endcase
						end

						8'h5b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_run_j_18 <= w_sys_tmp3994;

									end
								end

							endcase
						end

						8'h5d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_j_18 <= w_sys_tmp4067;

									end
								end

							endcase
						end

						8'h61: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_run_j_18 <= w_sys_tmp4083;

									end
								end

							endcase
						end

						8'h68: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_j_18 <= w_sys_tmp4161;

									end
								end

							endcase
						end

						8'h6c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_run_j_18 <= w_sys_tmp4175;

									end
								end

							endcase
						end

						8'h6e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_j_18 <= w_sys_tmp4236;

									end
								end

							endcase
						end

						8'h72: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_run_j_18 <= w_sys_tmp4252;

									end
								end

							endcase
						end

						8'h74: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_j_18 <= w_sys_tmp4325;

									end
								end

							endcase
						end

						8'h78: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_run_j_18 <= w_sys_tmp4341;

									end
								end

							endcase
						end

						8'h7a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_j_18 <= w_sys_tmp4414;

									end
								end

							endcase
						end

						8'h7e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_run_j_18 <= w_sys_tmp4430;

									end
								end

							endcase
						end

						8'h85: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_j_18 <= w_sys_tmp4508;

									end
								end

							endcase
						end

						8'h89: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_run_j_18 <= w_sys_tmp4522;

									end
								end

							endcase
						end

						8'h8b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_j_18 <= w_sys_tmp4583;

									end
								end

							endcase
						end

						8'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_run_j_18 <= w_sys_tmp4599;

									end
								end

							endcase
						end

						8'h91: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_j_18 <= w_sys_tmp4672;

									end
								end

							endcase
						end

						8'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_run_j_18 <= w_sys_tmp4688;

									end
								end

							endcase
						end

						8'h97: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_j_18 <= w_sys_tmp4761;

									end
								end

							endcase
						end

						8'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_run_j_18 <= w_sys_tmp4777;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_n_19 <= w_sys_intOne;

									end
								end

							endcase
						end

						8'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_n_19 <= w_sys_tmp53;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_mx_20 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_my_21 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_nlast_22 <= w_sys_intOne;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy0_j_23 <= r_run_j_18;

									end
								end

							endcase
						end

						8'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3) || (r_sys_run_step==9'h7) || (r_sys_run_step==9'hb) || (r_sys_run_step==9'hf) || (r_sys_run_step==9'h13) || (r_sys_run_step==9'h17) || (r_sys_run_step==9'h1b)) begin
										r_run_copy0_j_23 <= w_sys_tmp75;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy1_j_24 <= r_run_j_18;

									end
								end

							endcase
						end

						8'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2) || (r_sys_run_step==9'h6) || (r_sys_run_step==9'ha) || (r_sys_run_step==9'he) || (r_sys_run_step==9'h12) || (r_sys_run_step==9'h16) || (r_sys_run_step==9'h1a)) begin
										r_run_copy1_j_24 <= w_sys_tmp76;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy2_j_25 <= r_run_j_18;

									end
								end

							endcase
						end

						8'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1) || (r_sys_run_step==9'h5) || (r_sys_run_step==9'h9) || (r_sys_run_step==9'hd) || (r_sys_run_step==9'h11) || (r_sys_run_step==9'h15) || (r_sys_run_step==9'h19)) begin
										r_run_copy2_j_25 <= w_sys_tmp77;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h2e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy0_j_26 <= r_run_j_18;

									end
								end

							endcase
						end

						8'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_run_copy0_j_26 <= w_sys_tmp3480;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h34: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy0_j_27 <= r_run_j_18;

									end
								end

							endcase
						end

						8'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_run_copy0_j_27 <= w_sys_tmp3557;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h3a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy0_j_28 <= r_run_j_18;

									end
								end

							endcase
						end

						8'h3e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_run_copy0_j_28 <= w_sys_tmp3646;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h40: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy0_j_29 <= r_run_j_18;

									end
								end

							endcase
						end

						8'h44: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_run_copy0_j_29 <= w_sys_tmp3735;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h4b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy0_j_30 <= r_run_j_18;

									end
								end

							endcase
						end

						8'h4f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_run_copy0_j_30 <= w_sys_tmp3827;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h51: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy0_j_31 <= r_run_j_18;

									end
								end

							endcase
						end

						8'h55: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_run_copy0_j_31 <= w_sys_tmp3904;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h57: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy0_j_32 <= r_run_j_18;

									end
								end

							endcase
						end

						8'h5b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_run_copy0_j_32 <= w_sys_tmp3993;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h5d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy0_j_33 <= r_run_j_18;

									end
								end

							endcase
						end

						8'h61: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_run_copy0_j_33 <= w_sys_tmp4082;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h68: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy0_j_34 <= r_run_j_18;

									end
								end

							endcase
						end

						8'h6c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_run_copy0_j_34 <= w_sys_tmp4174;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h6e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy0_j_35 <= r_run_j_18;

									end
								end

							endcase
						end

						8'h72: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_run_copy0_j_35 <= w_sys_tmp4251;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h74: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy0_j_36 <= r_run_j_18;

									end
								end

							endcase
						end

						8'h78: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_run_copy0_j_36 <= w_sys_tmp4340;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h7a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy0_j_37 <= r_run_j_18;

									end
								end

							endcase
						end

						8'h7e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_run_copy0_j_37 <= w_sys_tmp4429;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h85: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy0_j_38 <= r_run_j_18;

									end
								end

							endcase
						end

						8'h89: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_run_copy0_j_38 <= w_sys_tmp4521;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h8b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy0_j_39 <= r_run_j_18;

									end
								end

							endcase
						end

						8'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_run_copy0_j_39 <= w_sys_tmp4598;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h91: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy0_j_40 <= r_run_j_18;

									end
								end

							endcase
						end

						8'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_run_copy0_j_40 <= w_sys_tmp4687;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h97: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy0_j_41 <= r_run_j_18;

									end
								end

							endcase
						end

						8'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_run_copy0_j_41 <= w_sys_tmp4776;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'h7: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub09_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub09_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc7)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2016[12:0] );

									end
									else
									if((r_sys_run_step==9'hc8)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2022[12:0] );

									end
									else
									if((r_sys_run_step==9'hb7)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp1920[12:0] );

									end
									else
									if((r_sys_run_step==9'hbb)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp1944[12:0] );

									end
									else
									if((r_sys_run_step==9'hae)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp1866[12:0] );

									end
									else
									if((r_sys_run_step==9'hb1)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp1884[12:0] );

									end
									else
									if((r_sys_run_step==9'hbe)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp1962[12:0] );

									end
									else
									if((r_sys_run_step==9'hb5)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp1908[12:0] );

									end
									else
									if((r_sys_run_step==9'hcb)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2055[12:0] );

									end
									else
									if((r_sys_run_step==9'hb2)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp1890[12:0] );

									end
									else
									if((r_sys_run_step==9'hb9)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp1932[12:0] );

									end
									else
									if((r_sys_run_step==9'hb3)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp1896[12:0] );

									end
									else
									if((r_sys_run_step==9'hca)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2034[12:0] );

									end
									else
									if((r_sys_run_step==9'hb8)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp1926[12:0] );

									end
									else
									if((r_sys_run_step==9'haa)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp1842[12:0] );

									end
									else
									if((r_sys_run_step==9'hbd)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp1956[12:0] );

									end
									else
									if((r_sys_run_step==9'haf)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp1872[12:0] );

									end
									else
									if((r_sys_run_step==9'hc3)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp1992[12:0] );

									end
									else
									if((r_sys_run_step==9'hb0)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp1878[12:0] );

									end
									else
									if((r_sys_run_step==9'hb4)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp1902[12:0] );

									end
									else
									if((r_sys_run_step==9'hb6)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp1914[12:0] );

									end
									else
									if((r_sys_run_step==9'hba)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp1938[12:0] );

									end
									else
									if((r_sys_run_step==9'hc0)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp1974[12:0] );

									end
									else
									if((r_sys_run_step==9'hac)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp1854[12:0] );

									end
									else
									if((r_sys_run_step==9'hc5)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2004[12:0] );

									end
									else
									if((r_sys_run_step==9'hc4)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp1998[12:0] );

									end
									else
									if((r_sys_run_step==9'hc1)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp1980[12:0] );

									end
									else
									if((r_sys_run_step==9'hc2)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp1986[12:0] );

									end
									else
									if((r_sys_run_step==9'hc9)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2028[12:0] );

									end
									else
									if((r_sys_run_step==9'hab)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp1848[12:0] );

									end
									else
									if((r_sys_run_step==9'hbf)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp1968[12:0] );

									end
									else
									if((r_sys_run_step==9'hbc)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp1950[12:0] );

									end
									else
									if((r_sys_run_step==9'hc6)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2010[12:0] );

									end
									else
									if((r_sys_run_step==9'had)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp1860[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'haa<=r_sys_run_step && r_sys_run_step<=9'hcb)) begin
										r_sub09_u_datain <= w_sys_tmp1034;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'haa<=r_sys_run_step && r_sys_run_step<=9'hcb)) begin
										r_sub09_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub09_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h72: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4246[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h72: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub09_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub08_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub08_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha6)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp2016[12:0] );

									end
									else
									if((r_sys_run_step==9'ha7)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp2022[12:0] );

									end
									else
									if((r_sys_run_step==9'h96)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1920[12:0] );

									end
									else
									if((r_sys_run_step==9'h9a)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1944[12:0] );

									end
									else
									if((r_sys_run_step==9'h8d)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1866[12:0] );

									end
									else
									if((r_sys_run_step==9'h90)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1884[12:0] );

									end
									else
									if((r_sys_run_step==9'h9d)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1962[12:0] );

									end
									else
									if((r_sys_run_step==9'h94)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1908[12:0] );

									end
									else
									if((r_sys_run_step==9'h91)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1890[12:0] );

									end
									else
									if((r_sys_run_step==9'h98)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1932[12:0] );

									end
									else
									if((r_sys_run_step==9'h92)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1896[12:0] );

									end
									else
									if((r_sys_run_step==9'ha9)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp2034[12:0] );

									end
									else
									if((r_sys_run_step==9'h97)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1926[12:0] );

									end
									else
									if((r_sys_run_step==9'h89)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1842[12:0] );

									end
									else
									if((r_sys_run_step==9'h9c)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1956[12:0] );

									end
									else
									if((r_sys_run_step==9'h8e)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1872[12:0] );

									end
									else
									if((r_sys_run_step==9'ha2)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1992[12:0] );

									end
									else
									if((r_sys_run_step==9'h8f)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1878[12:0] );

									end
									else
									if((r_sys_run_step==9'h93)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1902[12:0] );

									end
									else
									if((r_sys_run_step==9'h95)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1914[12:0] );

									end
									else
									if((r_sys_run_step==9'h99)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1938[12:0] );

									end
									else
									if((r_sys_run_step==9'h9f)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1974[12:0] );

									end
									else
									if((r_sys_run_step==9'h8b)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1854[12:0] );

									end
									else
									if((r_sys_run_step==9'ha4)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp2004[12:0] );

									end
									else
									if((r_sys_run_step==9'ha3)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1998[12:0] );

									end
									else
									if((r_sys_run_step==9'ha0)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1980[12:0] );

									end
									else
									if((r_sys_run_step==9'ha1)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1986[12:0] );

									end
									else
									if((r_sys_run_step==9'ha8)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp2028[12:0] );

									end
									else
									if((r_sys_run_step==9'h8a)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1848[12:0] );

									end
									else
									if((r_sys_run_step==9'h9e)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1968[12:0] );

									end
									else
									if((r_sys_run_step==9'h9b)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1950[12:0] );

									end
									else
									if((r_sys_run_step==9'ha5)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp2010[12:0] );

									end
									else
									if((r_sys_run_step==9'h8c)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1860[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h89<=r_sys_run_step && r_sys_run_step<=9'ha9)) begin
										r_sub08_u_datain <= w_sys_tmp1034;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h89<=r_sys_run_step && r_sys_run_step<=9'ha9)) begin
										r_sub08_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub08_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h6c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4171[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h6c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub08_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'h10: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub12_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub12_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12f)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2838[12:0] );

									end
									else
									if((r_sys_run_step==9'h11a)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2712[12:0] );

									end
									else
									if((r_sys_run_step==9'h11d)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2730[12:0] );

									end
									else
									if((r_sys_run_step==9'h118)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2700[12:0] );

									end
									else
									if((r_sys_run_step==9'h12d)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2826[12:0] );

									end
									else
									if((r_sys_run_step==9'h113)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2670[12:0] );

									end
									else
									if((r_sys_run_step==9'h120)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2748[12:0] );

									end
									else
									if((r_sys_run_step==9'h123)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2766[12:0] );

									end
									else
									if((r_sys_run_step==9'h119)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2706[12:0] );

									end
									else
									if((r_sys_run_step==9'h11e)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2736[12:0] );

									end
									else
									if((r_sys_run_step==9'h117)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2694[12:0] );

									end
									else
									if((r_sys_run_step==9'h110)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2652[12:0] );

									end
									else
									if((r_sys_run_step==9'h129)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2802[12:0] );

									end
									else
									if((r_sys_run_step==9'h116)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2688[12:0] );

									end
									else
									if((r_sys_run_step==9'h11b)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2718[12:0] );

									end
									else
									if((r_sys_run_step==9'h112)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2664[12:0] );

									end
									else
									if((r_sys_run_step==9'h12e)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2832[12:0] );

									end
									else
									if((r_sys_run_step==9'h12a)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2808[12:0] );

									end
									else
									if((r_sys_run_step==9'h11f)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2742[12:0] );

									end
									else
									if((r_sys_run_step==9'h115)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2682[12:0] );

									end
									else
									if((r_sys_run_step==9'h121)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2754[12:0] );

									end
									else
									if((r_sys_run_step==9'h124)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2772[12:0] );

									end
									else
									if((r_sys_run_step==9'h12c)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2820[12:0] );

									end
									else
									if((r_sys_run_step==9'h128)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2796[12:0] );

									end
									else
									if((r_sys_run_step==9'h126)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2784[12:0] );

									end
									else
									if((r_sys_run_step==9'h122)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2760[12:0] );

									end
									else
									if((r_sys_run_step==9'h127)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2790[12:0] );

									end
									else
									if((r_sys_run_step==9'h114)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2676[12:0] );

									end
									else
									if((r_sys_run_step==9'h125)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2778[12:0] );

									end
									else
									if((r_sys_run_step==9'h12b)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2814[12:0] );

									end
									else
									if((r_sys_run_step==9'h11c)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2724[12:0] );

									end
									else
									if((r_sys_run_step==9'h111)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2658[12:0] );

									end
									else
									if((r_sys_run_step==9'h130)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2844[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h110<=r_sys_run_step && r_sys_run_step<=9'h130)) begin
										r_sub12_u_datain <= w_sys_tmp1034;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h110<=r_sys_run_step && r_sys_run_step<=9'h130)) begin
										r_sub12_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub12_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h89: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp4518[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h89: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub12_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'h3: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7b)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp336[12:0] );

									end
									else
									if((r_sys_run_step==9'h7a)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp330[12:0] );

									end
									else
									if((r_sys_run_step==9'h7e)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp354[12:0] );

									end
									else
									if((r_sys_run_step==9'h7f)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp360[12:0] );

									end
									else
									if((r_sys_run_step==9'h71)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp276[12:0] );

									end
									else
									if((r_sys_run_step==9'h73)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp288[12:0] );

									end
									else
									if((r_sys_run_step==9'h6d)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp252[12:0] );

									end
									else
									if((r_sys_run_step==9'h68)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp222[12:0] );

									end
									else
									if((r_sys_run_step==9'h78)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp318[12:0] );

									end
									else
									if((r_sys_run_step==9'h81)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp372[12:0] );

									end
									else
									if((r_sys_run_step==9'h86)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp402[12:0] );

									end
									else
									if((r_sys_run_step==9'h69)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp228[12:0] );

									end
									else
									if((r_sys_run_step==9'h7d)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp348[12:0] );

									end
									else
									if((r_sys_run_step==9'h87)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp408[12:0] );

									end
									else
									if((r_sys_run_step==9'h7c)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp342[12:0] );

									end
									else
									if((r_sys_run_step==9'h6a)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp234[12:0] );

									end
									else
									if((r_sys_run_step==9'h76)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp306[12:0] );

									end
									else
									if((r_sys_run_step==9'h72)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp282[12:0] );

									end
									else
									if((r_sys_run_step==9'h67)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp216[12:0] );

									end
									else
									if((r_sys_run_step==9'h70)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp270[12:0] );

									end
									else
									if((r_sys_run_step==9'h75)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp300[12:0] );

									end
									else
									if((r_sys_run_step==9'h77)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp312[12:0] );

									end
									else
									if((r_sys_run_step==9'h6c)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp246[12:0] );

									end
									else
									if((r_sys_run_step==9'h85)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp396[12:0] );

									end
									else
									if((r_sys_run_step==9'h83)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp384[12:0] );

									end
									else
									if((r_sys_run_step==9'h6f)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp264[12:0] );

									end
									else
									if((r_sys_run_step==9'h84)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp390[12:0] );

									end
									else
									if((r_sys_run_step==9'h79)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp324[12:0] );

									end
									else
									if((r_sys_run_step==9'h82)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp378[12:0] );

									end
									else
									if((r_sys_run_step==9'h80)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp366[12:0] );

									end
									else
									if((r_sys_run_step==9'h6e)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp258[12:0] );

									end
									else
									if((r_sys_run_step==9'h74)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp294[12:0] );

									end
									else
									if((r_sys_run_step==9'h6b)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp240[12:0] );

									end
									else
									if((r_sys_run_step==9'h88)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp429[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h67<=r_sys_run_step && r_sys_run_step<=9'h88)) begin
										r_sub03_u_datain <= w_sys_tmp218;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h67<=r_sys_run_step && r_sys_run_step<=9'h88)) begin
										r_sub03_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub03_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h44: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp3730[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h44: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub03_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'h2: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h59)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp336[12:0] );

									end
									else
									if((r_sys_run_step==9'h58)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp330[12:0] );

									end
									else
									if((r_sys_run_step==9'h5c)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp354[12:0] );

									end
									else
									if((r_sys_run_step==9'h5d)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp360[12:0] );

									end
									else
									if((r_sys_run_step==9'h4f)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp276[12:0] );

									end
									else
									if((r_sys_run_step==9'h51)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp288[12:0] );

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp252[12:0] );

									end
									else
									if((r_sys_run_step==9'h46)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp222[12:0] );

									end
									else
									if((r_sys_run_step==9'h56)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp318[12:0] );

									end
									else
									if((r_sys_run_step==9'h5f)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp372[12:0] );

									end
									else
									if((r_sys_run_step==9'h64)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp402[12:0] );

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp228[12:0] );

									end
									else
									if((r_sys_run_step==9'h5b)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp348[12:0] );

									end
									else
									if((r_sys_run_step==9'h65)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp408[12:0] );

									end
									else
									if((r_sys_run_step==9'h5a)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp342[12:0] );

									end
									else
									if((r_sys_run_step==9'h48)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp234[12:0] );

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp306[12:0] );

									end
									else
									if((r_sys_run_step==9'h50)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp282[12:0] );

									end
									else
									if((r_sys_run_step==9'h45)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp216[12:0] );

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp270[12:0] );

									end
									else
									if((r_sys_run_step==9'h53)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp300[12:0] );

									end
									else
									if((r_sys_run_step==9'h55)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp312[12:0] );

									end
									else
									if((r_sys_run_step==9'h4a)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp246[12:0] );

									end
									else
									if((r_sys_run_step==9'h63)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp396[12:0] );

									end
									else
									if((r_sys_run_step==9'h61)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp384[12:0] );

									end
									else
									if((r_sys_run_step==9'h4d)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp264[12:0] );

									end
									else
									if((r_sys_run_step==9'h62)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp390[12:0] );

									end
									else
									if((r_sys_run_step==9'h57)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp324[12:0] );

									end
									else
									if((r_sys_run_step==9'h60)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp378[12:0] );

									end
									else
									if((r_sys_run_step==9'h5e)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp366[12:0] );

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp258[12:0] );

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp294[12:0] );

									end
									else
									if((r_sys_run_step==9'h49)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp240[12:0] );

									end
									else
									if((r_sys_run_step==9'h66)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp429[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h45<=r_sys_run_step && r_sys_run_step<=9'h66)) begin
										r_sub02_u_datain <= w_sys_tmp218;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h45<=r_sys_run_step && r_sys_run_step<=9'h66)) begin
										r_sub02_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub02_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h3e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3641[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h3e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub02_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'h9: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub11_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub11_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10b)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2016[12:0] );

									end
									else
									if((r_sys_run_step==9'h10c)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2022[12:0] );

									end
									else
									if((r_sys_run_step==9'hfb)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1920[12:0] );

									end
									else
									if((r_sys_run_step==9'hff)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1944[12:0] );

									end
									else
									if((r_sys_run_step==9'hf2)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1866[12:0] );

									end
									else
									if((r_sys_run_step==9'hf5)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1884[12:0] );

									end
									else
									if((r_sys_run_step==9'h102)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1962[12:0] );

									end
									else
									if((r_sys_run_step==9'hf9)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1908[12:0] );

									end
									else
									if((r_sys_run_step==9'h10f)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2055[12:0] );

									end
									else
									if((r_sys_run_step==9'hf6)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1890[12:0] );

									end
									else
									if((r_sys_run_step==9'hfd)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1932[12:0] );

									end
									else
									if((r_sys_run_step==9'hf7)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1896[12:0] );

									end
									else
									if((r_sys_run_step==9'h10e)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2034[12:0] );

									end
									else
									if((r_sys_run_step==9'hfc)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1926[12:0] );

									end
									else
									if((r_sys_run_step==9'hee)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1842[12:0] );

									end
									else
									if((r_sys_run_step==9'h101)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1956[12:0] );

									end
									else
									if((r_sys_run_step==9'hf3)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1872[12:0] );

									end
									else
									if((r_sys_run_step==9'h107)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1992[12:0] );

									end
									else
									if((r_sys_run_step==9'hf4)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1878[12:0] );

									end
									else
									if((r_sys_run_step==9'hf8)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1902[12:0] );

									end
									else
									if((r_sys_run_step==9'hfa)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1914[12:0] );

									end
									else
									if((r_sys_run_step==9'hfe)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1938[12:0] );

									end
									else
									if((r_sys_run_step==9'h104)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1974[12:0] );

									end
									else
									if((r_sys_run_step==9'hf0)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1854[12:0] );

									end
									else
									if((r_sys_run_step==9'h109)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2004[12:0] );

									end
									else
									if((r_sys_run_step==9'h108)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1998[12:0] );

									end
									else
									if((r_sys_run_step==9'h105)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1980[12:0] );

									end
									else
									if((r_sys_run_step==9'h106)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1986[12:0] );

									end
									else
									if((r_sys_run_step==9'h10d)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2028[12:0] );

									end
									else
									if((r_sys_run_step==9'hef)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1848[12:0] );

									end
									else
									if((r_sys_run_step==9'h103)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1968[12:0] );

									end
									else
									if((r_sys_run_step==9'h100)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1950[12:0] );

									end
									else
									if((r_sys_run_step==9'h10a)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2010[12:0] );

									end
									else
									if((r_sys_run_step==9'hf1)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1860[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'hee<=r_sys_run_step && r_sys_run_step<=9'h10f)) begin
										r_sub11_u_datain <= w_sys_tmp1034;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'hee<=r_sys_run_step && r_sys_run_step<=9'h10f)) begin
										r_sub11_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub11_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h7e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp4424[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h7e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub11_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'hb: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub14_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub14_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h172)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2838[12:0] );

									end
									else
									if((r_sys_run_step==9'h15d)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2712[12:0] );

									end
									else
									if((r_sys_run_step==9'h160)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2730[12:0] );

									end
									else
									if((r_sys_run_step==9'h15b)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2700[12:0] );

									end
									else
									if((r_sys_run_step==9'h170)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2826[12:0] );

									end
									else
									if((r_sys_run_step==9'h156)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2670[12:0] );

									end
									else
									if((r_sys_run_step==9'h163)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2748[12:0] );

									end
									else
									if((r_sys_run_step==9'h166)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2766[12:0] );

									end
									else
									if((r_sys_run_step==9'h15c)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2706[12:0] );

									end
									else
									if((r_sys_run_step==9'h161)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2736[12:0] );

									end
									else
									if((r_sys_run_step==9'h15a)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2694[12:0] );

									end
									else
									if((r_sys_run_step==9'h153)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2652[12:0] );

									end
									else
									if((r_sys_run_step==9'h16c)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2802[12:0] );

									end
									else
									if((r_sys_run_step==9'h174)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2865[12:0] );

									end
									else
									if((r_sys_run_step==9'h159)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2688[12:0] );

									end
									else
									if((r_sys_run_step==9'h15e)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2718[12:0] );

									end
									else
									if((r_sys_run_step==9'h155)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2664[12:0] );

									end
									else
									if((r_sys_run_step==9'h171)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2832[12:0] );

									end
									else
									if((r_sys_run_step==9'h16d)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2808[12:0] );

									end
									else
									if((r_sys_run_step==9'h162)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2742[12:0] );

									end
									else
									if((r_sys_run_step==9'h158)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2682[12:0] );

									end
									else
									if((r_sys_run_step==9'h164)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2754[12:0] );

									end
									else
									if((r_sys_run_step==9'h167)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2772[12:0] );

									end
									else
									if((r_sys_run_step==9'h16f)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2820[12:0] );

									end
									else
									if((r_sys_run_step==9'h16b)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2796[12:0] );

									end
									else
									if((r_sys_run_step==9'h169)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2784[12:0] );

									end
									else
									if((r_sys_run_step==9'h165)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2760[12:0] );

									end
									else
									if((r_sys_run_step==9'h16a)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2790[12:0] );

									end
									else
									if((r_sys_run_step==9'h157)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2676[12:0] );

									end
									else
									if((r_sys_run_step==9'h168)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2778[12:0] );

									end
									else
									if((r_sys_run_step==9'h16e)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2814[12:0] );

									end
									else
									if((r_sys_run_step==9'h15f)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2724[12:0] );

									end
									else
									if((r_sys_run_step==9'h154)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2658[12:0] );

									end
									else
									if((r_sys_run_step==9'h173)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp2844[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h153<=r_sys_run_step && r_sys_run_step<=9'h174)) begin
										r_sub14_u_datain <= w_sys_tmp1034;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h153<=r_sys_run_step && r_sys_run_step<=9'h174)) begin
										r_sub14_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub14_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp4682[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub14_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h37)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp336[12:0] );

									end
									else
									if((r_sys_run_step==9'h36)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp330[12:0] );

									end
									else
									if((r_sys_run_step==9'h3a)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp354[12:0] );

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp360[12:0] );

									end
									else
									if((r_sys_run_step==9'h2d)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp276[12:0] );

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp288[12:0] );

									end
									else
									if((r_sys_run_step==9'h29)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp252[12:0] );

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp222[12:0] );

									end
									else
									if((r_sys_run_step==9'h34)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp318[12:0] );

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp372[12:0] );

									end
									else
									if((r_sys_run_step==9'h42)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp402[12:0] );

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp228[12:0] );

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp348[12:0] );

									end
									else
									if((r_sys_run_step==9'h43)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp408[12:0] );

									end
									else
									if((r_sys_run_step==9'h38)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp342[12:0] );

									end
									else
									if((r_sys_run_step==9'h26)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp234[12:0] );

									end
									else
									if((r_sys_run_step==9'h32)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp306[12:0] );

									end
									else
									if((r_sys_run_step==9'h2e)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp282[12:0] );

									end
									else
									if((r_sys_run_step==9'h23)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp216[12:0] );

									end
									else
									if((r_sys_run_step==9'h2c)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp270[12:0] );

									end
									else
									if((r_sys_run_step==9'h31)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp300[12:0] );

									end
									else
									if((r_sys_run_step==9'h33)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp312[12:0] );

									end
									else
									if((r_sys_run_step==9'h28)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp246[12:0] );

									end
									else
									if((r_sys_run_step==9'h41)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp396[12:0] );

									end
									else
									if((r_sys_run_step==9'h3f)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp384[12:0] );

									end
									else
									if((r_sys_run_step==9'h2b)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp264[12:0] );

									end
									else
									if((r_sys_run_step==9'h40)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp390[12:0] );

									end
									else
									if((r_sys_run_step==9'h35)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp324[12:0] );

									end
									else
									if((r_sys_run_step==9'h3e)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp378[12:0] );

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp366[12:0] );

									end
									else
									if((r_sys_run_step==9'h2a)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp258[12:0] );

									end
									else
									if((r_sys_run_step==9'h30)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp294[12:0] );

									end
									else
									if((r_sys_run_step==9'h27)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp240[12:0] );

									end
									else
									if((r_sys_run_step==9'h44)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp429[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h23<=r_sys_run_step && r_sys_run_step<=9'h44)) begin
										r_sub01_u_datain <= w_sys_tmp218;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h23<=r_sys_run_step && r_sys_run_step<=9'h44)) begin
										r_sub01_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub01_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3552[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'ha: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub13_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub13_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h150)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2838[12:0] );

									end
									else
									if((r_sys_run_step==9'h13b)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2712[12:0] );

									end
									else
									if((r_sys_run_step==9'h13e)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2730[12:0] );

									end
									else
									if((r_sys_run_step==9'h139)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2700[12:0] );

									end
									else
									if((r_sys_run_step==9'h14e)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2826[12:0] );

									end
									else
									if((r_sys_run_step==9'h134)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2670[12:0] );

									end
									else
									if((r_sys_run_step==9'h141)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2748[12:0] );

									end
									else
									if((r_sys_run_step==9'h144)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2766[12:0] );

									end
									else
									if((r_sys_run_step==9'h13a)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2706[12:0] );

									end
									else
									if((r_sys_run_step==9'h13f)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2736[12:0] );

									end
									else
									if((r_sys_run_step==9'h138)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2694[12:0] );

									end
									else
									if((r_sys_run_step==9'h131)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2652[12:0] );

									end
									else
									if((r_sys_run_step==9'h14a)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2802[12:0] );

									end
									else
									if((r_sys_run_step==9'h152)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2865[12:0] );

									end
									else
									if((r_sys_run_step==9'h137)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2688[12:0] );

									end
									else
									if((r_sys_run_step==9'h13c)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2718[12:0] );

									end
									else
									if((r_sys_run_step==9'h133)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2664[12:0] );

									end
									else
									if((r_sys_run_step==9'h14f)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2832[12:0] );

									end
									else
									if((r_sys_run_step==9'h14b)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2808[12:0] );

									end
									else
									if((r_sys_run_step==9'h140)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2742[12:0] );

									end
									else
									if((r_sys_run_step==9'h136)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2682[12:0] );

									end
									else
									if((r_sys_run_step==9'h142)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2754[12:0] );

									end
									else
									if((r_sys_run_step==9'h145)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2772[12:0] );

									end
									else
									if((r_sys_run_step==9'h14d)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2820[12:0] );

									end
									else
									if((r_sys_run_step==9'h149)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2796[12:0] );

									end
									else
									if((r_sys_run_step==9'h147)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2784[12:0] );

									end
									else
									if((r_sys_run_step==9'h143)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2760[12:0] );

									end
									else
									if((r_sys_run_step==9'h148)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2790[12:0] );

									end
									else
									if((r_sys_run_step==9'h135)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2676[12:0] );

									end
									else
									if((r_sys_run_step==9'h146)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2778[12:0] );

									end
									else
									if((r_sys_run_step==9'h14c)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2814[12:0] );

									end
									else
									if((r_sys_run_step==9'h13d)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2724[12:0] );

									end
									else
									if((r_sys_run_step==9'h132)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2658[12:0] );

									end
									else
									if((r_sys_run_step==9'h151)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2844[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h131<=r_sys_run_step && r_sys_run_step<=9'h152)) begin
										r_sub13_u_datain <= w_sys_tmp1034;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h131<=r_sys_run_step && r_sys_run_step<=9'h152)) begin
										r_sub13_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub13_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp4593[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub13_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h16)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp336[12:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp330[12:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp354[12:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp360[12:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp276[12:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp288[12:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp252[12:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp222[12:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp318[12:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp372[12:0] );

									end
									else
									if((r_sys_run_step==9'h21)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp402[12:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp228[12:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp348[12:0] );

									end
									else
									if((r_sys_run_step==9'h22)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp408[12:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp342[12:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp234[12:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp306[12:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp282[12:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp216[12:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp270[12:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp300[12:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp312[12:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp246[12:0] );

									end
									else
									if((r_sys_run_step==9'h20)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp396[12:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp384[12:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp264[12:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp390[12:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp324[12:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp378[12:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp366[12:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp258[12:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp294[12:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp240[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h22)) begin
										r_sub00_u_datain <= w_sys_tmp218;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h22)) begin
										r_sub00_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub00_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3477[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'h6: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub07_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub07_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h79)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1140[12:0] );

									end
									else
									if((r_sys_run_step==9'h6c)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1062[12:0] );

									end
									else
									if((r_sys_run_step==9'h7f)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1176[12:0] );

									end
									else
									if((r_sys_run_step==9'h81)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1188[12:0] );

									end
									else
									if((r_sys_run_step==9'h84)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1206[12:0] );

									end
									else
									if((r_sys_run_step==9'h73)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1104[12:0] );

									end
									else
									if((r_sys_run_step==9'h74)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1110[12:0] );

									end
									else
									if((r_sys_run_step==9'h7b)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1152[12:0] );

									end
									else
									if((r_sys_run_step==9'h6f)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1080[12:0] );

									end
									else
									if((r_sys_run_step==9'h7d)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1164[12:0] );

									end
									else
									if((r_sys_run_step==9'h88)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1245[12:0] );

									end
									else
									if((r_sys_run_step==9'h87)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1224[12:0] );

									end
									else
									if((r_sys_run_step==9'h86)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1218[12:0] );

									end
									else
									if((r_sys_run_step==9'h71)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1092[12:0] );

									end
									else
									if((r_sys_run_step==9'h72)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1098[12:0] );

									end
									else
									if((r_sys_run_step==9'h85)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1212[12:0] );

									end
									else
									if((r_sys_run_step==9'h7c)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1158[12:0] );

									end
									else
									if((r_sys_run_step==9'h83)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1200[12:0] );

									end
									else
									if((r_sys_run_step==9'h6d)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1068[12:0] );

									end
									else
									if((r_sys_run_step==9'h7e)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1170[12:0] );

									end
									else
									if((r_sys_run_step==9'h78)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1134[12:0] );

									end
									else
									if((r_sys_run_step==9'h70)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1086[12:0] );

									end
									else
									if((r_sys_run_step==9'h77)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1128[12:0] );

									end
									else
									if((r_sys_run_step==9'h6a)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1050[12:0] );

									end
									else
									if((r_sys_run_step==9'h76)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1122[12:0] );

									end
									else
									if((r_sys_run_step==9'h67)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1032[12:0] );

									end
									else
									if((r_sys_run_step==9'h7a)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1146[12:0] );

									end
									else
									if((r_sys_run_step==9'h82)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1194[12:0] );

									end
									else
									if((r_sys_run_step==9'h75)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1116[12:0] );

									end
									else
									if((r_sys_run_step==9'h6b)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1056[12:0] );

									end
									else
									if((r_sys_run_step==9'h6e)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1074[12:0] );

									end
									else
									if((r_sys_run_step==9'h68)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1038[12:0] );

									end
									else
									if((r_sys_run_step==9'h69)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1044[12:0] );

									end
									else
									if((r_sys_run_step==9'h80)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1182[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h67<=r_sys_run_step && r_sys_run_step<=9'h88)) begin
										r_sub07_u_datain <= w_sys_tmp1034;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h67<=r_sys_run_step && r_sys_run_step<=9'h88)) begin
										r_sub07_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub07_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h61: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4077[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h61: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub07_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'h5: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub06_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub06_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h57)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1140[12:0] );

									end
									else
									if((r_sys_run_step==9'h4a)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1062[12:0] );

									end
									else
									if((r_sys_run_step==9'h5d)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1176[12:0] );

									end
									else
									if((r_sys_run_step==9'h5f)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1188[12:0] );

									end
									else
									if((r_sys_run_step==9'h62)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1206[12:0] );

									end
									else
									if((r_sys_run_step==9'h51)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1104[12:0] );

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1110[12:0] );

									end
									else
									if((r_sys_run_step==9'h59)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1152[12:0] );

									end
									else
									if((r_sys_run_step==9'h4d)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1080[12:0] );

									end
									else
									if((r_sys_run_step==9'h5b)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1164[12:0] );

									end
									else
									if((r_sys_run_step==9'h66)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1245[12:0] );

									end
									else
									if((r_sys_run_step==9'h65)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1224[12:0] );

									end
									else
									if((r_sys_run_step==9'h64)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1218[12:0] );

									end
									else
									if((r_sys_run_step==9'h4f)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1092[12:0] );

									end
									else
									if((r_sys_run_step==9'h50)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1098[12:0] );

									end
									else
									if((r_sys_run_step==9'h63)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1212[12:0] );

									end
									else
									if((r_sys_run_step==9'h5a)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1158[12:0] );

									end
									else
									if((r_sys_run_step==9'h61)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1200[12:0] );

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1068[12:0] );

									end
									else
									if((r_sys_run_step==9'h5c)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1170[12:0] );

									end
									else
									if((r_sys_run_step==9'h56)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1134[12:0] );

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1086[12:0] );

									end
									else
									if((r_sys_run_step==9'h55)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1128[12:0] );

									end
									else
									if((r_sys_run_step==9'h48)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1050[12:0] );

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1122[12:0] );

									end
									else
									if((r_sys_run_step==9'h45)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1032[12:0] );

									end
									else
									if((r_sys_run_step==9'h58)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1146[12:0] );

									end
									else
									if((r_sys_run_step==9'h60)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1194[12:0] );

									end
									else
									if((r_sys_run_step==9'h53)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1116[12:0] );

									end
									else
									if((r_sys_run_step==9'h49)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1056[12:0] );

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1074[12:0] );

									end
									else
									if((r_sys_run_step==9'h46)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1038[12:0] );

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1044[12:0] );

									end
									else
									if((r_sys_run_step==9'h5e)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1182[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h45<=r_sys_run_step && r_sys_run_step<=9'h66)) begin
										r_sub06_u_datain <= w_sys_tmp1034;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h45<=r_sys_run_step && r_sys_run_step<=9'h66)) begin
										r_sub06_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub06_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h5b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp3988[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h5b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub06_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'hc: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub15_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub15_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h194)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2838[12:0] );

									end
									else
									if((r_sys_run_step==9'h17f)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2712[12:0] );

									end
									else
									if((r_sys_run_step==9'h182)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2730[12:0] );

									end
									else
									if((r_sys_run_step==9'h17d)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2700[12:0] );

									end
									else
									if((r_sys_run_step==9'h192)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2826[12:0] );

									end
									else
									if((r_sys_run_step==9'h178)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2670[12:0] );

									end
									else
									if((r_sys_run_step==9'h185)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2748[12:0] );

									end
									else
									if((r_sys_run_step==9'h188)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2766[12:0] );

									end
									else
									if((r_sys_run_step==9'h17e)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2706[12:0] );

									end
									else
									if((r_sys_run_step==9'h183)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2736[12:0] );

									end
									else
									if((r_sys_run_step==9'h17c)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2694[12:0] );

									end
									else
									if((r_sys_run_step==9'h175)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2652[12:0] );

									end
									else
									if((r_sys_run_step==9'h18e)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2802[12:0] );

									end
									else
									if((r_sys_run_step==9'h196)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2865[12:0] );

									end
									else
									if((r_sys_run_step==9'h17b)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2688[12:0] );

									end
									else
									if((r_sys_run_step==9'h180)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2718[12:0] );

									end
									else
									if((r_sys_run_step==9'h177)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2664[12:0] );

									end
									else
									if((r_sys_run_step==9'h193)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2832[12:0] );

									end
									else
									if((r_sys_run_step==9'h18f)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2808[12:0] );

									end
									else
									if((r_sys_run_step==9'h184)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2742[12:0] );

									end
									else
									if((r_sys_run_step==9'h17a)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2682[12:0] );

									end
									else
									if((r_sys_run_step==9'h186)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2754[12:0] );

									end
									else
									if((r_sys_run_step==9'h189)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2772[12:0] );

									end
									else
									if((r_sys_run_step==9'h191)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2820[12:0] );

									end
									else
									if((r_sys_run_step==9'h18d)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2796[12:0] );

									end
									else
									if((r_sys_run_step==9'h18b)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2784[12:0] );

									end
									else
									if((r_sys_run_step==9'h187)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2760[12:0] );

									end
									else
									if((r_sys_run_step==9'h18c)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2790[12:0] );

									end
									else
									if((r_sys_run_step==9'h179)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2676[12:0] );

									end
									else
									if((r_sys_run_step==9'h18a)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2778[12:0] );

									end
									else
									if((r_sys_run_step==9'h190)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2814[12:0] );

									end
									else
									if((r_sys_run_step==9'h181)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2724[12:0] );

									end
									else
									if((r_sys_run_step==9'h176)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2658[12:0] );

									end
									else
									if((r_sys_run_step==9'h195)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp2844[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h175<=r_sys_run_step && r_sys_run_step<=9'h196)) begin
										r_sub15_u_datain <= w_sys_tmp1034;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h175<=r_sys_run_step && r_sys_run_step<=9'h196)) begin
										r_sub15_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub15_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp4771[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub15_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'h4: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub05_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub05_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h35)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1140[12:0] );

									end
									else
									if((r_sys_run_step==9'h28)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1062[12:0] );

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1176[12:0] );

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1188[12:0] );

									end
									else
									if((r_sys_run_step==9'h40)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1206[12:0] );

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1104[12:0] );

									end
									else
									if((r_sys_run_step==9'h30)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1110[12:0] );

									end
									else
									if((r_sys_run_step==9'h37)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1152[12:0] );

									end
									else
									if((r_sys_run_step==9'h2b)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1080[12:0] );

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1164[12:0] );

									end
									else
									if((r_sys_run_step==9'h44)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1245[12:0] );

									end
									else
									if((r_sys_run_step==9'h43)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1224[12:0] );

									end
									else
									if((r_sys_run_step==9'h42)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1218[12:0] );

									end
									else
									if((r_sys_run_step==9'h2d)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1092[12:0] );

									end
									else
									if((r_sys_run_step==9'h2e)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1098[12:0] );

									end
									else
									if((r_sys_run_step==9'h41)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1212[12:0] );

									end
									else
									if((r_sys_run_step==9'h38)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1158[12:0] );

									end
									else
									if((r_sys_run_step==9'h3f)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1200[12:0] );

									end
									else
									if((r_sys_run_step==9'h29)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1068[12:0] );

									end
									else
									if((r_sys_run_step==9'h3a)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1170[12:0] );

									end
									else
									if((r_sys_run_step==9'h34)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1134[12:0] );

									end
									else
									if((r_sys_run_step==9'h2c)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1086[12:0] );

									end
									else
									if((r_sys_run_step==9'h33)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1128[12:0] );

									end
									else
									if((r_sys_run_step==9'h26)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1050[12:0] );

									end
									else
									if((r_sys_run_step==9'h32)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1122[12:0] );

									end
									else
									if((r_sys_run_step==9'h23)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1032[12:0] );

									end
									else
									if((r_sys_run_step==9'h36)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1146[12:0] );

									end
									else
									if((r_sys_run_step==9'h3e)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1194[12:0] );

									end
									else
									if((r_sys_run_step==9'h31)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1116[12:0] );

									end
									else
									if((r_sys_run_step==9'h27)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1056[12:0] );

									end
									else
									if((r_sys_run_step==9'h2a)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1074[12:0] );

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1038[12:0] );

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1044[12:0] );

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1182[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h23<=r_sys_run_step && r_sys_run_step<=9'h44)) begin
										r_sub05_u_datain <= w_sys_tmp1034;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h23<=r_sys_run_step && r_sys_run_step<=9'h44)) begin
										r_sub05_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub05_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h55: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp3899[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h55: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub05_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'he: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub04_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub04_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1140[12:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1062[12:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1176[12:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1188[12:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1206[12:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1104[12:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1110[12:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1152[12:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1080[12:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1164[12:0] );

									end
									else
									if((r_sys_run_step==9'h22)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1224[12:0] );

									end
									else
									if((r_sys_run_step==9'h21)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1218[12:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1092[12:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1098[12:0] );

									end
									else
									if((r_sys_run_step==9'h20)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1212[12:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1158[12:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1200[12:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1068[12:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1170[12:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1134[12:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1086[12:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1128[12:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1050[12:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1122[12:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1032[12:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1146[12:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1194[12:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1116[12:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1056[12:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1074[12:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1038[12:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1044[12:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1182[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h22)) begin
										r_sub04_u_datain <= w_sys_tmp1034;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h22)) begin
										r_sub04_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub04_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h4f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp3824[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h4f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub04_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'h8: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub10_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub10_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he9)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2016[12:0] );

									end
									else
									if((r_sys_run_step==9'hea)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2022[12:0] );

									end
									else
									if((r_sys_run_step==9'hd9)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp1920[12:0] );

									end
									else
									if((r_sys_run_step==9'hdd)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp1944[12:0] );

									end
									else
									if((r_sys_run_step==9'hd0)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp1866[12:0] );

									end
									else
									if((r_sys_run_step==9'hd3)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp1884[12:0] );

									end
									else
									if((r_sys_run_step==9'he0)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp1962[12:0] );

									end
									else
									if((r_sys_run_step==9'hd7)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp1908[12:0] );

									end
									else
									if((r_sys_run_step==9'hed)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2055[12:0] );

									end
									else
									if((r_sys_run_step==9'hd4)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp1890[12:0] );

									end
									else
									if((r_sys_run_step==9'hdb)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp1932[12:0] );

									end
									else
									if((r_sys_run_step==9'hd5)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp1896[12:0] );

									end
									else
									if((r_sys_run_step==9'hec)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2034[12:0] );

									end
									else
									if((r_sys_run_step==9'hda)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp1926[12:0] );

									end
									else
									if((r_sys_run_step==9'hcc)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp1842[12:0] );

									end
									else
									if((r_sys_run_step==9'hdf)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp1956[12:0] );

									end
									else
									if((r_sys_run_step==9'hd1)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp1872[12:0] );

									end
									else
									if((r_sys_run_step==9'he5)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp1992[12:0] );

									end
									else
									if((r_sys_run_step==9'hd2)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp1878[12:0] );

									end
									else
									if((r_sys_run_step==9'hd6)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp1902[12:0] );

									end
									else
									if((r_sys_run_step==9'hd8)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp1914[12:0] );

									end
									else
									if((r_sys_run_step==9'hdc)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp1938[12:0] );

									end
									else
									if((r_sys_run_step==9'he2)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp1974[12:0] );

									end
									else
									if((r_sys_run_step==9'hce)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp1854[12:0] );

									end
									else
									if((r_sys_run_step==9'he7)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2004[12:0] );

									end
									else
									if((r_sys_run_step==9'he6)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp1998[12:0] );

									end
									else
									if((r_sys_run_step==9'he3)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp1980[12:0] );

									end
									else
									if((r_sys_run_step==9'he4)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp1986[12:0] );

									end
									else
									if((r_sys_run_step==9'heb)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2028[12:0] );

									end
									else
									if((r_sys_run_step==9'hcd)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp1848[12:0] );

									end
									else
									if((r_sys_run_step==9'he1)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp1968[12:0] );

									end
									else
									if((r_sys_run_step==9'hde)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp1950[12:0] );

									end
									else
									if((r_sys_run_step==9'he8)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2010[12:0] );

									end
									else
									if((r_sys_run_step==9'hcf)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp1860[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'hcc<=r_sys_run_step && r_sys_run_step<=9'hed)) begin
										r_sub10_u_datain <= w_sys_tmp1034;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'hcc<=r_sys_run_step && r_sys_run_step<=9'hed)) begin
										r_sub10_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub10_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h78: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp4335[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						8'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h78: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						8'h9d: begin
							r_sub10_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


endmodule
