/*
TimeStamp:	2016/10/19		18:57
*/


module c1(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy	
);

	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 8:0] r_sys_run_phase;
	reg         [ 4:0] r_sys_run_stage;
	reg         [ 6:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 4:0] w_sys_run_stage_p1;
	wire        [ 6:0] w_sys_run_step_p1;
	wire signed [14:0] w_fld_u_0_addr_0;
	wire        [31:0] w_fld_u_0_datain_0;
	wire        [31:0] w_fld_u_0_dataout_0;
	wire               w_fld_u_0_r_w_0;
	wire               w_fld_u_0_ce_0;
	reg  signed [14:0] r_fld_u_0_addr_1;
	reg         [31:0] r_fld_u_0_datain_1;
	wire        [31:0] w_fld_u_0_dataout_1;
	reg                r_fld_u_0_r_w_1;
	wire               w_fld_u_0_ce_1;
	reg  signed [31:0] r_run_k_17;
	reg  signed [31:0] r_run_j_18;
	reg  signed [31:0] r_run_n_19;
	reg  signed [31:0] r_run_mx_20;
	reg  signed [31:0] r_run_my_21;
	reg  signed [31:0] r_run_nlast_22;
	reg  signed [31:0] r_run_tmpj_23;
	reg  signed [31:0] r_run_copy0_j_24;
	reg  signed [31:0] r_run_copy0_j_25;
	reg  signed [31:0] r_run_copy0_j_26;
	reg  signed [31:0] r_run_copy0_j_27;
	reg  signed [31:0] r_run_copy0_j_28;
	reg  signed [31:0] r_run_copy0_j_29;
	reg  signed [31:0] r_run_copy0_j_30;
	reg  signed [31:0] r_run_copy0_j_31;
	reg  signed [31:0] r_run_copy0_j_32;
	reg  signed [31:0] r_run_copy0_j_33;
	reg  signed [31:0] r_run_copy0_j_34;
	reg  signed [31:0] r_run_copy0_j_35;
	reg  signed [31:0] r_run_copy0_j_36;
	reg  signed [31:0] r_run_copy0_j_37;
	reg  signed [31:0] r_run_copy0_j_38;
	reg  signed [31:0] r_run_copy0_j_39;
	reg  signed [31:0] r_run_copy0_j_40;
	reg  signed [31:0] r_run_copy1_j_41;
	reg  signed [31:0] r_run_copy2_j_42;
	reg  signed [31:0] r_run_copy3_j_43;
	reg  signed [31:0] r_run_copy4_j_44;
	reg  signed [31:0] r_run_copy5_j_45;
	reg  signed [31:0] r_run_copy6_j_46;
	reg  signed [31:0] r_run_copy7_j_47;
	reg  signed [31:0] r_run_copy8_j_48;
	reg  signed [31:0] r_run_copy9_j_49;
	reg  signed [31:0] r_run_copy10_j_50;
	reg  signed [31:0] r_run_copy0_j_51;
	reg  signed [31:0] r_run_copy0_j_52;
	reg  signed [31:0] r_run_copy1_j_53;
	reg  signed [31:0] r_run_copy0_j_54;
	reg  signed [31:0] r_run_copy1_j_55;
	reg  signed [31:0] r_run_copy0_j_56;
	reg  signed [31:0] r_run_copy1_j_57;
	reg  signed [31:0] r_run_copy0_j_58;
	reg  signed [31:0] r_run_copy0_j_59;
	reg  signed [31:0] r_run_copy1_j_60;
	reg  signed [31:0] r_run_copy0_j_61;
	reg  signed [31:0] r_run_copy1_j_62;
	reg  signed [31:0] r_run_copy0_j_63;
	reg  signed [31:0] r_run_copy1_j_64;
	reg  signed [31:0] r_run_copy0_j_65;
	reg  signed [31:0] r_run_copy0_j_66;
	reg  signed [31:0] r_run_copy1_j_67;
	reg  signed [31:0] r_run_copy0_j_68;
	reg  signed [31:0] r_run_copy1_j_69;
	reg  signed [31:0] r_run_copy0_j_70;
	reg  signed [31:0] r_run_copy1_j_71;
	reg  signed [31:0] r_run_copy0_j_72;
	reg  signed [31:0] r_run_copy0_j_73;
	reg  signed [31:0] r_run_copy1_j_74;
	reg  signed [31:0] r_run_copy0_j_75;
	reg  signed [31:0] r_run_copy1_j_76;
	reg  signed [31:0] r_run_copy0_j_77;
	reg  signed [31:0] r_run_copy1_j_78;
	reg                r_sub09_run_req;
	wire               w_sub09_run_busy;
	wire signed [12:0] w_sub09_u_addr;
	reg  signed [12:0] r_sub09_u_addr;
	wire        [31:0] w_sub09_u_datain;
	reg         [31:0] r_sub09_u_datain;
	wire        [31:0] w_sub09_u_dataout;
	wire               w_sub09_u_r_w;
	reg                r_sub09_u_r_w;
	wire signed [12:0] w_sub09_result_addr;
	reg  signed [12:0] r_sub09_result_addr;
	wire        [31:0] w_sub09_result_datain;
	reg         [31:0] r_sub09_result_datain;
	wire        [31:0] w_sub09_result_dataout;
	wire               w_sub09_result_r_w;
	reg                r_sub09_result_r_w;
	reg                r_sub08_run_req;
	wire               w_sub08_run_busy;
	wire signed [12:0] w_sub08_u_addr;
	reg  signed [12:0] r_sub08_u_addr;
	wire        [31:0] w_sub08_u_datain;
	reg         [31:0] r_sub08_u_datain;
	wire        [31:0] w_sub08_u_dataout;
	wire               w_sub08_u_r_w;
	reg                r_sub08_u_r_w;
	wire signed [12:0] w_sub08_result_addr;
	reg  signed [12:0] r_sub08_result_addr;
	wire        [31:0] w_sub08_result_datain;
	reg         [31:0] r_sub08_result_datain;
	wire        [31:0] w_sub08_result_dataout;
	wire               w_sub08_result_r_w;
	reg                r_sub08_result_r_w;
	reg                r_sub12_run_req;
	wire               w_sub12_run_busy;
	wire signed [12:0] w_sub12_u_addr;
	reg  signed [12:0] r_sub12_u_addr;
	wire        [31:0] w_sub12_u_datain;
	reg         [31:0] r_sub12_u_datain;
	wire        [31:0] w_sub12_u_dataout;
	wire               w_sub12_u_r_w;
	reg                r_sub12_u_r_w;
	wire signed [12:0] w_sub12_result_addr;
	reg  signed [12:0] r_sub12_result_addr;
	wire        [31:0] w_sub12_result_datain;
	reg         [31:0] r_sub12_result_datain;
	wire        [31:0] w_sub12_result_dataout;
	wire               w_sub12_result_r_w;
	reg                r_sub12_result_r_w;
	reg                r_sub03_run_req;
	wire               w_sub03_run_busy;
	wire signed [12:0] w_sub03_u_addr;
	reg  signed [12:0] r_sub03_u_addr;
	wire        [31:0] w_sub03_u_datain;
	reg         [31:0] r_sub03_u_datain;
	wire        [31:0] w_sub03_u_dataout;
	wire               w_sub03_u_r_w;
	reg                r_sub03_u_r_w;
	wire signed [12:0] w_sub03_result_addr;
	reg  signed [12:0] r_sub03_result_addr;
	wire        [31:0] w_sub03_result_datain;
	reg         [31:0] r_sub03_result_datain;
	wire        [31:0] w_sub03_result_dataout;
	wire               w_sub03_result_r_w;
	reg                r_sub03_result_r_w;
	reg                r_sub02_run_req;
	wire               w_sub02_run_busy;
	wire signed [12:0] w_sub02_u_addr;
	reg  signed [12:0] r_sub02_u_addr;
	wire        [31:0] w_sub02_u_datain;
	reg         [31:0] r_sub02_u_datain;
	wire        [31:0] w_sub02_u_dataout;
	wire               w_sub02_u_r_w;
	reg                r_sub02_u_r_w;
	wire signed [12:0] w_sub02_result_addr;
	reg  signed [12:0] r_sub02_result_addr;
	wire        [31:0] w_sub02_result_datain;
	reg         [31:0] r_sub02_result_datain;
	wire        [31:0] w_sub02_result_dataout;
	wire               w_sub02_result_r_w;
	reg                r_sub02_result_r_w;
	reg                r_sub11_run_req;
	wire               w_sub11_run_busy;
	wire signed [12:0] w_sub11_u_addr;
	reg  signed [12:0] r_sub11_u_addr;
	wire        [31:0] w_sub11_u_datain;
	reg         [31:0] r_sub11_u_datain;
	wire        [31:0] w_sub11_u_dataout;
	wire               w_sub11_u_r_w;
	reg                r_sub11_u_r_w;
	wire signed [12:0] w_sub11_result_addr;
	reg  signed [12:0] r_sub11_result_addr;
	wire        [31:0] w_sub11_result_datain;
	reg         [31:0] r_sub11_result_datain;
	wire        [31:0] w_sub11_result_dataout;
	wire               w_sub11_result_r_w;
	reg                r_sub11_result_r_w;
	reg                r_sub14_run_req;
	wire               w_sub14_run_busy;
	wire signed [12:0] w_sub14_u_addr;
	reg  signed [12:0] r_sub14_u_addr;
	wire        [31:0] w_sub14_u_datain;
	reg         [31:0] r_sub14_u_datain;
	wire        [31:0] w_sub14_u_dataout;
	wire               w_sub14_u_r_w;
	reg                r_sub14_u_r_w;
	wire signed [12:0] w_sub14_result_addr;
	reg  signed [12:0] r_sub14_result_addr;
	wire        [31:0] w_sub14_result_datain;
	reg         [31:0] r_sub14_result_datain;
	wire        [31:0] w_sub14_result_dataout;
	wire               w_sub14_result_r_w;
	reg                r_sub14_result_r_w;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [12:0] w_sub01_u_addr;
	reg  signed [12:0] r_sub01_u_addr;
	wire        [31:0] w_sub01_u_datain;
	reg         [31:0] r_sub01_u_datain;
	wire        [31:0] w_sub01_u_dataout;
	wire               w_sub01_u_r_w;
	reg                r_sub01_u_r_w;
	wire signed [12:0] w_sub01_result_addr;
	reg  signed [12:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub13_run_req;
	wire               w_sub13_run_busy;
	wire signed [12:0] w_sub13_u_addr;
	reg  signed [12:0] r_sub13_u_addr;
	wire        [31:0] w_sub13_u_datain;
	reg         [31:0] r_sub13_u_datain;
	wire        [31:0] w_sub13_u_dataout;
	wire               w_sub13_u_r_w;
	reg                r_sub13_u_r_w;
	wire signed [12:0] w_sub13_result_addr;
	reg  signed [12:0] r_sub13_result_addr;
	wire        [31:0] w_sub13_result_datain;
	reg         [31:0] r_sub13_result_datain;
	wire        [31:0] w_sub13_result_dataout;
	wire               w_sub13_result_r_w;
	reg                r_sub13_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [12:0] w_sub00_u_addr;
	reg  signed [12:0] r_sub00_u_addr;
	wire        [31:0] w_sub00_u_datain;
	reg         [31:0] r_sub00_u_datain;
	wire        [31:0] w_sub00_u_dataout;
	wire               w_sub00_u_r_w;
	reg                r_sub00_u_r_w;
	wire signed [12:0] w_sub00_result_addr;
	reg  signed [12:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	reg                r_sub07_run_req;
	wire               w_sub07_run_busy;
	wire signed [12:0] w_sub07_u_addr;
	reg  signed [12:0] r_sub07_u_addr;
	wire        [31:0] w_sub07_u_datain;
	reg         [31:0] r_sub07_u_datain;
	wire        [31:0] w_sub07_u_dataout;
	wire               w_sub07_u_r_w;
	reg                r_sub07_u_r_w;
	wire signed [12:0] w_sub07_result_addr;
	reg  signed [12:0] r_sub07_result_addr;
	wire        [31:0] w_sub07_result_datain;
	reg         [31:0] r_sub07_result_datain;
	wire        [31:0] w_sub07_result_dataout;
	wire               w_sub07_result_r_w;
	reg                r_sub07_result_r_w;
	reg                r_sub06_run_req;
	wire               w_sub06_run_busy;
	wire signed [12:0] w_sub06_u_addr;
	reg  signed [12:0] r_sub06_u_addr;
	wire        [31:0] w_sub06_u_datain;
	reg         [31:0] r_sub06_u_datain;
	wire        [31:0] w_sub06_u_dataout;
	wire               w_sub06_u_r_w;
	reg                r_sub06_u_r_w;
	wire signed [12:0] w_sub06_result_addr;
	reg  signed [12:0] r_sub06_result_addr;
	wire        [31:0] w_sub06_result_datain;
	reg         [31:0] r_sub06_result_datain;
	wire        [31:0] w_sub06_result_dataout;
	wire               w_sub06_result_r_w;
	reg                r_sub06_result_r_w;
	reg                r_sub15_run_req;
	wire               w_sub15_run_busy;
	wire signed [12:0] w_sub15_u_addr;
	reg  signed [12:0] r_sub15_u_addr;
	wire        [31:0] w_sub15_u_datain;
	reg         [31:0] r_sub15_u_datain;
	wire        [31:0] w_sub15_u_dataout;
	wire               w_sub15_u_r_w;
	reg                r_sub15_u_r_w;
	wire signed [12:0] w_sub15_result_addr;
	reg  signed [12:0] r_sub15_result_addr;
	wire        [31:0] w_sub15_result_datain;
	reg         [31:0] r_sub15_result_datain;
	wire        [31:0] w_sub15_result_dataout;
	wire               w_sub15_result_r_w;
	reg                r_sub15_result_r_w;
	reg                r_sub05_run_req;
	wire               w_sub05_run_busy;
	wire signed [12:0] w_sub05_u_addr;
	reg  signed [12:0] r_sub05_u_addr;
	wire        [31:0] w_sub05_u_datain;
	reg         [31:0] r_sub05_u_datain;
	wire        [31:0] w_sub05_u_dataout;
	wire               w_sub05_u_r_w;
	reg                r_sub05_u_r_w;
	wire signed [12:0] w_sub05_result_addr;
	reg  signed [12:0] r_sub05_result_addr;
	wire        [31:0] w_sub05_result_datain;
	reg         [31:0] r_sub05_result_datain;
	wire        [31:0] w_sub05_result_dataout;
	wire               w_sub05_result_r_w;
	reg                r_sub05_result_r_w;
	reg                r_sub04_run_req;
	wire               w_sub04_run_busy;
	wire signed [12:0] w_sub04_u_addr;
	reg  signed [12:0] r_sub04_u_addr;
	wire        [31:0] w_sub04_u_datain;
	reg         [31:0] r_sub04_u_datain;
	wire        [31:0] w_sub04_u_dataout;
	wire               w_sub04_u_r_w;
	reg                r_sub04_u_r_w;
	wire signed [12:0] w_sub04_result_addr;
	reg  signed [12:0] r_sub04_result_addr;
	wire        [31:0] w_sub04_result_datain;
	reg         [31:0] r_sub04_result_datain;
	wire        [31:0] w_sub04_result_dataout;
	wire               w_sub04_result_r_w;
	reg                r_sub04_result_r_w;
	reg                r_sub10_run_req;
	wire               w_sub10_run_busy;
	wire signed [12:0] w_sub10_u_addr;
	reg  signed [12:0] r_sub10_u_addr;
	wire        [31:0] w_sub10_u_datain;
	reg         [31:0] r_sub10_u_datain;
	wire        [31:0] w_sub10_u_dataout;
	wire               w_sub10_u_r_w;
	reg                r_sub10_u_r_w;
	wire signed [12:0] w_sub10_result_addr;
	reg  signed [12:0] r_sub10_result_addr;
	wire        [31:0] w_sub10_result_datain;
	reg         [31:0] r_sub10_result_datain;
	wire        [31:0] w_sub10_result_dataout;
	wire               w_sub10_result_r_w;
	reg                r_sub10_result_r_w;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	wire signed [31:0] w_sys_tmp1;
	wire signed [31:0] w_sys_tmp3;
	wire               w_sys_tmp4;
	wire               w_sys_tmp5;
	wire signed [31:0] w_sys_tmp6;
	wire               w_sys_tmp7;
	wire               w_sys_tmp8;
	wire signed [31:0] w_sys_tmp11;
	wire signed [31:0] w_sys_tmp12;
	wire signed [31:0] w_sys_tmp13;
	wire        [31:0] w_sys_tmp14;
	wire signed [31:0] w_sys_tmp15;
	wire               w_sys_tmp52;
	wire               w_sys_tmp53;
	wire signed [31:0] w_sys_tmp54;
	wire signed [31:0] w_sys_tmp55;
	wire               w_sys_tmp56;
	wire               w_sys_tmp57;
	wire signed [31:0] w_sys_tmp58;
	wire signed [31:0] w_sys_tmp61;
	wire signed [31:0] w_sys_tmp62;
	wire signed [31:0] w_sys_tmp63;
	wire        [31:0] w_sys_tmp64;
	wire signed [31:0] w_sys_tmp65;
	wire signed [31:0] w_sys_tmp66;
	wire signed [31:0] w_sys_tmp68;
	wire signed [31:0] w_sys_tmp69;
	wire signed [31:0] w_sys_tmp130;
	wire               w_sys_tmp131;
	wire               w_sys_tmp132;
	wire signed [31:0] w_sys_tmp133;
	wire signed [31:0] w_sys_tmp135;
	wire signed [31:0] w_sys_tmp136;
	wire signed [31:0] w_sys_tmp138;
	wire signed [31:0] w_sys_tmp139;
	wire signed [31:0] w_sys_tmp140;
	wire        [31:0] w_sys_tmp141;
	wire signed [31:0] w_sys_tmp142;
	wire signed [31:0] w_sys_tmp143;
	wire signed [31:0] w_sys_tmp145;
	wire signed [31:0] w_sys_tmp146;
	wire signed [31:0] w_sys_tmp219;
	wire               w_sys_tmp220;
	wire               w_sys_tmp221;
	wire signed [31:0] w_sys_tmp222;
	wire signed [31:0] w_sys_tmp224;
	wire signed [31:0] w_sys_tmp225;
	wire signed [31:0] w_sys_tmp227;
	wire signed [31:0] w_sys_tmp228;
	wire signed [31:0] w_sys_tmp229;
	wire        [31:0] w_sys_tmp230;
	wire signed [31:0] w_sys_tmp231;
	wire signed [31:0] w_sys_tmp232;
	wire signed [31:0] w_sys_tmp234;
	wire signed [31:0] w_sys_tmp235;
	wire signed [31:0] w_sys_tmp308;
	wire               w_sys_tmp309;
	wire               w_sys_tmp310;
	wire signed [31:0] w_sys_tmp311;
	wire signed [31:0] w_sys_tmp313;
	wire signed [31:0] w_sys_tmp314;
	wire signed [31:0] w_sys_tmp316;
	wire signed [31:0] w_sys_tmp317;
	wire signed [31:0] w_sys_tmp318;
	wire        [31:0] w_sys_tmp319;
	wire signed [31:0] w_sys_tmp320;
	wire signed [31:0] w_sys_tmp321;
	wire signed [31:0] w_sys_tmp323;
	wire signed [31:0] w_sys_tmp324;
	wire signed [31:0] w_sys_tmp397;
	wire               w_sys_tmp398;
	wire               w_sys_tmp399;
	wire signed [31:0] w_sys_tmp400;
	wire signed [31:0] w_sys_tmp401;
	wire               w_sys_tmp402;
	wire               w_sys_tmp403;
	wire signed [31:0] w_sys_tmp404;
	wire signed [31:0] w_sys_tmp407;
	wire signed [31:0] w_sys_tmp408;
	wire signed [31:0] w_sys_tmp409;
	wire        [31:0] w_sys_tmp410;
	wire signed [31:0] w_sys_tmp411;
	wire signed [31:0] w_sys_tmp412;
	wire signed [31:0] w_sys_tmp414;
	wire signed [31:0] w_sys_tmp415;
	wire signed [31:0] w_sys_tmp476;
	wire               w_sys_tmp477;
	wire               w_sys_tmp478;
	wire signed [31:0] w_sys_tmp479;
	wire signed [31:0] w_sys_tmp481;
	wire signed [31:0] w_sys_tmp482;
	wire signed [31:0] w_sys_tmp484;
	wire signed [31:0] w_sys_tmp485;
	wire signed [31:0] w_sys_tmp486;
	wire        [31:0] w_sys_tmp487;
	wire signed [31:0] w_sys_tmp488;
	wire signed [31:0] w_sys_tmp489;
	wire signed [31:0] w_sys_tmp491;
	wire signed [31:0] w_sys_tmp492;
	wire signed [31:0] w_sys_tmp565;
	wire               w_sys_tmp566;
	wire               w_sys_tmp567;
	wire signed [31:0] w_sys_tmp568;
	wire signed [31:0] w_sys_tmp570;
	wire signed [31:0] w_sys_tmp571;
	wire signed [31:0] w_sys_tmp573;
	wire signed [31:0] w_sys_tmp574;
	wire signed [31:0] w_sys_tmp575;
	wire        [31:0] w_sys_tmp576;
	wire signed [31:0] w_sys_tmp577;
	wire signed [31:0] w_sys_tmp578;
	wire signed [31:0] w_sys_tmp580;
	wire signed [31:0] w_sys_tmp581;
	wire signed [31:0] w_sys_tmp654;
	wire               w_sys_tmp655;
	wire               w_sys_tmp656;
	wire signed [31:0] w_sys_tmp657;
	wire signed [31:0] w_sys_tmp659;
	wire signed [31:0] w_sys_tmp660;
	wire signed [31:0] w_sys_tmp662;
	wire signed [31:0] w_sys_tmp663;
	wire signed [31:0] w_sys_tmp664;
	wire        [31:0] w_sys_tmp665;
	wire signed [31:0] w_sys_tmp666;
	wire signed [31:0] w_sys_tmp667;
	wire signed [31:0] w_sys_tmp669;
	wire signed [31:0] w_sys_tmp670;
	wire signed [31:0] w_sys_tmp743;
	wire               w_sys_tmp744;
	wire               w_sys_tmp745;
	wire signed [31:0] w_sys_tmp746;
	wire signed [31:0] w_sys_tmp747;
	wire               w_sys_tmp748;
	wire               w_sys_tmp749;
	wire signed [31:0] w_sys_tmp750;
	wire signed [31:0] w_sys_tmp753;
	wire signed [31:0] w_sys_tmp754;
	wire signed [31:0] w_sys_tmp755;
	wire        [31:0] w_sys_tmp756;
	wire signed [31:0] w_sys_tmp757;
	wire signed [31:0] w_sys_tmp758;
	wire signed [31:0] w_sys_tmp760;
	wire signed [31:0] w_sys_tmp761;
	wire signed [31:0] w_sys_tmp822;
	wire               w_sys_tmp823;
	wire               w_sys_tmp824;
	wire signed [31:0] w_sys_tmp825;
	wire signed [31:0] w_sys_tmp827;
	wire signed [31:0] w_sys_tmp828;
	wire signed [31:0] w_sys_tmp830;
	wire signed [31:0] w_sys_tmp831;
	wire signed [31:0] w_sys_tmp832;
	wire        [31:0] w_sys_tmp833;
	wire signed [31:0] w_sys_tmp834;
	wire signed [31:0] w_sys_tmp835;
	wire signed [31:0] w_sys_tmp837;
	wire signed [31:0] w_sys_tmp838;
	wire signed [31:0] w_sys_tmp911;
	wire               w_sys_tmp912;
	wire               w_sys_tmp913;
	wire signed [31:0] w_sys_tmp914;
	wire signed [31:0] w_sys_tmp916;
	wire signed [31:0] w_sys_tmp917;
	wire signed [31:0] w_sys_tmp919;
	wire signed [31:0] w_sys_tmp920;
	wire signed [31:0] w_sys_tmp921;
	wire        [31:0] w_sys_tmp922;
	wire signed [31:0] w_sys_tmp923;
	wire signed [31:0] w_sys_tmp924;
	wire signed [31:0] w_sys_tmp926;
	wire signed [31:0] w_sys_tmp927;
	wire signed [31:0] w_sys_tmp1000;
	wire               w_sys_tmp1001;
	wire               w_sys_tmp1002;
	wire signed [31:0] w_sys_tmp1003;
	wire signed [31:0] w_sys_tmp1005;
	wire signed [31:0] w_sys_tmp1006;
	wire signed [31:0] w_sys_tmp1008;
	wire signed [31:0] w_sys_tmp1009;
	wire signed [31:0] w_sys_tmp1010;
	wire        [31:0] w_sys_tmp1011;
	wire signed [31:0] w_sys_tmp1012;
	wire signed [31:0] w_sys_tmp1013;
	wire signed [31:0] w_sys_tmp1015;
	wire signed [31:0] w_sys_tmp1016;
	wire signed [31:0] w_sys_tmp1089;
	wire               w_sys_tmp1090;
	wire               w_sys_tmp1091;
	wire signed [31:0] w_sys_tmp1092;
	wire signed [31:0] w_sys_tmp1093;
	wire               w_sys_tmp1094;
	wire               w_sys_tmp1095;
	wire signed [31:0] w_sys_tmp1096;
	wire signed [31:0] w_sys_tmp1099;
	wire signed [31:0] w_sys_tmp1100;
	wire signed [31:0] w_sys_tmp1101;
	wire        [31:0] w_sys_tmp1102;
	wire signed [31:0] w_sys_tmp1103;
	wire signed [31:0] w_sys_tmp1104;
	wire signed [31:0] w_sys_tmp1106;
	wire signed [31:0] w_sys_tmp1107;
	wire signed [31:0] w_sys_tmp1168;
	wire               w_sys_tmp1169;
	wire               w_sys_tmp1170;
	wire signed [31:0] w_sys_tmp1171;
	wire signed [31:0] w_sys_tmp1173;
	wire signed [31:0] w_sys_tmp1174;
	wire signed [31:0] w_sys_tmp1176;
	wire signed [31:0] w_sys_tmp1177;
	wire signed [31:0] w_sys_tmp1178;
	wire        [31:0] w_sys_tmp1179;
	wire signed [31:0] w_sys_tmp1180;
	wire signed [31:0] w_sys_tmp1181;
	wire signed [31:0] w_sys_tmp1183;
	wire signed [31:0] w_sys_tmp1184;
	wire signed [31:0] w_sys_tmp1257;
	wire               w_sys_tmp1258;
	wire               w_sys_tmp1259;
	wire signed [31:0] w_sys_tmp1260;
	wire signed [31:0] w_sys_tmp1262;
	wire signed [31:0] w_sys_tmp1263;
	wire signed [31:0] w_sys_tmp1265;
	wire signed [31:0] w_sys_tmp1266;
	wire signed [31:0] w_sys_tmp1267;
	wire        [31:0] w_sys_tmp1268;
	wire signed [31:0] w_sys_tmp1269;
	wire signed [31:0] w_sys_tmp1270;
	wire signed [31:0] w_sys_tmp1272;
	wire signed [31:0] w_sys_tmp1273;
	wire signed [31:0] w_sys_tmp1346;
	wire               w_sys_tmp1347;
	wire               w_sys_tmp1348;
	wire signed [31:0] w_sys_tmp1349;
	wire signed [31:0] w_sys_tmp1351;
	wire signed [31:0] w_sys_tmp1352;
	wire signed [31:0] w_sys_tmp1354;
	wire signed [31:0] w_sys_tmp1355;
	wire signed [31:0] w_sys_tmp1356;
	wire        [31:0] w_sys_tmp1357;
	wire signed [31:0] w_sys_tmp1358;
	wire signed [31:0] w_sys_tmp1359;
	wire signed [31:0] w_sys_tmp1361;
	wire signed [31:0] w_sys_tmp1362;
	wire               w_sys_tmp1435;
	wire               w_sys_tmp1436;
	wire signed [31:0] w_sys_tmp1437;
	wire signed [31:0] w_sys_tmp1438;
	wire               w_sys_tmp1439;
	wire               w_sys_tmp1440;
	wire signed [31:0] w_sys_tmp1441;
	wire signed [31:0] w_sys_tmp1444;
	wire signed [31:0] w_sys_tmp1445;
	wire        [31:0] w_sys_tmp1446;
	wire signed [31:0] w_sys_tmp1447;
	wire signed [31:0] w_sys_tmp1448;
	wire signed [31:0] w_sys_tmp1450;
	wire signed [31:0] w_sys_tmp1451;
	wire        [31:0] w_sys_tmp1452;
	wire signed [31:0] w_sys_tmp1453;
	wire signed [31:0] w_sys_tmp1454;
	wire signed [31:0] w_sys_tmp1456;
	wire signed [31:0] w_sys_tmp1457;
	wire        [31:0] w_sys_tmp1474;
	wire signed [31:0] w_sys_tmp1477;
	wire signed [31:0] w_sys_tmp1478;
	wire               w_sys_tmp1479;
	wire               w_sys_tmp1480;
	wire signed [31:0] w_sys_tmp1481;
	wire signed [31:0] w_sys_tmp1484;
	wire signed [31:0] w_sys_tmp1485;
	wire        [31:0] w_sys_tmp1486;
	wire signed [31:0] w_sys_tmp1487;
	wire signed [31:0] w_sys_tmp1488;
	wire signed [31:0] w_sys_tmp1490;
	wire signed [31:0] w_sys_tmp1491;
	wire        [31:0] w_sys_tmp1492;
	wire signed [31:0] w_sys_tmp1493;
	wire signed [31:0] w_sys_tmp1494;
	wire signed [31:0] w_sys_tmp1496;
	wire signed [31:0] w_sys_tmp1497;
	wire        [31:0] w_sys_tmp1514;
	wire signed [31:0] w_sys_tmp1517;
	wire signed [31:0] w_sys_tmp1518;
	wire               w_sys_tmp1519;
	wire               w_sys_tmp1520;
	wire signed [31:0] w_sys_tmp1521;
	wire signed [31:0] w_sys_tmp1524;
	wire signed [31:0] w_sys_tmp1525;
	wire        [31:0] w_sys_tmp1526;
	wire signed [31:0] w_sys_tmp1527;
	wire signed [31:0] w_sys_tmp1528;
	wire signed [31:0] w_sys_tmp1530;
	wire signed [31:0] w_sys_tmp1531;
	wire        [31:0] w_sys_tmp1532;
	wire signed [31:0] w_sys_tmp1533;
	wire signed [31:0] w_sys_tmp1534;
	wire signed [31:0] w_sys_tmp1536;
	wire signed [31:0] w_sys_tmp1537;
	wire        [31:0] w_sys_tmp1554;
	wire signed [31:0] w_sys_tmp1557;
	wire signed [31:0] w_sys_tmp1558;
	wire               w_sys_tmp1559;
	wire               w_sys_tmp1560;
	wire signed [31:0] w_sys_tmp1561;
	wire signed [31:0] w_sys_tmp1564;
	wire signed [31:0] w_sys_tmp1565;
	wire        [31:0] w_sys_tmp1566;
	wire signed [31:0] w_sys_tmp1567;
	wire signed [31:0] w_sys_tmp1568;
	wire signed [31:0] w_sys_tmp1570;
	wire signed [31:0] w_sys_tmp1571;
	wire        [31:0] w_sys_tmp1572;
	wire signed [31:0] w_sys_tmp1573;
	wire signed [31:0] w_sys_tmp1574;
	wire signed [31:0] w_sys_tmp1576;
	wire signed [31:0] w_sys_tmp1577;
	wire        [31:0] w_sys_tmp1594;
	wire signed [31:0] w_sys_tmp1595;
	wire signed [31:0] w_sys_tmp1596;
	wire signed [31:0] w_sys_tmp1597;
	wire signed [31:0] w_sys_tmp1598;
	wire               w_sys_tmp1599;
	wire               w_sys_tmp1600;
	wire signed [31:0] w_sys_tmp1601;
	wire signed [31:0] w_sys_tmp1604;
	wire signed [31:0] w_sys_tmp1605;
	wire signed [31:0] w_sys_tmp1606;
	wire signed [31:0] w_sys_tmp1607;
	wire        [31:0] w_sys_tmp1608;
	wire signed [31:0] w_sys_tmp1609;
	wire signed [31:0] w_sys_tmp1610;
	wire signed [31:0] w_sys_tmp1614;
	wire signed [31:0] w_sys_tmp1615;
	wire signed [31:0] w_sys_tmp1617;
	wire        [31:0] w_sys_tmp1618;
	wire signed [31:0] w_sys_tmp1619;
	wire signed [31:0] w_sys_tmp1620;
	wire signed [31:0] w_sys_tmp1624;
	wire signed [31:0] w_sys_tmp1625;
	wire signed [31:0] w_sys_tmp1627;
	wire signed [31:0] w_sys_tmp1628;
	wire signed [31:0] w_sys_tmp1629;
	wire signed [31:0] w_sys_tmp1633;
	wire signed [31:0] w_sys_tmp1634;
	wire signed [31:0] w_sys_tmp1636;
	wire signed [31:0] w_sys_tmp1638;
	wire signed [31:0] w_sys_tmp1639;
	wire signed [31:0] w_sys_tmp1643;
	wire signed [31:0] w_sys_tmp1644;
	wire signed [31:0] w_sys_tmp1646;
	wire signed [31:0] w_sys_tmp1647;
	wire signed [31:0] w_sys_tmp1648;
	wire signed [31:0] w_sys_tmp1652;
	wire signed [31:0] w_sys_tmp1653;
	wire signed [31:0] w_sys_tmp1655;
	wire        [31:0] w_sys_tmp1656;
	wire signed [31:0] w_sys_tmp1657;
	wire signed [31:0] w_sys_tmp1658;
	wire signed [31:0] w_sys_tmp1661;
	wire signed [31:0] w_sys_tmp1662;
	wire signed [31:0] w_sys_tmp1663;
	wire signed [31:0] w_sys_tmp1664;
	wire signed [31:0] w_sys_tmp1665;
	wire signed [31:0] w_sys_tmp1666;
	wire signed [31:0] w_sys_tmp1667;
	wire signed [31:0] w_sys_tmp1668;
	wire signed [31:0] w_sys_tmp1669;
	wire signed [31:0] w_sys_tmp1670;
	wire signed [31:0] w_sys_tmp1671;
	wire signed [31:0] w_sys_tmp1672;
	wire signed [31:0] w_sys_tmp2099;
	wire               w_sys_tmp2100;
	wire               w_sys_tmp2101;
	wire signed [31:0] w_sys_tmp2102;
	wire signed [31:0] w_sys_tmp2104;
	wire signed [31:0] w_sys_tmp2105;
	wire signed [31:0] w_sys_tmp2107;
	wire signed [31:0] w_sys_tmp2108;
	wire signed [31:0] w_sys_tmp2109;
	wire signed [31:0] w_sys_tmp2110;
	wire        [31:0] w_sys_tmp2111;
	wire signed [31:0] w_sys_tmp2112;
	wire signed [31:0] w_sys_tmp2113;
	wire signed [31:0] w_sys_tmp2114;
	wire signed [31:0] w_sys_tmp2118;
	wire signed [31:0] w_sys_tmp2121;
	wire        [31:0] w_sys_tmp2122;
	wire signed [31:0] w_sys_tmp2128;
	wire signed [31:0] w_sys_tmp2131;
	wire signed [31:0] w_sys_tmp2132;
	wire signed [31:0] w_sys_tmp2138;
	wire signed [31:0] w_sys_tmp2141;
	wire signed [31:0] w_sys_tmp2148;
	wire signed [31:0] w_sys_tmp2151;
	wire signed [31:0] w_sys_tmp2152;
	wire signed [31:0] w_sys_tmp2158;
	wire signed [31:0] w_sys_tmp2161;
	wire        [31:0] w_sys_tmp2162;
	wire signed [31:0] w_sys_tmp2167;
	wire signed [31:0] w_sys_tmp2546;
	wire               w_sys_tmp2547;
	wire               w_sys_tmp2548;
	wire signed [31:0] w_sys_tmp2549;
	wire signed [31:0] w_sys_tmp2551;
	wire signed [31:0] w_sys_tmp2552;
	wire signed [31:0] w_sys_tmp2554;
	wire signed [31:0] w_sys_tmp2555;
	wire signed [31:0] w_sys_tmp2556;
	wire signed [31:0] w_sys_tmp2557;
	wire        [31:0] w_sys_tmp2558;
	wire signed [31:0] w_sys_tmp2559;
	wire signed [31:0] w_sys_tmp2560;
	wire signed [31:0] w_sys_tmp2561;
	wire signed [31:0] w_sys_tmp2565;
	wire signed [31:0] w_sys_tmp2568;
	wire        [31:0] w_sys_tmp2569;
	wire signed [31:0] w_sys_tmp2575;
	wire signed [31:0] w_sys_tmp2578;
	wire signed [31:0] w_sys_tmp2579;
	wire signed [31:0] w_sys_tmp2585;
	wire signed [31:0] w_sys_tmp2588;
	wire signed [31:0] w_sys_tmp2595;
	wire signed [31:0] w_sys_tmp2598;
	wire signed [31:0] w_sys_tmp2599;
	wire signed [31:0] w_sys_tmp2605;
	wire signed [31:0] w_sys_tmp2608;
	wire        [31:0] w_sys_tmp2609;
	wire signed [31:0] w_sys_tmp2614;
	wire signed [31:0] w_sys_tmp2993;
	wire               w_sys_tmp2994;
	wire               w_sys_tmp2995;
	wire signed [31:0] w_sys_tmp2996;
	wire signed [31:0] w_sys_tmp2998;
	wire signed [31:0] w_sys_tmp2999;
	wire signed [31:0] w_sys_tmp3001;
	wire signed [31:0] w_sys_tmp3002;
	wire signed [31:0] w_sys_tmp3003;
	wire signed [31:0] w_sys_tmp3004;
	wire        [31:0] w_sys_tmp3005;
	wire signed [31:0] w_sys_tmp3006;
	wire signed [31:0] w_sys_tmp3007;
	wire signed [31:0] w_sys_tmp3008;
	wire signed [31:0] w_sys_tmp3012;
	wire signed [31:0] w_sys_tmp3015;
	wire        [31:0] w_sys_tmp3016;
	wire signed [31:0] w_sys_tmp3022;
	wire signed [31:0] w_sys_tmp3025;
	wire signed [31:0] w_sys_tmp3026;
	wire signed [31:0] w_sys_tmp3032;
	wire signed [31:0] w_sys_tmp3035;
	wire signed [31:0] w_sys_tmp3042;
	wire signed [31:0] w_sys_tmp3045;
	wire signed [31:0] w_sys_tmp3046;
	wire signed [31:0] w_sys_tmp3052;
	wire signed [31:0] w_sys_tmp3055;
	wire        [31:0] w_sys_tmp3056;
	wire signed [31:0] w_sys_tmp3061;
	wire signed [31:0] w_sys_tmp3440;
	wire               w_sys_tmp3441;
	wire               w_sys_tmp3442;
	wire signed [31:0] w_sys_tmp3443;
	wire signed [31:0] w_sys_tmp3444;
	wire signed [31:0] w_sys_tmp3445;
	wire               w_sys_tmp3446;
	wire               w_sys_tmp3447;
	wire signed [31:0] w_sys_tmp3448;
	wire signed [31:0] w_sys_tmp3451;
	wire signed [31:0] w_sys_tmp3452;
	wire signed [31:0] w_sys_tmp3453;
	wire        [31:0] w_sys_tmp3454;
	wire signed [31:0] w_sys_tmp3455;
	wire signed [31:0] w_sys_tmp3456;
	wire signed [31:0] w_sys_tmp3458;
	wire signed [31:0] w_sys_tmp3459;
	wire signed [31:0] w_sys_tmp3520;
	wire               w_sys_tmp3521;
	wire               w_sys_tmp3522;
	wire signed [31:0] w_sys_tmp3523;
	wire signed [31:0] w_sys_tmp3525;
	wire signed [31:0] w_sys_tmp3526;
	wire signed [31:0] w_sys_tmp3528;
	wire signed [31:0] w_sys_tmp3529;
	wire signed [31:0] w_sys_tmp3530;
	wire        [31:0] w_sys_tmp3531;
	wire signed [31:0] w_sys_tmp3532;
	wire signed [31:0] w_sys_tmp3533;
	wire signed [31:0] w_sys_tmp3535;
	wire signed [31:0] w_sys_tmp3536;
	wire signed [31:0] w_sys_tmp3537;
	wire signed [31:0] w_sys_tmp3616;
	wire               w_sys_tmp3617;
	wire               w_sys_tmp3618;
	wire signed [31:0] w_sys_tmp3619;
	wire signed [31:0] w_sys_tmp3621;
	wire signed [31:0] w_sys_tmp3622;
	wire signed [31:0] w_sys_tmp3624;
	wire signed [31:0] w_sys_tmp3625;
	wire signed [31:0] w_sys_tmp3626;
	wire        [31:0] w_sys_tmp3627;
	wire signed [31:0] w_sys_tmp3628;
	wire signed [31:0] w_sys_tmp3629;
	wire signed [31:0] w_sys_tmp3631;
	wire signed [31:0] w_sys_tmp3632;
	wire signed [31:0] w_sys_tmp3633;
	wire signed [31:0] w_sys_tmp3712;
	wire               w_sys_tmp3713;
	wire               w_sys_tmp3714;
	wire signed [31:0] w_sys_tmp3715;
	wire signed [31:0] w_sys_tmp3717;
	wire signed [31:0] w_sys_tmp3718;
	wire signed [31:0] w_sys_tmp3720;
	wire signed [31:0] w_sys_tmp3721;
	wire signed [31:0] w_sys_tmp3722;
	wire        [31:0] w_sys_tmp3723;
	wire signed [31:0] w_sys_tmp3724;
	wire signed [31:0] w_sys_tmp3725;
	wire signed [31:0] w_sys_tmp3727;
	wire signed [31:0] w_sys_tmp3728;
	wire signed [31:0] w_sys_tmp3729;
	wire signed [31:0] w_sys_tmp3808;
	wire               w_sys_tmp3809;
	wire               w_sys_tmp3810;
	wire signed [31:0] w_sys_tmp3811;
	wire signed [31:0] w_sys_tmp3812;
	wire signed [31:0] w_sys_tmp3813;
	wire               w_sys_tmp3814;
	wire               w_sys_tmp3815;
	wire signed [31:0] w_sys_tmp3816;
	wire signed [31:0] w_sys_tmp3819;
	wire signed [31:0] w_sys_tmp3820;
	wire signed [31:0] w_sys_tmp3821;
	wire        [31:0] w_sys_tmp3822;
	wire signed [31:0] w_sys_tmp3823;
	wire signed [31:0] w_sys_tmp3824;
	wire signed [31:0] w_sys_tmp3826;
	wire signed [31:0] w_sys_tmp3827;
	wire signed [31:0] w_sys_tmp3888;
	wire               w_sys_tmp3889;
	wire               w_sys_tmp3890;
	wire signed [31:0] w_sys_tmp3891;
	wire signed [31:0] w_sys_tmp3893;
	wire signed [31:0] w_sys_tmp3894;
	wire signed [31:0] w_sys_tmp3896;
	wire signed [31:0] w_sys_tmp3897;
	wire signed [31:0] w_sys_tmp3898;
	wire        [31:0] w_sys_tmp3899;
	wire signed [31:0] w_sys_tmp3900;
	wire signed [31:0] w_sys_tmp3901;
	wire signed [31:0] w_sys_tmp3903;
	wire signed [31:0] w_sys_tmp3904;
	wire signed [31:0] w_sys_tmp3905;
	wire signed [31:0] w_sys_tmp3984;
	wire               w_sys_tmp3985;
	wire               w_sys_tmp3986;
	wire signed [31:0] w_sys_tmp3987;
	wire signed [31:0] w_sys_tmp3989;
	wire signed [31:0] w_sys_tmp3990;
	wire signed [31:0] w_sys_tmp3992;
	wire signed [31:0] w_sys_tmp3993;
	wire signed [31:0] w_sys_tmp3994;
	wire        [31:0] w_sys_tmp3995;
	wire signed [31:0] w_sys_tmp3996;
	wire signed [31:0] w_sys_tmp3997;
	wire signed [31:0] w_sys_tmp3999;
	wire signed [31:0] w_sys_tmp4000;
	wire signed [31:0] w_sys_tmp4001;
	wire signed [31:0] w_sys_tmp4080;
	wire               w_sys_tmp4081;
	wire               w_sys_tmp4082;
	wire signed [31:0] w_sys_tmp4083;
	wire signed [31:0] w_sys_tmp4085;
	wire signed [31:0] w_sys_tmp4086;
	wire signed [31:0] w_sys_tmp4088;
	wire signed [31:0] w_sys_tmp4089;
	wire signed [31:0] w_sys_tmp4090;
	wire        [31:0] w_sys_tmp4091;
	wire signed [31:0] w_sys_tmp4092;
	wire signed [31:0] w_sys_tmp4093;
	wire signed [31:0] w_sys_tmp4095;
	wire signed [31:0] w_sys_tmp4096;
	wire signed [31:0] w_sys_tmp4097;
	wire signed [31:0] w_sys_tmp4176;
	wire               w_sys_tmp4177;
	wire               w_sys_tmp4178;
	wire signed [31:0] w_sys_tmp4179;
	wire signed [31:0] w_sys_tmp4180;
	wire signed [31:0] w_sys_tmp4181;
	wire               w_sys_tmp4182;
	wire               w_sys_tmp4183;
	wire signed [31:0] w_sys_tmp4184;
	wire signed [31:0] w_sys_tmp4187;
	wire signed [31:0] w_sys_tmp4188;
	wire signed [31:0] w_sys_tmp4189;
	wire        [31:0] w_sys_tmp4190;
	wire signed [31:0] w_sys_tmp4191;
	wire signed [31:0] w_sys_tmp4192;
	wire signed [31:0] w_sys_tmp4194;
	wire signed [31:0] w_sys_tmp4195;
	wire signed [31:0] w_sys_tmp4256;
	wire               w_sys_tmp4257;
	wire               w_sys_tmp4258;
	wire signed [31:0] w_sys_tmp4259;
	wire signed [31:0] w_sys_tmp4261;
	wire signed [31:0] w_sys_tmp4262;
	wire signed [31:0] w_sys_tmp4264;
	wire signed [31:0] w_sys_tmp4265;
	wire signed [31:0] w_sys_tmp4266;
	wire        [31:0] w_sys_tmp4267;
	wire signed [31:0] w_sys_tmp4268;
	wire signed [31:0] w_sys_tmp4269;
	wire signed [31:0] w_sys_tmp4271;
	wire signed [31:0] w_sys_tmp4272;
	wire signed [31:0] w_sys_tmp4273;
	wire signed [31:0] w_sys_tmp4352;
	wire               w_sys_tmp4353;
	wire               w_sys_tmp4354;
	wire signed [31:0] w_sys_tmp4355;
	wire signed [31:0] w_sys_tmp4357;
	wire signed [31:0] w_sys_tmp4358;
	wire signed [31:0] w_sys_tmp4360;
	wire signed [31:0] w_sys_tmp4361;
	wire signed [31:0] w_sys_tmp4362;
	wire        [31:0] w_sys_tmp4363;
	wire signed [31:0] w_sys_tmp4364;
	wire signed [31:0] w_sys_tmp4365;
	wire signed [31:0] w_sys_tmp4367;
	wire signed [31:0] w_sys_tmp4368;
	wire signed [31:0] w_sys_tmp4369;
	wire signed [31:0] w_sys_tmp4448;
	wire               w_sys_tmp4449;
	wire               w_sys_tmp4450;
	wire signed [31:0] w_sys_tmp4451;
	wire signed [31:0] w_sys_tmp4453;
	wire signed [31:0] w_sys_tmp4454;
	wire signed [31:0] w_sys_tmp4456;
	wire signed [31:0] w_sys_tmp4457;
	wire signed [31:0] w_sys_tmp4458;
	wire        [31:0] w_sys_tmp4459;
	wire signed [31:0] w_sys_tmp4460;
	wire signed [31:0] w_sys_tmp4461;
	wire signed [31:0] w_sys_tmp4463;
	wire signed [31:0] w_sys_tmp4464;
	wire signed [31:0] w_sys_tmp4465;
	wire signed [31:0] w_sys_tmp4544;
	wire               w_sys_tmp4545;
	wire               w_sys_tmp4546;
	wire signed [31:0] w_sys_tmp4547;
	wire signed [31:0] w_sys_tmp4548;
	wire signed [31:0] w_sys_tmp4549;
	wire               w_sys_tmp4550;
	wire               w_sys_tmp4551;
	wire signed [31:0] w_sys_tmp4552;
	wire signed [31:0] w_sys_tmp4555;
	wire signed [31:0] w_sys_tmp4556;
	wire signed [31:0] w_sys_tmp4557;
	wire        [31:0] w_sys_tmp4558;
	wire signed [31:0] w_sys_tmp4559;
	wire signed [31:0] w_sys_tmp4560;
	wire signed [31:0] w_sys_tmp4562;
	wire signed [31:0] w_sys_tmp4563;
	wire signed [31:0] w_sys_tmp4624;
	wire               w_sys_tmp4625;
	wire               w_sys_tmp4626;
	wire signed [31:0] w_sys_tmp4627;
	wire signed [31:0] w_sys_tmp4629;
	wire signed [31:0] w_sys_tmp4630;
	wire signed [31:0] w_sys_tmp4632;
	wire signed [31:0] w_sys_tmp4633;
	wire signed [31:0] w_sys_tmp4634;
	wire        [31:0] w_sys_tmp4635;
	wire signed [31:0] w_sys_tmp4636;
	wire signed [31:0] w_sys_tmp4637;
	wire signed [31:0] w_sys_tmp4639;
	wire signed [31:0] w_sys_tmp4640;
	wire signed [31:0] w_sys_tmp4641;
	wire signed [31:0] w_sys_tmp4720;
	wire               w_sys_tmp4721;
	wire               w_sys_tmp4722;
	wire signed [31:0] w_sys_tmp4723;
	wire signed [31:0] w_sys_tmp4725;
	wire signed [31:0] w_sys_tmp4726;
	wire signed [31:0] w_sys_tmp4728;
	wire signed [31:0] w_sys_tmp4729;
	wire signed [31:0] w_sys_tmp4730;
	wire        [31:0] w_sys_tmp4731;
	wire signed [31:0] w_sys_tmp4732;
	wire signed [31:0] w_sys_tmp4733;
	wire signed [31:0] w_sys_tmp4735;
	wire signed [31:0] w_sys_tmp4736;
	wire signed [31:0] w_sys_tmp4737;
	wire signed [31:0] w_sys_tmp4816;
	wire               w_sys_tmp4817;
	wire               w_sys_tmp4818;
	wire signed [31:0] w_sys_tmp4819;
	wire signed [31:0] w_sys_tmp4821;
	wire signed [31:0] w_sys_tmp4822;
	wire signed [31:0] w_sys_tmp4824;
	wire signed [31:0] w_sys_tmp4825;
	wire signed [31:0] w_sys_tmp4826;
	wire        [31:0] w_sys_tmp4827;
	wire signed [31:0] w_sys_tmp4828;
	wire signed [31:0] w_sys_tmp4829;
	wire signed [31:0] w_sys_tmp4831;
	wire signed [31:0] w_sys_tmp4832;
	wire signed [31:0] w_sys_tmp4833;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 5'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 7'h1);
	assign w_fld_u_0_addr_0 = 15'sh0;
	assign w_fld_u_0_datain_0 = 32'h0;
	assign w_fld_u_0_r_w_0 = 1'h0;
	assign w_fld_u_0_ce_0 = w_sys_ce;
	assign w_fld_u_0_ce_1 = w_sys_ce;
	assign w_sub09_u_addr = ( (|r_sys_processing_methodID) ? r_sub09_u_addr : 13'sh0 ) ;
	assign w_sub09_u_datain = ( (|r_sys_processing_methodID) ? r_sub09_u_datain : 32'h0 ) ;
	assign w_sub09_u_r_w = ( (|r_sys_processing_methodID) ? r_sub09_u_r_w : 1'h0 ) ;
	assign w_sub09_result_addr = ( (|r_sys_processing_methodID) ? r_sub09_result_addr : 13'sh0 ) ;
	assign w_sub09_result_datain = ( (|r_sys_processing_methodID) ? r_sub09_result_datain : 32'h0 ) ;
	assign w_sub09_result_r_w = ( (|r_sys_processing_methodID) ? r_sub09_result_r_w : 1'h0 ) ;
	assign w_sub08_u_addr = ( (|r_sys_processing_methodID) ? r_sub08_u_addr : 13'sh0 ) ;
	assign w_sub08_u_datain = ( (|r_sys_processing_methodID) ? r_sub08_u_datain : 32'h0 ) ;
	assign w_sub08_u_r_w = ( (|r_sys_processing_methodID) ? r_sub08_u_r_w : 1'h0 ) ;
	assign w_sub08_result_addr = ( (|r_sys_processing_methodID) ? r_sub08_result_addr : 13'sh0 ) ;
	assign w_sub08_result_datain = ( (|r_sys_processing_methodID) ? r_sub08_result_datain : 32'h0 ) ;
	assign w_sub08_result_r_w = ( (|r_sys_processing_methodID) ? r_sub08_result_r_w : 1'h0 ) ;
	assign w_sub12_u_addr = ( (|r_sys_processing_methodID) ? r_sub12_u_addr : 13'sh0 ) ;
	assign w_sub12_u_datain = ( (|r_sys_processing_methodID) ? r_sub12_u_datain : 32'h0 ) ;
	assign w_sub12_u_r_w = ( (|r_sys_processing_methodID) ? r_sub12_u_r_w : 1'h0 ) ;
	assign w_sub12_result_addr = ( (|r_sys_processing_methodID) ? r_sub12_result_addr : 13'sh0 ) ;
	assign w_sub12_result_datain = ( (|r_sys_processing_methodID) ? r_sub12_result_datain : 32'h0 ) ;
	assign w_sub12_result_r_w = ( (|r_sys_processing_methodID) ? r_sub12_result_r_w : 1'h0 ) ;
	assign w_sub03_u_addr = ( (|r_sys_processing_methodID) ? r_sub03_u_addr : 13'sh0 ) ;
	assign w_sub03_u_datain = ( (|r_sys_processing_methodID) ? r_sub03_u_datain : 32'h0 ) ;
	assign w_sub03_u_r_w = ( (|r_sys_processing_methodID) ? r_sub03_u_r_w : 1'h0 ) ;
	assign w_sub03_result_addr = ( (|r_sys_processing_methodID) ? r_sub03_result_addr : 13'sh0 ) ;
	assign w_sub03_result_datain = ( (|r_sys_processing_methodID) ? r_sub03_result_datain : 32'h0 ) ;
	assign w_sub03_result_r_w = ( (|r_sys_processing_methodID) ? r_sub03_result_r_w : 1'h0 ) ;
	assign w_sub02_u_addr = ( (|r_sys_processing_methodID) ? r_sub02_u_addr : 13'sh0 ) ;
	assign w_sub02_u_datain = ( (|r_sys_processing_methodID) ? r_sub02_u_datain : 32'h0 ) ;
	assign w_sub02_u_r_w = ( (|r_sys_processing_methodID) ? r_sub02_u_r_w : 1'h0 ) ;
	assign w_sub02_result_addr = ( (|r_sys_processing_methodID) ? r_sub02_result_addr : 13'sh0 ) ;
	assign w_sub02_result_datain = ( (|r_sys_processing_methodID) ? r_sub02_result_datain : 32'h0 ) ;
	assign w_sub02_result_r_w = ( (|r_sys_processing_methodID) ? r_sub02_result_r_w : 1'h0 ) ;
	assign w_sub11_u_addr = ( (|r_sys_processing_methodID) ? r_sub11_u_addr : 13'sh0 ) ;
	assign w_sub11_u_datain = ( (|r_sys_processing_methodID) ? r_sub11_u_datain : 32'h0 ) ;
	assign w_sub11_u_r_w = ( (|r_sys_processing_methodID) ? r_sub11_u_r_w : 1'h0 ) ;
	assign w_sub11_result_addr = ( (|r_sys_processing_methodID) ? r_sub11_result_addr : 13'sh0 ) ;
	assign w_sub11_result_datain = ( (|r_sys_processing_methodID) ? r_sub11_result_datain : 32'h0 ) ;
	assign w_sub11_result_r_w = ( (|r_sys_processing_methodID) ? r_sub11_result_r_w : 1'h0 ) ;
	assign w_sub14_u_addr = ( (|r_sys_processing_methodID) ? r_sub14_u_addr : 13'sh0 ) ;
	assign w_sub14_u_datain = ( (|r_sys_processing_methodID) ? r_sub14_u_datain : 32'h0 ) ;
	assign w_sub14_u_r_w = ( (|r_sys_processing_methodID) ? r_sub14_u_r_w : 1'h0 ) ;
	assign w_sub14_result_addr = ( (|r_sys_processing_methodID) ? r_sub14_result_addr : 13'sh0 ) ;
	assign w_sub14_result_datain = ( (|r_sys_processing_methodID) ? r_sub14_result_datain : 32'h0 ) ;
	assign w_sub14_result_r_w = ( (|r_sys_processing_methodID) ? r_sub14_result_r_w : 1'h0 ) ;
	assign w_sub01_u_addr = ( (|r_sys_processing_methodID) ? r_sub01_u_addr : 13'sh0 ) ;
	assign w_sub01_u_datain = ( (|r_sys_processing_methodID) ? r_sub01_u_datain : 32'h0 ) ;
	assign w_sub01_u_r_w = ( (|r_sys_processing_methodID) ? r_sub01_u_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 13'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub13_u_addr = ( (|r_sys_processing_methodID) ? r_sub13_u_addr : 13'sh0 ) ;
	assign w_sub13_u_datain = ( (|r_sys_processing_methodID) ? r_sub13_u_datain : 32'h0 ) ;
	assign w_sub13_u_r_w = ( (|r_sys_processing_methodID) ? r_sub13_u_r_w : 1'h0 ) ;
	assign w_sub13_result_addr = ( (|r_sys_processing_methodID) ? r_sub13_result_addr : 13'sh0 ) ;
	assign w_sub13_result_datain = ( (|r_sys_processing_methodID) ? r_sub13_result_datain : 32'h0 ) ;
	assign w_sub13_result_r_w = ( (|r_sys_processing_methodID) ? r_sub13_result_r_w : 1'h0 ) ;
	assign w_sub00_u_addr = ( (|r_sys_processing_methodID) ? r_sub00_u_addr : 13'sh0 ) ;
	assign w_sub00_u_datain = ( (|r_sys_processing_methodID) ? r_sub00_u_datain : 32'h0 ) ;
	assign w_sub00_u_r_w = ( (|r_sys_processing_methodID) ? r_sub00_u_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 13'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sub07_u_addr = ( (|r_sys_processing_methodID) ? r_sub07_u_addr : 13'sh0 ) ;
	assign w_sub07_u_datain = ( (|r_sys_processing_methodID) ? r_sub07_u_datain : 32'h0 ) ;
	assign w_sub07_u_r_w = ( (|r_sys_processing_methodID) ? r_sub07_u_r_w : 1'h0 ) ;
	assign w_sub07_result_addr = ( (|r_sys_processing_methodID) ? r_sub07_result_addr : 13'sh0 ) ;
	assign w_sub07_result_datain = ( (|r_sys_processing_methodID) ? r_sub07_result_datain : 32'h0 ) ;
	assign w_sub07_result_r_w = ( (|r_sys_processing_methodID) ? r_sub07_result_r_w : 1'h0 ) ;
	assign w_sub06_u_addr = ( (|r_sys_processing_methodID) ? r_sub06_u_addr : 13'sh0 ) ;
	assign w_sub06_u_datain = ( (|r_sys_processing_methodID) ? r_sub06_u_datain : 32'h0 ) ;
	assign w_sub06_u_r_w = ( (|r_sys_processing_methodID) ? r_sub06_u_r_w : 1'h0 ) ;
	assign w_sub06_result_addr = ( (|r_sys_processing_methodID) ? r_sub06_result_addr : 13'sh0 ) ;
	assign w_sub06_result_datain = ( (|r_sys_processing_methodID) ? r_sub06_result_datain : 32'h0 ) ;
	assign w_sub06_result_r_w = ( (|r_sys_processing_methodID) ? r_sub06_result_r_w : 1'h0 ) ;
	assign w_sub15_u_addr = ( (|r_sys_processing_methodID) ? r_sub15_u_addr : 13'sh0 ) ;
	assign w_sub15_u_datain = ( (|r_sys_processing_methodID) ? r_sub15_u_datain : 32'h0 ) ;
	assign w_sub15_u_r_w = ( (|r_sys_processing_methodID) ? r_sub15_u_r_w : 1'h0 ) ;
	assign w_sub15_result_addr = ( (|r_sys_processing_methodID) ? r_sub15_result_addr : 13'sh0 ) ;
	assign w_sub15_result_datain = ( (|r_sys_processing_methodID) ? r_sub15_result_datain : 32'h0 ) ;
	assign w_sub15_result_r_w = ( (|r_sys_processing_methodID) ? r_sub15_result_r_w : 1'h0 ) ;
	assign w_sub05_u_addr = ( (|r_sys_processing_methodID) ? r_sub05_u_addr : 13'sh0 ) ;
	assign w_sub05_u_datain = ( (|r_sys_processing_methodID) ? r_sub05_u_datain : 32'h0 ) ;
	assign w_sub05_u_r_w = ( (|r_sys_processing_methodID) ? r_sub05_u_r_w : 1'h0 ) ;
	assign w_sub05_result_addr = ( (|r_sys_processing_methodID) ? r_sub05_result_addr : 13'sh0 ) ;
	assign w_sub05_result_datain = ( (|r_sys_processing_methodID) ? r_sub05_result_datain : 32'h0 ) ;
	assign w_sub05_result_r_w = ( (|r_sys_processing_methodID) ? r_sub05_result_r_w : 1'h0 ) ;
	assign w_sub04_u_addr = ( (|r_sys_processing_methodID) ? r_sub04_u_addr : 13'sh0 ) ;
	assign w_sub04_u_datain = ( (|r_sys_processing_methodID) ? r_sub04_u_datain : 32'h0 ) ;
	assign w_sub04_u_r_w = ( (|r_sys_processing_methodID) ? r_sub04_u_r_w : 1'h0 ) ;
	assign w_sub04_result_addr = ( (|r_sys_processing_methodID) ? r_sub04_result_addr : 13'sh0 ) ;
	assign w_sub04_result_datain = ( (|r_sys_processing_methodID) ? r_sub04_result_datain : 32'h0 ) ;
	assign w_sub04_result_r_w = ( (|r_sys_processing_methodID) ? r_sub04_result_r_w : 1'h0 ) ;
	assign w_sub10_u_addr = ( (|r_sys_processing_methodID) ? r_sub10_u_addr : 13'sh0 ) ;
	assign w_sub10_u_datain = ( (|r_sys_processing_methodID) ? r_sub10_u_datain : 32'h0 ) ;
	assign w_sub10_u_r_w = ( (|r_sys_processing_methodID) ? r_sub10_u_r_w : 1'h0 ) ;
	assign w_sub10_result_addr = ( (|r_sys_processing_methodID) ? r_sub10_result_addr : 13'sh0 ) ;
	assign w_sub10_result_datain = ( (|r_sys_processing_methodID) ? r_sub10_result_datain : 32'h0 ) ;
	assign w_sub10_result_r_w = ( (|r_sys_processing_methodID) ? r_sub10_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh00000081;
	assign w_sys_tmp3 = 32'sh00000190;
	assign w_sys_tmp4 = ( !w_sys_tmp5 );
	assign w_sys_tmp5 = (r_run_my_21 < r_run_k_17);
	assign w_sys_tmp6 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp7 = ( !w_sys_tmp8 );
	assign w_sys_tmp8 = (r_run_mx_20 < r_run_j_18);
	assign w_sys_tmp11 = (w_sys_tmp12 + r_run_k_17);
	assign w_sys_tmp12 = (r_run_j_18 * w_sys_tmp13);
	assign w_sys_tmp13 = 32'sh00000081;
	assign w_sys_tmp14 = 32'h0;
	assign w_sys_tmp15 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp52 = ( !w_sys_tmp53 );
	assign w_sys_tmp53 = (w_sys_tmp54 < r_run_k_17);
	assign w_sys_tmp54 = 32'sh00000021;
	assign w_sys_tmp55 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp56 = ( !w_sys_tmp57 );
	assign w_sys_tmp57 = (w_sys_tmp58 < r_run_j_18);
	assign w_sys_tmp58 = 32'sh00000021;
	assign w_sys_tmp61 = (w_sys_tmp62 + r_run_k_17);
	assign w_sys_tmp62 = (r_run_j_18 * w_sys_tmp63);
	assign w_sys_tmp63 = 32'sh00000081;
	assign w_sys_tmp64 = w_fld_u_0_dataout_1;
	assign w_sys_tmp65 = (w_sys_tmp66 + r_run_k_17);
	assign w_sys_tmp66 = (r_run_copy0_j_24 * w_sys_tmp63);
	assign w_sys_tmp68 = (r_run_copy0_j_24 + w_sys_intOne);
	assign w_sys_tmp69 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp130 = 32'sh00000020;
	assign w_sys_tmp131 = ( !w_sys_tmp132 );
	assign w_sys_tmp132 = (w_sys_tmp133 < r_run_j_18);
	assign w_sys_tmp133 = 32'sh00000041;
	assign w_sys_tmp135 = (r_run_j_18 - w_sys_tmp136);
	assign w_sys_tmp136 = 32'sh0000001f;
	assign w_sys_tmp138 = (w_sys_tmp139 + r_run_k_17);
	assign w_sys_tmp139 = (r_run_tmpj_23 * w_sys_tmp140);
	assign w_sys_tmp140 = 32'sh00000081;
	assign w_sys_tmp141 = w_fld_u_0_dataout_1;
	assign w_sys_tmp142 = (w_sys_tmp143 + r_run_k_17);
	assign w_sys_tmp143 = (r_run_copy0_j_25 * w_sys_tmp140);
	assign w_sys_tmp145 = (r_run_copy0_j_25 + w_sys_intOne);
	assign w_sys_tmp146 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp219 = 32'sh00000040;
	assign w_sys_tmp220 = ( !w_sys_tmp221 );
	assign w_sys_tmp221 = (w_sys_tmp222 < r_run_j_18);
	assign w_sys_tmp222 = 32'sh00000061;
	assign w_sys_tmp224 = (r_run_j_18 - w_sys_tmp225);
	assign w_sys_tmp225 = 32'sh0000003f;
	assign w_sys_tmp227 = (w_sys_tmp228 + r_run_k_17);
	assign w_sys_tmp228 = (r_run_tmpj_23 * w_sys_tmp229);
	assign w_sys_tmp229 = 32'sh00000081;
	assign w_sys_tmp230 = w_fld_u_0_dataout_1;
	assign w_sys_tmp231 = (w_sys_tmp232 + r_run_k_17);
	assign w_sys_tmp232 = (r_run_copy0_j_26 * w_sys_tmp229);
	assign w_sys_tmp234 = (r_run_copy0_j_26 + w_sys_intOne);
	assign w_sys_tmp235 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp308 = 32'sh00000060;
	assign w_sys_tmp309 = ( !w_sys_tmp310 );
	assign w_sys_tmp310 = (w_sys_tmp311 < r_run_j_18);
	assign w_sys_tmp311 = 32'sh00000081;
	assign w_sys_tmp313 = (r_run_j_18 - w_sys_tmp314);
	assign w_sys_tmp314 = 32'sh0000005f;
	assign w_sys_tmp316 = (w_sys_tmp317 + r_run_k_17);
	assign w_sys_tmp317 = (r_run_tmpj_23 * w_sys_tmp318);
	assign w_sys_tmp318 = 32'sh00000081;
	assign w_sys_tmp319 = w_fld_u_0_dataout_1;
	assign w_sys_tmp320 = (w_sys_tmp321 + r_run_k_17);
	assign w_sys_tmp321 = (r_run_copy0_j_27 * w_sys_tmp318);
	assign w_sys_tmp323 = (r_run_copy0_j_27 + w_sys_intOne);
	assign w_sys_tmp324 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp397 = 32'sh00000020;
	assign w_sys_tmp398 = ( !w_sys_tmp399 );
	assign w_sys_tmp399 = (w_sys_tmp400 < r_run_k_17);
	assign w_sys_tmp400 = 32'sh00000041;
	assign w_sys_tmp401 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp402 = ( !w_sys_tmp403 );
	assign w_sys_tmp403 = (w_sys_tmp404 < r_run_j_18);
	assign w_sys_tmp404 = 32'sh00000021;
	assign w_sys_tmp407 = (w_sys_tmp408 + r_run_k_17);
	assign w_sys_tmp408 = (r_run_j_18 * w_sys_tmp409);
	assign w_sys_tmp409 = 32'sh00000081;
	assign w_sys_tmp410 = w_fld_u_0_dataout_1;
	assign w_sys_tmp411 = (w_sys_tmp412 + r_run_k_17);
	assign w_sys_tmp412 = (r_run_copy0_j_28 * w_sys_tmp409);
	assign w_sys_tmp414 = (r_run_copy0_j_28 + w_sys_intOne);
	assign w_sys_tmp415 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp476 = 32'sh00000020;
	assign w_sys_tmp477 = ( !w_sys_tmp478 );
	assign w_sys_tmp478 = (w_sys_tmp479 < r_run_j_18);
	assign w_sys_tmp479 = 32'sh00000041;
	assign w_sys_tmp481 = (r_run_j_18 - w_sys_tmp482);
	assign w_sys_tmp482 = 32'sh0000001f;
	assign w_sys_tmp484 = (w_sys_tmp485 + r_run_k_17);
	assign w_sys_tmp485 = (r_run_tmpj_23 * w_sys_tmp486);
	assign w_sys_tmp486 = 32'sh00000081;
	assign w_sys_tmp487 = w_fld_u_0_dataout_1;
	assign w_sys_tmp488 = (w_sys_tmp489 + r_run_k_17);
	assign w_sys_tmp489 = (r_run_copy0_j_29 * w_sys_tmp486);
	assign w_sys_tmp491 = (r_run_copy0_j_29 + w_sys_intOne);
	assign w_sys_tmp492 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp565 = 32'sh00000040;
	assign w_sys_tmp566 = ( !w_sys_tmp567 );
	assign w_sys_tmp567 = (w_sys_tmp568 < r_run_j_18);
	assign w_sys_tmp568 = 32'sh00000061;
	assign w_sys_tmp570 = (r_run_j_18 - w_sys_tmp571);
	assign w_sys_tmp571 = 32'sh0000003f;
	assign w_sys_tmp573 = (w_sys_tmp574 + r_run_k_17);
	assign w_sys_tmp574 = (r_run_tmpj_23 * w_sys_tmp575);
	assign w_sys_tmp575 = 32'sh00000081;
	assign w_sys_tmp576 = w_fld_u_0_dataout_1;
	assign w_sys_tmp577 = (w_sys_tmp578 + r_run_k_17);
	assign w_sys_tmp578 = (r_run_copy0_j_30 * w_sys_tmp575);
	assign w_sys_tmp580 = (r_run_copy0_j_30 + w_sys_intOne);
	assign w_sys_tmp581 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp654 = 32'sh00000060;
	assign w_sys_tmp655 = ( !w_sys_tmp656 );
	assign w_sys_tmp656 = (w_sys_tmp657 < r_run_j_18);
	assign w_sys_tmp657 = 32'sh00000081;
	assign w_sys_tmp659 = (r_run_j_18 - w_sys_tmp660);
	assign w_sys_tmp660 = 32'sh0000005f;
	assign w_sys_tmp662 = (w_sys_tmp663 + r_run_k_17);
	assign w_sys_tmp663 = (r_run_tmpj_23 * w_sys_tmp664);
	assign w_sys_tmp664 = 32'sh00000081;
	assign w_sys_tmp665 = w_fld_u_0_dataout_1;
	assign w_sys_tmp666 = (w_sys_tmp667 + r_run_k_17);
	assign w_sys_tmp667 = (r_run_copy0_j_31 * w_sys_tmp664);
	assign w_sys_tmp669 = (r_run_copy0_j_31 + w_sys_intOne);
	assign w_sys_tmp670 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp743 = 32'sh00000040;
	assign w_sys_tmp744 = ( !w_sys_tmp745 );
	assign w_sys_tmp745 = (w_sys_tmp746 < r_run_k_17);
	assign w_sys_tmp746 = 32'sh00000061;
	assign w_sys_tmp747 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp748 = ( !w_sys_tmp749 );
	assign w_sys_tmp749 = (w_sys_tmp750 < r_run_j_18);
	assign w_sys_tmp750 = 32'sh00000021;
	assign w_sys_tmp753 = (w_sys_tmp754 + r_run_k_17);
	assign w_sys_tmp754 = (r_run_j_18 * w_sys_tmp755);
	assign w_sys_tmp755 = 32'sh00000081;
	assign w_sys_tmp756 = w_fld_u_0_dataout_1;
	assign w_sys_tmp757 = (w_sys_tmp758 + r_run_k_17);
	assign w_sys_tmp758 = (r_run_copy0_j_32 * w_sys_tmp755);
	assign w_sys_tmp760 = (r_run_copy0_j_32 + w_sys_intOne);
	assign w_sys_tmp761 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp822 = 32'sh00000020;
	assign w_sys_tmp823 = ( !w_sys_tmp824 );
	assign w_sys_tmp824 = (w_sys_tmp825 < r_run_j_18);
	assign w_sys_tmp825 = 32'sh00000041;
	assign w_sys_tmp827 = (r_run_j_18 - w_sys_tmp828);
	assign w_sys_tmp828 = 32'sh0000001f;
	assign w_sys_tmp830 = (w_sys_tmp831 + r_run_k_17);
	assign w_sys_tmp831 = (r_run_tmpj_23 * w_sys_tmp832);
	assign w_sys_tmp832 = 32'sh00000081;
	assign w_sys_tmp833 = w_fld_u_0_dataout_1;
	assign w_sys_tmp834 = (w_sys_tmp835 + r_run_k_17);
	assign w_sys_tmp835 = (r_run_copy0_j_33 * w_sys_tmp832);
	assign w_sys_tmp837 = (r_run_copy0_j_33 + w_sys_intOne);
	assign w_sys_tmp838 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp911 = 32'sh00000040;
	assign w_sys_tmp912 = ( !w_sys_tmp913 );
	assign w_sys_tmp913 = (w_sys_tmp914 < r_run_j_18);
	assign w_sys_tmp914 = 32'sh00000061;
	assign w_sys_tmp916 = (r_run_j_18 - w_sys_tmp917);
	assign w_sys_tmp917 = 32'sh0000003f;
	assign w_sys_tmp919 = (w_sys_tmp920 + r_run_k_17);
	assign w_sys_tmp920 = (r_run_tmpj_23 * w_sys_tmp921);
	assign w_sys_tmp921 = 32'sh00000081;
	assign w_sys_tmp922 = w_fld_u_0_dataout_1;
	assign w_sys_tmp923 = (w_sys_tmp924 + r_run_k_17);
	assign w_sys_tmp924 = (r_run_copy0_j_34 * w_sys_tmp921);
	assign w_sys_tmp926 = (r_run_copy0_j_34 + w_sys_intOne);
	assign w_sys_tmp927 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp1000 = 32'sh00000060;
	assign w_sys_tmp1001 = ( !w_sys_tmp1002 );
	assign w_sys_tmp1002 = (w_sys_tmp1003 < r_run_j_18);
	assign w_sys_tmp1003 = 32'sh00000081;
	assign w_sys_tmp1005 = (r_run_j_18 - w_sys_tmp1006);
	assign w_sys_tmp1006 = 32'sh0000005f;
	assign w_sys_tmp1008 = (w_sys_tmp1009 + r_run_k_17);
	assign w_sys_tmp1009 = (r_run_tmpj_23 * w_sys_tmp1010);
	assign w_sys_tmp1010 = 32'sh00000081;
	assign w_sys_tmp1011 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1012 = (w_sys_tmp1013 + r_run_k_17);
	assign w_sys_tmp1013 = (r_run_copy0_j_35 * w_sys_tmp1010);
	assign w_sys_tmp1015 = (r_run_copy0_j_35 + w_sys_intOne);
	assign w_sys_tmp1016 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp1089 = 32'sh00000060;
	assign w_sys_tmp1090 = ( !w_sys_tmp1091 );
	assign w_sys_tmp1091 = (w_sys_tmp1092 < r_run_k_17);
	assign w_sys_tmp1092 = 32'sh00000081;
	assign w_sys_tmp1093 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp1094 = ( !w_sys_tmp1095 );
	assign w_sys_tmp1095 = (w_sys_tmp1096 < r_run_j_18);
	assign w_sys_tmp1096 = 32'sh00000021;
	assign w_sys_tmp1099 = (w_sys_tmp1100 + r_run_k_17);
	assign w_sys_tmp1100 = (r_run_j_18 * w_sys_tmp1101);
	assign w_sys_tmp1101 = 32'sh00000081;
	assign w_sys_tmp1102 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1103 = (w_sys_tmp1104 + r_run_k_17);
	assign w_sys_tmp1104 = (r_run_copy0_j_36 * w_sys_tmp1101);
	assign w_sys_tmp1106 = (r_run_copy0_j_36 + w_sys_intOne);
	assign w_sys_tmp1107 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp1168 = 32'sh00000020;
	assign w_sys_tmp1169 = ( !w_sys_tmp1170 );
	assign w_sys_tmp1170 = (w_sys_tmp1171 < r_run_j_18);
	assign w_sys_tmp1171 = 32'sh00000041;
	assign w_sys_tmp1173 = (r_run_j_18 - w_sys_tmp1174);
	assign w_sys_tmp1174 = 32'sh0000001f;
	assign w_sys_tmp1176 = (w_sys_tmp1177 + r_run_k_17);
	assign w_sys_tmp1177 = (r_run_tmpj_23 * w_sys_tmp1178);
	assign w_sys_tmp1178 = 32'sh00000081;
	assign w_sys_tmp1179 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1180 = (w_sys_tmp1181 + r_run_k_17);
	assign w_sys_tmp1181 = (r_run_copy0_j_37 * w_sys_tmp1178);
	assign w_sys_tmp1183 = (r_run_copy0_j_37 + w_sys_intOne);
	assign w_sys_tmp1184 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp1257 = 32'sh00000040;
	assign w_sys_tmp1258 = ( !w_sys_tmp1259 );
	assign w_sys_tmp1259 = (w_sys_tmp1260 < r_run_j_18);
	assign w_sys_tmp1260 = 32'sh00000061;
	assign w_sys_tmp1262 = (r_run_j_18 - w_sys_tmp1263);
	assign w_sys_tmp1263 = 32'sh0000003f;
	assign w_sys_tmp1265 = (w_sys_tmp1266 + r_run_k_17);
	assign w_sys_tmp1266 = (r_run_tmpj_23 * w_sys_tmp1267);
	assign w_sys_tmp1267 = 32'sh00000081;
	assign w_sys_tmp1268 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1269 = (w_sys_tmp1270 + r_run_k_17);
	assign w_sys_tmp1270 = (r_run_copy0_j_38 * w_sys_tmp1267);
	assign w_sys_tmp1272 = (r_run_copy0_j_38 + w_sys_intOne);
	assign w_sys_tmp1273 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp1346 = 32'sh00000060;
	assign w_sys_tmp1347 = ( !w_sys_tmp1348 );
	assign w_sys_tmp1348 = (w_sys_tmp1349 < r_run_j_18);
	assign w_sys_tmp1349 = 32'sh00000081;
	assign w_sys_tmp1351 = (r_run_j_18 - w_sys_tmp1352);
	assign w_sys_tmp1352 = 32'sh0000005f;
	assign w_sys_tmp1354 = (w_sys_tmp1355 + r_run_k_17);
	assign w_sys_tmp1355 = (r_run_tmpj_23 * w_sys_tmp1356);
	assign w_sys_tmp1356 = 32'sh00000081;
	assign w_sys_tmp1357 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1358 = (w_sys_tmp1359 + r_run_k_17);
	assign w_sys_tmp1359 = (r_run_copy0_j_39 * w_sys_tmp1356);
	assign w_sys_tmp1361 = (r_run_copy0_j_39 + w_sys_intOne);
	assign w_sys_tmp1362 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp1435 = ( !w_sys_tmp1436 );
	assign w_sys_tmp1436 = (r_run_nlast_22 < r_run_n_19);
	assign w_sys_tmp1437 = (r_run_n_19 + w_sys_intOne);
	assign w_sys_tmp1438 = 32'sh00000002;
	assign w_sys_tmp1439 = ( !w_sys_tmp1440 );
	assign w_sys_tmp1440 = (w_sys_tmp1441 < r_run_k_17);
	assign w_sys_tmp1441 = 32'sh00000020;
	assign w_sys_tmp1444 = (w_sys_tmp1445 + r_run_k_17);
	assign w_sys_tmp1445 = 32'sh000010a1;
	assign w_sys_tmp1446 = w_sub01_result_dataout;
	assign w_sys_tmp1447 = (w_sys_tmp1448 + r_run_k_17);
	assign w_sys_tmp1448 = 32'sh00000102;
	assign w_sys_tmp1450 = (w_sys_tmp1451 + r_run_k_17);
	assign w_sys_tmp1451 = 32'sh00000081;
	assign w_sys_tmp1452 = w_sub00_result_dataout;
	assign w_sys_tmp1453 = (w_sys_tmp1454 + r_run_k_17);
	assign w_sys_tmp1454 = 32'sh00001020;
	assign w_sys_tmp1456 = (w_sys_tmp1457 + r_run_k_17);
	assign w_sys_tmp1457 = 32'sh00001122;
	assign w_sys_tmp1474 = w_sub02_result_dataout;
	assign w_sys_tmp1477 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp1478 = 32'sh00000021;
	assign w_sys_tmp1479 = ( !w_sys_tmp1480 );
	assign w_sys_tmp1480 = (w_sys_tmp1481 < r_run_k_17);
	assign w_sys_tmp1481 = 32'sh00000040;
	assign w_sys_tmp1484 = (w_sys_tmp1485 + r_run_k_17);
	assign w_sys_tmp1485 = 32'sh000010a1;
	assign w_sys_tmp1486 = w_sub05_result_dataout;
	assign w_sys_tmp1487 = (w_sys_tmp1488 + r_run_k_17);
	assign w_sys_tmp1488 = 32'sh00000102;
	assign w_sys_tmp1490 = (w_sys_tmp1491 + r_run_k_17);
	assign w_sys_tmp1491 = 32'sh00000081;
	assign w_sys_tmp1492 = w_sub04_result_dataout;
	assign w_sys_tmp1493 = (w_sys_tmp1494 + r_run_k_17);
	assign w_sys_tmp1494 = 32'sh00001020;
	assign w_sys_tmp1496 = (w_sys_tmp1497 + r_run_k_17);
	assign w_sys_tmp1497 = 32'sh00001122;
	assign w_sys_tmp1514 = w_sub06_result_dataout;
	assign w_sys_tmp1517 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp1518 = 32'sh00000041;
	assign w_sys_tmp1519 = ( !w_sys_tmp1520 );
	assign w_sys_tmp1520 = (w_sys_tmp1521 < r_run_k_17);
	assign w_sys_tmp1521 = 32'sh00000060;
	assign w_sys_tmp1524 = (w_sys_tmp1525 + r_run_k_17);
	assign w_sys_tmp1525 = 32'sh000010a1;
	assign w_sys_tmp1526 = w_sub09_result_dataout;
	assign w_sys_tmp1527 = (w_sys_tmp1528 + r_run_k_17);
	assign w_sys_tmp1528 = 32'sh00000102;
	assign w_sys_tmp1530 = (w_sys_tmp1531 + r_run_k_17);
	assign w_sys_tmp1531 = 32'sh00000081;
	assign w_sys_tmp1532 = w_sub08_result_dataout;
	assign w_sys_tmp1533 = (w_sys_tmp1534 + r_run_k_17);
	assign w_sys_tmp1534 = 32'sh00001020;
	assign w_sys_tmp1536 = (w_sys_tmp1537 + r_run_k_17);
	assign w_sys_tmp1537 = 32'sh00001122;
	assign w_sys_tmp1554 = w_sub10_result_dataout;
	assign w_sys_tmp1557 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp1558 = 32'sh00000061;
	assign w_sys_tmp1559 = ( !w_sys_tmp1560 );
	assign w_sys_tmp1560 = (w_sys_tmp1561 < r_run_k_17);
	assign w_sys_tmp1561 = 32'sh00000080;
	assign w_sys_tmp1564 = (w_sys_tmp1565 + r_run_k_17);
	assign w_sys_tmp1565 = 32'sh000010a1;
	assign w_sys_tmp1566 = w_sub13_result_dataout;
	assign w_sys_tmp1567 = (w_sys_tmp1568 + r_run_k_17);
	assign w_sys_tmp1568 = 32'sh00000102;
	assign w_sys_tmp1570 = (w_sys_tmp1571 + r_run_k_17);
	assign w_sys_tmp1571 = 32'sh00000081;
	assign w_sys_tmp1572 = w_sub12_result_dataout;
	assign w_sys_tmp1573 = (w_sys_tmp1574 + r_run_k_17);
	assign w_sys_tmp1574 = 32'sh00001020;
	assign w_sys_tmp1576 = (w_sys_tmp1577 + r_run_k_17);
	assign w_sys_tmp1577 = 32'sh00001122;
	assign w_sys_tmp1594 = w_sub14_result_dataout;
	assign w_sys_tmp1595 = (w_sys_tmp1596 + r_run_k_17);
	assign w_sys_tmp1596 = 32'sh00000183;
	assign w_sys_tmp1597 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp1598 = 32'sh00000002;
	assign w_sys_tmp1599 = ( !w_sys_tmp1600 );
	assign w_sys_tmp1600 = (w_sys_tmp1601 < r_run_j_18);
	assign w_sys_tmp1601 = 32'sh00000020;
	assign w_sys_tmp1604 = (w_sys_tmp1605 + w_sys_tmp1607);
	assign w_sys_tmp1605 = (r_run_j_18 * w_sys_tmp1606);
	assign w_sys_tmp1606 = 32'sh00000081;
	assign w_sys_tmp1607 = 32'sh00000021;
	assign w_sys_tmp1608 = w_sub04_result_dataout;
	assign w_sys_tmp1609 = (w_sys_tmp1610 + w_sys_tmp1607);
	assign w_sys_tmp1610 = (r_run_copy10_j_50 * w_sys_tmp1606);
	assign w_sys_tmp1614 = (w_sys_tmp1615 + w_sys_tmp1617);
	assign w_sys_tmp1615 = (r_run_copy9_j_49 * w_sys_tmp1606);
	assign w_sys_tmp1617 = 32'sh00000020;
	assign w_sys_tmp1618 = w_sub00_result_dataout;
	assign w_sys_tmp1619 = (w_sys_tmp1620 + w_sys_tmp1617);
	assign w_sys_tmp1620 = (r_run_copy8_j_48 * w_sys_tmp1606);
	assign w_sys_tmp1624 = (w_sys_tmp1625 + w_sys_tmp1627);
	assign w_sys_tmp1625 = (r_run_copy7_j_47 * w_sys_tmp1606);
	assign w_sys_tmp1627 = 32'sh00000041;
	assign w_sys_tmp1628 = (w_sys_tmp1629 + w_sys_tmp1627);
	assign w_sys_tmp1629 = (r_run_copy6_j_46 * w_sys_tmp1606);
	assign w_sys_tmp1633 = (w_sys_tmp1634 + w_sys_tmp1636);
	assign w_sys_tmp1634 = (r_run_copy5_j_45 * w_sys_tmp1606);
	assign w_sys_tmp1636 = 32'sh00000040;
	assign w_sys_tmp1638 = (w_sys_tmp1639 + w_sys_tmp1636);
	assign w_sys_tmp1639 = (r_run_copy4_j_44 * w_sys_tmp1606);
	assign w_sys_tmp1643 = (w_sys_tmp1644 + w_sys_tmp1646);
	assign w_sys_tmp1644 = (r_run_copy3_j_43 * w_sys_tmp1606);
	assign w_sys_tmp1646 = 32'sh00000061;
	assign w_sys_tmp1647 = (w_sys_tmp1648 + w_sys_tmp1646);
	assign w_sys_tmp1648 = (r_run_copy2_j_42 * w_sys_tmp1606);
	assign w_sys_tmp1652 = (w_sys_tmp1653 + w_sys_tmp1655);
	assign w_sys_tmp1653 = (r_run_copy1_j_41 * w_sys_tmp1606);
	assign w_sys_tmp1655 = 32'sh00000060;
	assign w_sys_tmp1656 = w_sub08_result_dataout;
	assign w_sys_tmp1657 = (w_sys_tmp1658 + w_sys_tmp1655);
	assign w_sys_tmp1658 = (r_run_copy0_j_40 * w_sys_tmp1606);
	assign w_sys_tmp1661 = (r_run_copy0_j_40 + w_sys_intOne);
	assign w_sys_tmp1662 = (r_run_copy1_j_41 + w_sys_intOne);
	assign w_sys_tmp1663 = (r_run_copy2_j_42 + w_sys_intOne);
	assign w_sys_tmp1664 = (r_run_copy3_j_43 + w_sys_intOne);
	assign w_sys_tmp1665 = (r_run_copy4_j_44 + w_sys_intOne);
	assign w_sys_tmp1666 = (r_run_copy5_j_45 + w_sys_intOne);
	assign w_sys_tmp1667 = (r_run_copy6_j_46 + w_sys_intOne);
	assign w_sys_tmp1668 = (r_run_copy7_j_47 + w_sys_intOne);
	assign w_sys_tmp1669 = (r_run_copy8_j_48 + w_sys_intOne);
	assign w_sys_tmp1670 = (r_run_copy9_j_49 + w_sys_intOne);
	assign w_sys_tmp1671 = (r_run_copy10_j_50 + w_sys_intOne);
	assign w_sys_tmp1672 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp2099 = 32'sh00000021;
	assign w_sys_tmp2100 = ( !w_sys_tmp2101 );
	assign w_sys_tmp2101 = (w_sys_tmp2102 < r_run_j_18);
	assign w_sys_tmp2102 = 32'sh00000040;
	assign w_sys_tmp2104 = (r_run_j_18 - w_sys_tmp2105);
	assign w_sys_tmp2105 = 32'sh0000001f;
	assign w_sys_tmp2107 = (w_sys_tmp2108 + w_sys_tmp2110);
	assign w_sys_tmp2108 = (r_run_tmpj_23 * w_sys_tmp2109);
	assign w_sys_tmp2109 = 32'sh00000081;
	assign w_sys_tmp2110 = 32'sh00000021;
	assign w_sys_tmp2111 = w_sub05_result_dataout;
	assign w_sys_tmp2112 = (w_sys_tmp2113 + w_sys_tmp2110);
	assign w_sys_tmp2113 = (w_sys_tmp2114 * w_sys_tmp2109);
	assign w_sys_tmp2114 = w_sys_tmp2104;
	assign w_sys_tmp2118 = (w_sys_tmp2108 + w_sys_tmp2121);
	assign w_sys_tmp2121 = 32'sh00000020;
	assign w_sys_tmp2122 = w_sub01_result_dataout;
	assign w_sys_tmp2128 = (w_sys_tmp2108 + w_sys_tmp2131);
	assign w_sys_tmp2131 = 32'sh00000041;
	assign w_sys_tmp2132 = (w_sys_tmp2113 + w_sys_tmp2131);
	assign w_sys_tmp2138 = (w_sys_tmp2108 + w_sys_tmp2141);
	assign w_sys_tmp2141 = 32'sh00000040;
	assign w_sys_tmp2148 = (w_sys_tmp2108 + w_sys_tmp2151);
	assign w_sys_tmp2151 = 32'sh00000061;
	assign w_sys_tmp2152 = (w_sys_tmp2113 + w_sys_tmp2151);
	assign w_sys_tmp2158 = (w_sys_tmp2108 + w_sys_tmp2161);
	assign w_sys_tmp2161 = 32'sh00000060;
	assign w_sys_tmp2162 = w_sub09_result_dataout;
	assign w_sys_tmp2167 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp2546 = 32'sh00000041;
	assign w_sys_tmp2547 = ( !w_sys_tmp2548 );
	assign w_sys_tmp2548 = (w_sys_tmp2549 < r_run_j_18);
	assign w_sys_tmp2549 = 32'sh00000060;
	assign w_sys_tmp2551 = (r_run_j_18 - w_sys_tmp2552);
	assign w_sys_tmp2552 = 32'sh0000003f;
	assign w_sys_tmp2554 = (w_sys_tmp2555 + w_sys_tmp2557);
	assign w_sys_tmp2555 = (r_run_tmpj_23 * w_sys_tmp2556);
	assign w_sys_tmp2556 = 32'sh00000081;
	assign w_sys_tmp2557 = 32'sh00000021;
	assign w_sys_tmp2558 = w_sub06_result_dataout;
	assign w_sys_tmp2559 = (w_sys_tmp2560 + w_sys_tmp2557);
	assign w_sys_tmp2560 = (w_sys_tmp2561 * w_sys_tmp2556);
	assign w_sys_tmp2561 = w_sys_tmp2551;
	assign w_sys_tmp2565 = (w_sys_tmp2555 + w_sys_tmp2568);
	assign w_sys_tmp2568 = 32'sh00000020;
	assign w_sys_tmp2569 = w_sub02_result_dataout;
	assign w_sys_tmp2575 = (w_sys_tmp2555 + w_sys_tmp2578);
	assign w_sys_tmp2578 = 32'sh00000041;
	assign w_sys_tmp2579 = (w_sys_tmp2560 + w_sys_tmp2578);
	assign w_sys_tmp2585 = (w_sys_tmp2555 + w_sys_tmp2588);
	assign w_sys_tmp2588 = 32'sh00000040;
	assign w_sys_tmp2595 = (w_sys_tmp2555 + w_sys_tmp2598);
	assign w_sys_tmp2598 = 32'sh00000061;
	assign w_sys_tmp2599 = (w_sys_tmp2560 + w_sys_tmp2598);
	assign w_sys_tmp2605 = (w_sys_tmp2555 + w_sys_tmp2608);
	assign w_sys_tmp2608 = 32'sh00000060;
	assign w_sys_tmp2609 = w_sub10_result_dataout;
	assign w_sys_tmp2614 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp2993 = 32'sh00000061;
	assign w_sys_tmp2994 = ( !w_sys_tmp2995 );
	assign w_sys_tmp2995 = (w_sys_tmp2996 < r_run_j_18);
	assign w_sys_tmp2996 = 32'sh00000080;
	assign w_sys_tmp2998 = (r_run_j_18 - w_sys_tmp2999);
	assign w_sys_tmp2999 = 32'sh0000005f;
	assign w_sys_tmp3001 = (w_sys_tmp3002 + w_sys_tmp3004);
	assign w_sys_tmp3002 = (r_run_tmpj_23 * w_sys_tmp3003);
	assign w_sys_tmp3003 = 32'sh00000081;
	assign w_sys_tmp3004 = 32'sh00000021;
	assign w_sys_tmp3005 = w_sub07_result_dataout;
	assign w_sys_tmp3006 = (w_sys_tmp3007 + w_sys_tmp3004);
	assign w_sys_tmp3007 = (w_sys_tmp3008 * w_sys_tmp3003);
	assign w_sys_tmp3008 = w_sys_tmp2998;
	assign w_sys_tmp3012 = (w_sys_tmp3002 + w_sys_tmp3015);
	assign w_sys_tmp3015 = 32'sh00000020;
	assign w_sys_tmp3016 = w_sub03_result_dataout;
	assign w_sys_tmp3022 = (w_sys_tmp3002 + w_sys_tmp3025);
	assign w_sys_tmp3025 = 32'sh00000041;
	assign w_sys_tmp3026 = (w_sys_tmp3007 + w_sys_tmp3025);
	assign w_sys_tmp3032 = (w_sys_tmp3002 + w_sys_tmp3035);
	assign w_sys_tmp3035 = 32'sh00000040;
	assign w_sys_tmp3042 = (w_sys_tmp3002 + w_sys_tmp3045);
	assign w_sys_tmp3045 = 32'sh00000061;
	assign w_sys_tmp3046 = (w_sys_tmp3007 + w_sys_tmp3045);
	assign w_sys_tmp3052 = (w_sys_tmp3002 + w_sys_tmp3055);
	assign w_sys_tmp3055 = 32'sh00000060;
	assign w_sys_tmp3056 = w_sub11_result_dataout;
	assign w_sys_tmp3061 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp3440 = 32'sh00000002;
	assign w_sys_tmp3441 = ( !w_sys_tmp3442 );
	assign w_sys_tmp3442 = (w_sys_tmp3443 < r_run_k_17);
	assign w_sys_tmp3443 = 32'sh00000020;
	assign w_sys_tmp3444 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp3445 = 32'sh00000002;
	assign w_sys_tmp3446 = ( !w_sys_tmp3447 );
	assign w_sys_tmp3447 = (w_sys_tmp3448 < r_run_j_18);
	assign w_sys_tmp3448 = 32'sh00000020;
	assign w_sys_tmp3451 = (w_sys_tmp3452 + r_run_k_17);
	assign w_sys_tmp3452 = (r_run_j_18 * w_sys_tmp3453);
	assign w_sys_tmp3453 = 32'sh00000081;
	assign w_sys_tmp3454 = w_sub00_result_dataout;
	assign w_sys_tmp3455 = (w_sys_tmp3456 + r_run_k_17);
	assign w_sys_tmp3456 = (r_run_copy0_j_51 * w_sys_tmp3453);
	assign w_sys_tmp3458 = (r_run_copy0_j_51 + w_sys_intOne);
	assign w_sys_tmp3459 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp3520 = 32'sh00000021;
	assign w_sys_tmp3521 = ( !w_sys_tmp3522 );
	assign w_sys_tmp3522 = (w_sys_tmp3523 < r_run_j_18);
	assign w_sys_tmp3523 = 32'sh00000040;
	assign w_sys_tmp3525 = (r_run_j_18 - w_sys_tmp3526);
	assign w_sys_tmp3526 = 32'sh0000001f;
	assign w_sys_tmp3528 = (w_sys_tmp3529 + r_run_k_17);
	assign w_sys_tmp3529 = (r_run_copy1_j_53 * w_sys_tmp3530);
	assign w_sys_tmp3530 = 32'sh00000081;
	assign w_sys_tmp3531 = w_sub01_result_dataout;
	assign w_sys_tmp3532 = (w_sys_tmp3533 + r_run_k_17);
	assign w_sys_tmp3533 = (r_run_copy0_j_52 * w_sys_tmp3530);
	assign w_sys_tmp3535 = (r_run_copy0_j_52 + w_sys_intOne);
	assign w_sys_tmp3536 = (r_run_copy1_j_53 + w_sys_intOne);
	assign w_sys_tmp3537 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp3616 = 32'sh00000041;
	assign w_sys_tmp3617 = ( !w_sys_tmp3618 );
	assign w_sys_tmp3618 = (w_sys_tmp3619 < r_run_j_18);
	assign w_sys_tmp3619 = 32'sh00000060;
	assign w_sys_tmp3621 = (r_run_j_18 - w_sys_tmp3622);
	assign w_sys_tmp3622 = 32'sh0000003f;
	assign w_sys_tmp3624 = (w_sys_tmp3625 + r_run_k_17);
	assign w_sys_tmp3625 = (r_run_copy1_j_55 * w_sys_tmp3626);
	assign w_sys_tmp3626 = 32'sh00000081;
	assign w_sys_tmp3627 = w_sub02_result_dataout;
	assign w_sys_tmp3628 = (w_sys_tmp3629 + r_run_k_17);
	assign w_sys_tmp3629 = (r_run_copy0_j_54 * w_sys_tmp3626);
	assign w_sys_tmp3631 = (r_run_copy0_j_54 + w_sys_intOne);
	assign w_sys_tmp3632 = (r_run_copy1_j_55 + w_sys_intOne);
	assign w_sys_tmp3633 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp3712 = 32'sh00000061;
	assign w_sys_tmp3713 = ( !w_sys_tmp3714 );
	assign w_sys_tmp3714 = (w_sys_tmp3715 < r_run_j_18);
	assign w_sys_tmp3715 = 32'sh00000080;
	assign w_sys_tmp3717 = (r_run_j_18 - w_sys_tmp3718);
	assign w_sys_tmp3718 = 32'sh0000005f;
	assign w_sys_tmp3720 = (w_sys_tmp3721 + r_run_k_17);
	assign w_sys_tmp3721 = (r_run_copy1_j_57 * w_sys_tmp3722);
	assign w_sys_tmp3722 = 32'sh00000081;
	assign w_sys_tmp3723 = w_sub03_result_dataout;
	assign w_sys_tmp3724 = (w_sys_tmp3725 + r_run_k_17);
	assign w_sys_tmp3725 = (r_run_copy0_j_56 * w_sys_tmp3722);
	assign w_sys_tmp3727 = (r_run_copy0_j_56 + w_sys_intOne);
	assign w_sys_tmp3728 = (r_run_copy1_j_57 + w_sys_intOne);
	assign w_sys_tmp3729 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp3808 = 32'sh00000021;
	assign w_sys_tmp3809 = ( !w_sys_tmp3810 );
	assign w_sys_tmp3810 = (w_sys_tmp3811 < r_run_k_17);
	assign w_sys_tmp3811 = 32'sh00000040;
	assign w_sys_tmp3812 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp3813 = 32'sh00000002;
	assign w_sys_tmp3814 = ( !w_sys_tmp3815 );
	assign w_sys_tmp3815 = (w_sys_tmp3816 < r_run_j_18);
	assign w_sys_tmp3816 = 32'sh00000020;
	assign w_sys_tmp3819 = (w_sys_tmp3820 + r_run_k_17);
	assign w_sys_tmp3820 = (r_run_j_18 * w_sys_tmp3821);
	assign w_sys_tmp3821 = 32'sh00000081;
	assign w_sys_tmp3822 = w_sub04_result_dataout;
	assign w_sys_tmp3823 = (w_sys_tmp3824 + r_run_k_17);
	assign w_sys_tmp3824 = (r_run_copy0_j_58 * w_sys_tmp3821);
	assign w_sys_tmp3826 = (r_run_copy0_j_58 + w_sys_intOne);
	assign w_sys_tmp3827 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp3888 = 32'sh00000021;
	assign w_sys_tmp3889 = ( !w_sys_tmp3890 );
	assign w_sys_tmp3890 = (w_sys_tmp3891 < r_run_j_18);
	assign w_sys_tmp3891 = 32'sh00000040;
	assign w_sys_tmp3893 = (r_run_j_18 - w_sys_tmp3894);
	assign w_sys_tmp3894 = 32'sh0000001f;
	assign w_sys_tmp3896 = (w_sys_tmp3897 + r_run_k_17);
	assign w_sys_tmp3897 = (r_run_copy1_j_60 * w_sys_tmp3898);
	assign w_sys_tmp3898 = 32'sh00000081;
	assign w_sys_tmp3899 = w_sub05_result_dataout;
	assign w_sys_tmp3900 = (w_sys_tmp3901 + r_run_k_17);
	assign w_sys_tmp3901 = (r_run_copy0_j_59 * w_sys_tmp3898);
	assign w_sys_tmp3903 = (r_run_copy0_j_59 + w_sys_intOne);
	assign w_sys_tmp3904 = (r_run_copy1_j_60 + w_sys_intOne);
	assign w_sys_tmp3905 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp3984 = 32'sh00000041;
	assign w_sys_tmp3985 = ( !w_sys_tmp3986 );
	assign w_sys_tmp3986 = (w_sys_tmp3987 < r_run_j_18);
	assign w_sys_tmp3987 = 32'sh00000060;
	assign w_sys_tmp3989 = (r_run_j_18 - w_sys_tmp3990);
	assign w_sys_tmp3990 = 32'sh0000003f;
	assign w_sys_tmp3992 = (w_sys_tmp3993 + r_run_k_17);
	assign w_sys_tmp3993 = (r_run_copy1_j_62 * w_sys_tmp3994);
	assign w_sys_tmp3994 = 32'sh00000081;
	assign w_sys_tmp3995 = w_sub06_result_dataout;
	assign w_sys_tmp3996 = (w_sys_tmp3997 + r_run_k_17);
	assign w_sys_tmp3997 = (r_run_copy0_j_61 * w_sys_tmp3994);
	assign w_sys_tmp3999 = (r_run_copy0_j_61 + w_sys_intOne);
	assign w_sys_tmp4000 = (r_run_copy1_j_62 + w_sys_intOne);
	assign w_sys_tmp4001 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp4080 = 32'sh00000061;
	assign w_sys_tmp4081 = ( !w_sys_tmp4082 );
	assign w_sys_tmp4082 = (w_sys_tmp4083 < r_run_j_18);
	assign w_sys_tmp4083 = 32'sh00000080;
	assign w_sys_tmp4085 = (r_run_j_18 - w_sys_tmp4086);
	assign w_sys_tmp4086 = 32'sh0000005f;
	assign w_sys_tmp4088 = (w_sys_tmp4089 + r_run_k_17);
	assign w_sys_tmp4089 = (r_run_copy1_j_64 * w_sys_tmp4090);
	assign w_sys_tmp4090 = 32'sh00000081;
	assign w_sys_tmp4091 = w_sub07_result_dataout;
	assign w_sys_tmp4092 = (w_sys_tmp4093 + r_run_k_17);
	assign w_sys_tmp4093 = (r_run_copy0_j_63 * w_sys_tmp4090);
	assign w_sys_tmp4095 = (r_run_copy0_j_63 + w_sys_intOne);
	assign w_sys_tmp4096 = (r_run_copy1_j_64 + w_sys_intOne);
	assign w_sys_tmp4097 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp4176 = 32'sh00000041;
	assign w_sys_tmp4177 = ( !w_sys_tmp4178 );
	assign w_sys_tmp4178 = (w_sys_tmp4179 < r_run_k_17);
	assign w_sys_tmp4179 = 32'sh00000060;
	assign w_sys_tmp4180 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp4181 = 32'sh00000002;
	assign w_sys_tmp4182 = ( !w_sys_tmp4183 );
	assign w_sys_tmp4183 = (w_sys_tmp4184 < r_run_j_18);
	assign w_sys_tmp4184 = 32'sh00000020;
	assign w_sys_tmp4187 = (w_sys_tmp4188 + r_run_k_17);
	assign w_sys_tmp4188 = (r_run_j_18 * w_sys_tmp4189);
	assign w_sys_tmp4189 = 32'sh00000081;
	assign w_sys_tmp4190 = w_sub08_result_dataout;
	assign w_sys_tmp4191 = (w_sys_tmp4192 + r_run_k_17);
	assign w_sys_tmp4192 = (r_run_copy0_j_65 * w_sys_tmp4189);
	assign w_sys_tmp4194 = (r_run_copy0_j_65 + w_sys_intOne);
	assign w_sys_tmp4195 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp4256 = 32'sh00000021;
	assign w_sys_tmp4257 = ( !w_sys_tmp4258 );
	assign w_sys_tmp4258 = (w_sys_tmp4259 < r_run_j_18);
	assign w_sys_tmp4259 = 32'sh00000040;
	assign w_sys_tmp4261 = (r_run_j_18 - w_sys_tmp4262);
	assign w_sys_tmp4262 = 32'sh0000001f;
	assign w_sys_tmp4264 = (w_sys_tmp4265 + r_run_k_17);
	assign w_sys_tmp4265 = (r_run_copy1_j_67 * w_sys_tmp4266);
	assign w_sys_tmp4266 = 32'sh00000081;
	assign w_sys_tmp4267 = w_sub09_result_dataout;
	assign w_sys_tmp4268 = (w_sys_tmp4269 + r_run_k_17);
	assign w_sys_tmp4269 = (r_run_copy0_j_66 * w_sys_tmp4266);
	assign w_sys_tmp4271 = (r_run_copy0_j_66 + w_sys_intOne);
	assign w_sys_tmp4272 = (r_run_copy1_j_67 + w_sys_intOne);
	assign w_sys_tmp4273 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp4352 = 32'sh00000041;
	assign w_sys_tmp4353 = ( !w_sys_tmp4354 );
	assign w_sys_tmp4354 = (w_sys_tmp4355 < r_run_j_18);
	assign w_sys_tmp4355 = 32'sh00000060;
	assign w_sys_tmp4357 = (r_run_j_18 - w_sys_tmp4358);
	assign w_sys_tmp4358 = 32'sh0000003f;
	assign w_sys_tmp4360 = (w_sys_tmp4361 + r_run_k_17);
	assign w_sys_tmp4361 = (r_run_copy1_j_69 * w_sys_tmp4362);
	assign w_sys_tmp4362 = 32'sh00000081;
	assign w_sys_tmp4363 = w_sub10_result_dataout;
	assign w_sys_tmp4364 = (w_sys_tmp4365 + r_run_k_17);
	assign w_sys_tmp4365 = (r_run_copy0_j_68 * w_sys_tmp4362);
	assign w_sys_tmp4367 = (r_run_copy0_j_68 + w_sys_intOne);
	assign w_sys_tmp4368 = (r_run_copy1_j_69 + w_sys_intOne);
	assign w_sys_tmp4369 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp4448 = 32'sh00000061;
	assign w_sys_tmp4449 = ( !w_sys_tmp4450 );
	assign w_sys_tmp4450 = (w_sys_tmp4451 < r_run_j_18);
	assign w_sys_tmp4451 = 32'sh00000080;
	assign w_sys_tmp4453 = (r_run_j_18 - w_sys_tmp4454);
	assign w_sys_tmp4454 = 32'sh0000005f;
	assign w_sys_tmp4456 = (w_sys_tmp4457 + r_run_k_17);
	assign w_sys_tmp4457 = (r_run_copy1_j_71 * w_sys_tmp4458);
	assign w_sys_tmp4458 = 32'sh00000081;
	assign w_sys_tmp4459 = w_sub11_result_dataout;
	assign w_sys_tmp4460 = (w_sys_tmp4461 + r_run_k_17);
	assign w_sys_tmp4461 = (r_run_copy0_j_70 * w_sys_tmp4458);
	assign w_sys_tmp4463 = (r_run_copy0_j_70 + w_sys_intOne);
	assign w_sys_tmp4464 = (r_run_copy1_j_71 + w_sys_intOne);
	assign w_sys_tmp4465 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp4544 = 32'sh00000061;
	assign w_sys_tmp4545 = ( !w_sys_tmp4546 );
	assign w_sys_tmp4546 = (w_sys_tmp4547 < r_run_k_17);
	assign w_sys_tmp4547 = 32'sh00000080;
	assign w_sys_tmp4548 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp4549 = 32'sh00000002;
	assign w_sys_tmp4550 = ( !w_sys_tmp4551 );
	assign w_sys_tmp4551 = (w_sys_tmp4552 < r_run_j_18);
	assign w_sys_tmp4552 = 32'sh00000020;
	assign w_sys_tmp4555 = (w_sys_tmp4556 + r_run_k_17);
	assign w_sys_tmp4556 = (r_run_j_18 * w_sys_tmp4557);
	assign w_sys_tmp4557 = 32'sh00000081;
	assign w_sys_tmp4558 = w_sub12_result_dataout;
	assign w_sys_tmp4559 = (w_sys_tmp4560 + r_run_k_17);
	assign w_sys_tmp4560 = (r_run_copy0_j_72 * w_sys_tmp4557);
	assign w_sys_tmp4562 = (r_run_copy0_j_72 + w_sys_intOne);
	assign w_sys_tmp4563 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp4624 = 32'sh00000021;
	assign w_sys_tmp4625 = ( !w_sys_tmp4626 );
	assign w_sys_tmp4626 = (w_sys_tmp4627 < r_run_j_18);
	assign w_sys_tmp4627 = 32'sh00000040;
	assign w_sys_tmp4629 = (r_run_j_18 - w_sys_tmp4630);
	assign w_sys_tmp4630 = 32'sh0000001f;
	assign w_sys_tmp4632 = (w_sys_tmp4633 + r_run_k_17);
	assign w_sys_tmp4633 = (r_run_copy1_j_74 * w_sys_tmp4634);
	assign w_sys_tmp4634 = 32'sh00000081;
	assign w_sys_tmp4635 = w_sub13_result_dataout;
	assign w_sys_tmp4636 = (w_sys_tmp4637 + r_run_k_17);
	assign w_sys_tmp4637 = (r_run_copy0_j_73 * w_sys_tmp4634);
	assign w_sys_tmp4639 = (r_run_copy0_j_73 + w_sys_intOne);
	assign w_sys_tmp4640 = (r_run_copy1_j_74 + w_sys_intOne);
	assign w_sys_tmp4641 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp4720 = 32'sh00000041;
	assign w_sys_tmp4721 = ( !w_sys_tmp4722 );
	assign w_sys_tmp4722 = (w_sys_tmp4723 < r_run_j_18);
	assign w_sys_tmp4723 = 32'sh00000060;
	assign w_sys_tmp4725 = (r_run_j_18 - w_sys_tmp4726);
	assign w_sys_tmp4726 = 32'sh0000003f;
	assign w_sys_tmp4728 = (w_sys_tmp4729 + r_run_k_17);
	assign w_sys_tmp4729 = (r_run_copy1_j_76 * w_sys_tmp4730);
	assign w_sys_tmp4730 = 32'sh00000081;
	assign w_sys_tmp4731 = w_sub14_result_dataout;
	assign w_sys_tmp4732 = (w_sys_tmp4733 + r_run_k_17);
	assign w_sys_tmp4733 = (r_run_copy0_j_75 * w_sys_tmp4730);
	assign w_sys_tmp4735 = (r_run_copy0_j_75 + w_sys_intOne);
	assign w_sys_tmp4736 = (r_run_copy1_j_76 + w_sys_intOne);
	assign w_sys_tmp4737 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp4816 = 32'sh00000061;
	assign w_sys_tmp4817 = ( !w_sys_tmp4818 );
	assign w_sys_tmp4818 = (w_sys_tmp4819 < r_run_j_18);
	assign w_sys_tmp4819 = 32'sh00000080;
	assign w_sys_tmp4821 = (r_run_j_18 - w_sys_tmp4822);
	assign w_sys_tmp4822 = 32'sh0000005f;
	assign w_sys_tmp4824 = (w_sys_tmp4825 + r_run_k_17);
	assign w_sys_tmp4825 = (r_run_copy1_j_78 * w_sys_tmp4826);
	assign w_sys_tmp4826 = 32'sh00000081;
	assign w_sys_tmp4827 = w_sub15_result_dataout;
	assign w_sys_tmp4828 = (w_sys_tmp4829 + r_run_k_17);
	assign w_sys_tmp4829 = (r_run_copy0_j_77 * w_sys_tmp4826);
	assign w_sys_tmp4831 = (r_run_copy0_j_77 + w_sys_intOne);
	assign w_sys_tmp4832 = (r_run_copy1_j_78 + w_sys_intOne);
	assign w_sys_tmp4833 = (r_run_j_18 + w_sys_intOne);


	sub09
		sub09_inst(
			.i_fld_result_1_addr_0 (w_sub09_result_addr),
			.i_fld_result_1_datain_0 (w_sub09_result_datain),
			.o_fld_result_1_dataout_0 (w_sub09_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub09_result_r_w),
			.i_fld_u_0_addr_0 (w_sub09_u_addr),
			.i_fld_u_0_datain_0 (w_sub09_u_datain),
			.o_fld_u_0_dataout_0 (w_sub09_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub09_u_r_w),
			.o_run_busy (w_sub09_run_busy),
			.i_run_req (r_sub09_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub08
		sub08_inst(
			.i_fld_result_1_addr_0 (w_sub08_result_addr),
			.i_fld_result_1_datain_0 (w_sub08_result_datain),
			.o_fld_result_1_dataout_0 (w_sub08_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub08_result_r_w),
			.i_fld_u_0_addr_0 (w_sub08_u_addr),
			.i_fld_u_0_datain_0 (w_sub08_u_datain),
			.o_fld_u_0_dataout_0 (w_sub08_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub08_u_r_w),
			.o_run_busy (w_sub08_run_busy),
			.i_run_req (r_sub08_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub12
		sub12_inst(
			.i_fld_result_1_addr_0 (w_sub12_result_addr),
			.i_fld_result_1_datain_0 (w_sub12_result_datain),
			.o_fld_result_1_dataout_0 (w_sub12_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub12_result_r_w),
			.i_fld_u_0_addr_0 (w_sub12_u_addr),
			.i_fld_u_0_datain_0 (w_sub12_u_datain),
			.o_fld_u_0_dataout_0 (w_sub12_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub12_u_r_w),
			.o_run_busy (w_sub12_run_busy),
			.i_run_req (r_sub12_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub03
		sub03_inst(
			.i_fld_result_1_addr_0 (w_sub03_result_addr),
			.i_fld_result_1_datain_0 (w_sub03_result_datain),
			.o_fld_result_1_dataout_0 (w_sub03_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub03_result_r_w),
			.i_fld_u_0_addr_0 (w_sub03_u_addr),
			.i_fld_u_0_datain_0 (w_sub03_u_datain),
			.o_fld_u_0_dataout_0 (w_sub03_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub03_u_r_w),
			.o_run_busy (w_sub03_run_busy),
			.i_run_req (r_sub03_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub02
		sub02_inst(
			.i_fld_result_1_addr_0 (w_sub02_result_addr),
			.i_fld_result_1_datain_0 (w_sub02_result_datain),
			.o_fld_result_1_dataout_0 (w_sub02_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub02_result_r_w),
			.i_fld_u_0_addr_0 (w_sub02_u_addr),
			.i_fld_u_0_datain_0 (w_sub02_u_datain),
			.o_fld_u_0_dataout_0 (w_sub02_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub02_u_r_w),
			.o_run_busy (w_sub02_run_busy),
			.i_run_req (r_sub02_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub11
		sub11_inst(
			.i_fld_result_1_addr_0 (w_sub11_result_addr),
			.i_fld_result_1_datain_0 (w_sub11_result_datain),
			.o_fld_result_1_dataout_0 (w_sub11_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub11_result_r_w),
			.i_fld_u_0_addr_0 (w_sub11_u_addr),
			.i_fld_u_0_datain_0 (w_sub11_u_datain),
			.o_fld_u_0_dataout_0 (w_sub11_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub11_u_r_w),
			.o_run_busy (w_sub11_run_busy),
			.i_run_req (r_sub11_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub14
		sub14_inst(
			.i_fld_result_1_addr_0 (w_sub14_result_addr),
			.i_fld_result_1_datain_0 (w_sub14_result_datain),
			.o_fld_result_1_dataout_0 (w_sub14_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub14_result_r_w),
			.i_fld_u_0_addr_0 (w_sub14_u_addr),
			.i_fld_u_0_datain_0 (w_sub14_u_datain),
			.o_fld_u_0_dataout_0 (w_sub14_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub14_u_r_w),
			.o_run_busy (w_sub14_run_busy),
			.i_run_req (r_sub14_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub01
		sub01_inst(
			.i_fld_result_1_addr_0 (w_sub01_result_addr),
			.i_fld_result_1_datain_0 (w_sub01_result_datain),
			.o_fld_result_1_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub01_result_r_w),
			.i_fld_u_0_addr_0 (w_sub01_u_addr),
			.i_fld_u_0_datain_0 (w_sub01_u_datain),
			.o_fld_u_0_dataout_0 (w_sub01_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub01_u_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub13
		sub13_inst(
			.i_fld_result_1_addr_0 (w_sub13_result_addr),
			.i_fld_result_1_datain_0 (w_sub13_result_datain),
			.o_fld_result_1_dataout_0 (w_sub13_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub13_result_r_w),
			.i_fld_u_0_addr_0 (w_sub13_u_addr),
			.i_fld_u_0_datain_0 (w_sub13_u_datain),
			.o_fld_u_0_dataout_0 (w_sub13_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub13_u_r_w),
			.o_run_busy (w_sub13_run_busy),
			.i_run_req (r_sub13_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub00
		sub00_inst(
			.i_fld_result_1_addr_0 (w_sub00_result_addr),
			.i_fld_result_1_datain_0 (w_sub00_result_datain),
			.o_fld_result_1_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub00_result_r_w),
			.i_fld_u_0_addr_0 (w_sub00_u_addr),
			.i_fld_u_0_datain_0 (w_sub00_u_datain),
			.o_fld_u_0_dataout_0 (w_sub00_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub00_u_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub07
		sub07_inst(
			.i_fld_result_1_addr_0 (w_sub07_result_addr),
			.i_fld_result_1_datain_0 (w_sub07_result_datain),
			.o_fld_result_1_dataout_0 (w_sub07_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub07_result_r_w),
			.i_fld_u_0_addr_0 (w_sub07_u_addr),
			.i_fld_u_0_datain_0 (w_sub07_u_datain),
			.o_fld_u_0_dataout_0 (w_sub07_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub07_u_r_w),
			.o_run_busy (w_sub07_run_busy),
			.i_run_req (r_sub07_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub06
		sub06_inst(
			.i_fld_result_1_addr_0 (w_sub06_result_addr),
			.i_fld_result_1_datain_0 (w_sub06_result_datain),
			.o_fld_result_1_dataout_0 (w_sub06_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub06_result_r_w),
			.i_fld_u_0_addr_0 (w_sub06_u_addr),
			.i_fld_u_0_datain_0 (w_sub06_u_datain),
			.o_fld_u_0_dataout_0 (w_sub06_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub06_u_r_w),
			.o_run_busy (w_sub06_run_busy),
			.i_run_req (r_sub06_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub15
		sub15_inst(
			.i_fld_result_1_addr_0 (w_sub15_result_addr),
			.i_fld_result_1_datain_0 (w_sub15_result_datain),
			.o_fld_result_1_dataout_0 (w_sub15_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub15_result_r_w),
			.i_fld_u_0_addr_0 (w_sub15_u_addr),
			.i_fld_u_0_datain_0 (w_sub15_u_datain),
			.o_fld_u_0_dataout_0 (w_sub15_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub15_u_r_w),
			.o_run_busy (w_sub15_run_busy),
			.i_run_req (r_sub15_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub05
		sub05_inst(
			.i_fld_result_1_addr_0 (w_sub05_result_addr),
			.i_fld_result_1_datain_0 (w_sub05_result_datain),
			.o_fld_result_1_dataout_0 (w_sub05_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub05_result_r_w),
			.i_fld_u_0_addr_0 (w_sub05_u_addr),
			.i_fld_u_0_datain_0 (w_sub05_u_datain),
			.o_fld_u_0_dataout_0 (w_sub05_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub05_u_r_w),
			.o_run_busy (w_sub05_run_busy),
			.i_run_req (r_sub05_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub04
		sub04_inst(
			.i_fld_result_1_addr_0 (w_sub04_result_addr),
			.i_fld_result_1_datain_0 (w_sub04_result_datain),
			.o_fld_result_1_dataout_0 (w_sub04_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub04_result_r_w),
			.i_fld_u_0_addr_0 (w_sub04_u_addr),
			.i_fld_u_0_datain_0 (w_sub04_u_datain),
			.o_fld_u_0_dataout_0 (w_sub04_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub04_u_r_w),
			.o_run_busy (w_sub04_run_busy),
			.i_run_req (r_sub04_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub10
		sub10_inst(
			.i_fld_result_1_addr_0 (w_sub10_result_addr),
			.i_fld_result_1_datain_0 (w_sub10_result_datain),
			.o_fld_result_1_dataout_0 (w_sub10_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub10_result_r_w),
			.i_fld_u_0_addr_0 (w_sub10_u_addr),
			.i_fld_u_0_datain_0 (w_sub10_u_datain),
			.o_fld_u_0_dataout_0 (w_sub10_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub10_u_r_w),
			.o_run_busy (w_sub10_run_busy),
			.i_run_req (r_sub10_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_u_0(
			.clk (clock),
			.ce_0 (w_fld_u_0_ce_0),
			.addr_0 (w_fld_u_0_addr_0),
			.datain_0 (w_fld_u_0_datain_0),
			.dataout_0 (w_fld_u_0_dataout_0),
			.r_w_0 (w_fld_u_0_r_w_0),
			.ce_1 (w_fld_u_0_ce_1),
			.addr_1 (r_fld_u_0_addr_1),
			.datain_1 (r_fld_u_0_datain_1),
			.dataout_1 (w_fld_u_0_dataout_1),
			.r_w_1 (r_fld_u_0_r_w_1)
		);

	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						9'h12f: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 9'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h0: begin
							r_sys_run_phase <= 9'h2;
						end

						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h4;

									end
								end

							endcase
						end

						9'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h5;

									end
								end

							endcase
						end

						9'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4) ? 9'h9 : 9'hf);

									end
								end

							endcase
						end

						9'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h5;

									end
								end

							endcase
						end

						9'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'ha;

									end
								end

							endcase
						end

						9'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7) ? 9'hd : 9'h6);

									end
								end

							endcase
						end

						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_run_phase <= 9'ha;

									end
								end

							endcase
						end

						9'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h10;

									end
								end

							endcase
						end

						9'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp52) ? 9'h14 : 9'h2c);

									end
								end

							endcase
						end

						9'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h10;

									end
								end

							endcase
						end

						9'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h15;

									end
								end

							endcase
						end

						9'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp56) ? 9'h18 : 9'h1a);

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h15;

									end
								end

							endcase
						end

						9'h1a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h1b;

									end
								end

							endcase
						end

						9'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp131) ? 9'h1e : 9'h20);

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h1b;

									end
								end

							endcase
						end

						9'h20: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h21;

									end
								end

							endcase
						end

						9'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp220) ? 9'h24 : 9'h26);

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h21;

									end
								end

							endcase
						end

						9'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h27;

									end
								end

							endcase
						end

						9'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp309) ? 9'h2a : 9'h11);

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h27;

									end
								end

							endcase
						end

						9'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h2d;

									end
								end

							endcase
						end

						9'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp398) ? 9'h31 : 9'h49);

									end
								end

							endcase
						end

						9'h2e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h2d;

									end
								end

							endcase
						end

						9'h31: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h32;

									end
								end

							endcase
						end

						9'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp402) ? 9'h35 : 9'h37);

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h32;

									end
								end

							endcase
						end

						9'h37: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h38;

									end
								end

							endcase
						end

						9'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp477) ? 9'h3b : 9'h3d);

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h38;

									end
								end

							endcase
						end

						9'h3d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h3e;

									end
								end

							endcase
						end

						9'h3e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp566) ? 9'h41 : 9'h43);

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h3e;

									end
								end

							endcase
						end

						9'h43: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h44;

									end
								end

							endcase
						end

						9'h44: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp655) ? 9'h47 : 9'h2e);

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h44;

									end
								end

							endcase
						end

						9'h49: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h4a;

									end
								end

							endcase
						end

						9'h4a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp744) ? 9'h4e : 9'h66);

									end
								end

							endcase
						end

						9'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h4a;

									end
								end

							endcase
						end

						9'h4e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h4f;

									end
								end

							endcase
						end

						9'h4f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp748) ? 9'h52 : 9'h54);

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h4f;

									end
								end

							endcase
						end

						9'h54: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h55;

									end
								end

							endcase
						end

						9'h55: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp823) ? 9'h58 : 9'h5a);

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h55;

									end
								end

							endcase
						end

						9'h5a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h5b;

									end
								end

							endcase
						end

						9'h5b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp912) ? 9'h5e : 9'h60);

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h5b;

									end
								end

							endcase
						end

						9'h60: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h61;

									end
								end

							endcase
						end

						9'h61: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1001) ? 9'h64 : 9'h4b);

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h61;

									end
								end

							endcase
						end

						9'h66: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h67;

									end
								end

							endcase
						end

						9'h67: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1090) ? 9'h6b : 9'h83);

									end
								end

							endcase
						end

						9'h68: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h67;

									end
								end

							endcase
						end

						9'h6b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h6c;

									end
								end

							endcase
						end

						9'h6c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1094) ? 9'h6f : 9'h71);

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h6c;

									end
								end

							endcase
						end

						9'h71: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h72;

									end
								end

							endcase
						end

						9'h72: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1169) ? 9'h75 : 9'h77);

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h72;

									end
								end

							endcase
						end

						9'h77: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h78;

									end
								end

							endcase
						end

						9'h78: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1258) ? 9'h7b : 9'h7d);

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h78;

									end
								end

							endcase
						end

						9'h7d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h7e;

									end
								end

							endcase
						end

						9'h7e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1347) ? 9'h81 : 9'h68);

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h7e;

									end
								end

							endcase
						end

						9'h83: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h84;

									end
								end

							endcase
						end

						9'h84: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1435) ? 9'h87 : 9'hbb);

									end
								end

							endcase
						end

						9'h85: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h84;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h10: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_phase <= 9'h89;

									end
								end

							endcase
						end

						9'h89: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_phase <= 9'h8b;

									end
								end

							endcase
						end

						9'h8b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h8c;

									end
								end

							endcase
						end

						9'h8c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1439) ? 9'h8f : 9'h91);

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_phase <= 9'h8c;

									end
								end

							endcase
						end

						9'h91: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h92;

									end
								end

							endcase
						end

						9'h92: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1479) ? 9'h95 : 9'h97);

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_phase <= 9'h92;

									end
								end

							endcase
						end

						9'h97: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h98;

									end
								end

							endcase
						end

						9'h98: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1519) ? 9'h9b : 9'h9d);

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_phase <= 9'h98;

									end
								end

							endcase
						end

						9'h9d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h9e;

									end
								end

							endcase
						end

						9'h9e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1559) ? 9'ha1 : 9'ha3);

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_phase <= 9'h9e;

									end
								end

							endcase
						end

						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'ha4;

									end
								end

							endcase
						end

						9'ha4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1599) ? 9'ha7 : 9'ha9);

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3d)) begin
										r_sys_run_phase <= 9'ha4;

									end
								end

							endcase
						end

						9'ha9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'haa;

									end
								end

							endcase
						end

						9'haa: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2100) ? 9'had : 9'haf);

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5b)) begin
										r_sys_run_phase <= 9'haa;

									end
								end

							endcase
						end

						9'haf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hb0;

									end
								end

							endcase
						end

						9'hb0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2547) ? 9'hb3 : 9'hb5);

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5b)) begin
										r_sys_run_phase <= 9'hb0;

									end
								end

							endcase
						end

						9'hb5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hb6;

									end
								end

							endcase
						end

						9'hb6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2994) ? 9'hb9 : 9'h85);

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5b)) begin
										r_sys_run_phase <= 9'hb6;

									end
								end

							endcase
						end

						9'hbb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hbc;

									end
								end

							endcase
						end

						9'hbc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3441) ? 9'hc0 : 9'hd8);

									end
								end

							endcase
						end

						9'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hbc;

									end
								end

							endcase
						end

						9'hc0: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hc1;

									end
								end

							endcase
						end

						9'hc1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3446) ? 9'hc4 : 9'hc6);

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'hc1;

									end
								end

							endcase
						end

						9'hc6: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hc7;

									end
								end

							endcase
						end

						9'hc7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3521) ? 9'hca : 9'hcc);

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'hc7;

									end
								end

							endcase
						end

						9'hcc: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hcd;

									end
								end

							endcase
						end

						9'hcd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3617) ? 9'hd0 : 9'hd2);

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'hcd;

									end
								end

							endcase
						end

						9'hd2: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hd3;

									end
								end

							endcase
						end

						9'hd3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3713) ? 9'hd6 : 9'hbd);

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'hd3;

									end
								end

							endcase
						end

						9'hd8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hd9;

									end
								end

							endcase
						end

						9'hd9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3809) ? 9'hdd : 9'hf5);

									end
								end

							endcase
						end

						9'hda: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hd9;

									end
								end

							endcase
						end

						9'hdd: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hde;

									end
								end

							endcase
						end

						9'hde: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3814) ? 9'he1 : 9'he3);

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'hde;

									end
								end

							endcase
						end

						9'he3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'he4;

									end
								end

							endcase
						end

						9'he4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3889) ? 9'he7 : 9'he9);

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'he4;

									end
								end

							endcase
						end

						9'he9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hea;

									end
								end

							endcase
						end

						9'hea: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3985) ? 9'hed : 9'hef);

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'hea;

									end
								end

							endcase
						end

						9'hef: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hf0;

									end
								end

							endcase
						end

						9'hf0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4081) ? 9'hf3 : 9'hda);

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'hf0;

									end
								end

							endcase
						end

						9'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hf6;

									end
								end

							endcase
						end

						9'hf6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4177) ? 9'hfa : 9'h112);

									end
								end

							endcase
						end

						9'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hf6;

									end
								end

							endcase
						end

						9'hfa: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hfb;

									end
								end

							endcase
						end

						9'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4182) ? 9'hfe : 9'h100);

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'hfb;

									end
								end

							endcase
						end

						9'h100: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h101;

									end
								end

							endcase
						end

						9'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4257) ? 9'h104 : 9'h106);

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h101;

									end
								end

							endcase
						end

						9'h106: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h107;

									end
								end

							endcase
						end

						9'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4353) ? 9'h10a : 9'h10c);

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h107;

									end
								end

							endcase
						end

						9'h10c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h10d;

									end
								end

							endcase
						end

						9'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4449) ? 9'h110 : 9'hf7);

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h10d;

									end
								end

							endcase
						end

						9'h112: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h113;

									end
								end

							endcase
						end

						9'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4545) ? 9'h117 : 9'h12f);

									end
								end

							endcase
						end

						9'h114: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h113;

									end
								end

							endcase
						end

						9'h117: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h118;

									end
								end

							endcase
						end

						9'h118: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4550) ? 9'h11b : 9'h11d);

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h118;

									end
								end

							endcase
						end

						9'h11d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h11e;

									end
								end

							endcase
						end

						9'h11e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4625) ? 9'h121 : 9'h123);

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h11e;

									end
								end

							endcase
						end

						9'h123: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h124;

									end
								end

							endcase
						end

						9'h124: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4721) ? 9'h127 : 9'h129);

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h124;

									end
								end

							endcase
						end

						9'h129: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h12a;

									end
								end

							endcase
						end

						9'h12a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4817) ? 9'h12d : 9'h114);

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h12a;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sys_run_phase <= 9'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 5'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h2e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h31: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h37: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h3e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h43: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h44: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h49: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h4a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h4e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h4f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h54: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h55: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h5a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h5b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h60: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h61: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h66: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h67: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h68: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h6c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h72: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h78: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h7d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h7e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h83: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h84: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h85: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h89: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h8b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h8c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h91: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h92: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h97: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h98: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h9d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h9e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'haa: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5b)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'haf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hb0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5b)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hb5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hb6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5b)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hbb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hbc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hc0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hc1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hc6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hc7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hcc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hcd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hda: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hdd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hde: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'he3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'he4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'he9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hea: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hfa: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h100: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h106: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h10c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h112: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h114: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h117: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h118: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h11d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h11e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h123: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h124: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h129: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h12a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 7'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h5)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h2e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h31: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h37: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h3e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h43: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h44: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h49: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h4a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h4e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h4f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h54: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h55: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h5a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h5b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h60: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h61: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h66: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h67: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h68: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h6c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h72: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h78: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h7d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h7e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h83: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h84: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h85: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h89: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub00_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub01_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub02_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub03_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub04_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub05_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub06_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub07_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub08_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub09_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub10_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub11_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub12_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub13_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub14_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub15_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h8b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h8c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'hc)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h91: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h92: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'hc)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h97: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h98: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'hc)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h9d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h9e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'hc)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'ha3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'ha4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3d)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'ha9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'haa: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h5a)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h5b)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'haf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hb0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5b)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h5a)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hb5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hb6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5b)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h5a)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hbb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hbc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hc0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hc1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hc6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hc7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hcc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hcd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hd2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hd3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hd8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hd9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hda: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hdd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hde: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'he3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'he4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'he9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hea: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hf0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hf6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hfa: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h100: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h106: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h10c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h112: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h114: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h117: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h118: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h11d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h11e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h123: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h124: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h129: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h12a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						9'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						9'h12f: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp11[14:0] );

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp65[14:0] );

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp142[14:0] );

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp231[14:0] );

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp320[14:0] );

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp411[14:0] );

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp488[14:0] );

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp577[14:0] );

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp666[14:0] );

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp757[14:0] );

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp834[14:0] );

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp923[14:0] );

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1012[14:0] );

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1103[14:0] );

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1180[14:0] );

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1269[14:0] );

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1358[14:0] );

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3451[14:0] );

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3528[14:0] );

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3624[14:0] );

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3720[14:0] );

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3819[14:0] );

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3896[14:0] );

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3992[14:0] );

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4088[14:0] );

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4187[14:0] );

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4264[14:0] );

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4360[14:0] );

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4456[14:0] );

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4555[14:0] );

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4632[14:0] );

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4728[14:0] );

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4824[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp14;

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp3454;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp3531;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp3627;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp3723;

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp3822;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp3899;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp3995;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp4091;

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp4190;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp4267;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp4363;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp4459;

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp4558;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp4635;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp4731;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp4827;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h12f: begin
							r_fld_u_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_17 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_17 <= w_sys_tmp6;

									end
								end

							endcase
						end

						9'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_17 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_17 <= w_sys_tmp55;

									end
								end

							endcase
						end

						9'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_17 <= w_sys_tmp397;

									end
								end

							endcase
						end

						9'h2e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_17 <= w_sys_tmp401;

									end
								end

							endcase
						end

						9'h49: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_17 <= w_sys_tmp743;

									end
								end

							endcase
						end

						9'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_17 <= w_sys_tmp747;

									end
								end

							endcase
						end

						9'h66: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_17 <= w_sys_tmp1089;

									end
								end

							endcase
						end

						9'h68: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_17 <= w_sys_tmp1093;

									end
								end

							endcase
						end

						9'h8b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_17 <= w_sys_tmp1438;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_run_k_17 <= w_sys_tmp1477;

									end
								end

							endcase
						end

						9'h91: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_17 <= w_sys_tmp1478;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_run_k_17 <= w_sys_tmp1517;

									end
								end

							endcase
						end

						9'h97: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_17 <= w_sys_tmp1518;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_run_k_17 <= w_sys_tmp1557;

									end
								end

							endcase
						end

						9'h9d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_17 <= w_sys_tmp1558;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_run_k_17 <= w_sys_tmp1597;

									end
								end

							endcase
						end

						9'hbb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_17 <= w_sys_tmp3440;

									end
								end

							endcase
						end

						9'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_17 <= w_sys_tmp3444;

									end
								end

							endcase
						end

						9'hd8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_17 <= w_sys_tmp3808;

									end
								end

							endcase
						end

						9'hda: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_17 <= w_sys_tmp3812;

									end
								end

							endcase
						end

						9'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_17 <= w_sys_tmp4176;

									end
								end

							endcase
						end

						9'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_17 <= w_sys_tmp4180;

									end
								end

							endcase
						end

						9'h112: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_17 <= w_sys_tmp4544;

									end
								end

							endcase
						end

						9'h114: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_17 <= w_sys_tmp4548;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_18 <= w_sys_tmp15;

									end
								end

							endcase
						end

						9'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_j_18 <= w_sys_tmp69;

									end
								end

							endcase
						end

						9'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp130;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_run_j_18 <= w_sys_tmp146;

									end
								end

							endcase
						end

						9'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp219;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_run_j_18 <= w_sys_tmp235;

									end
								end

							endcase
						end

						9'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp308;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_run_j_18 <= w_sys_tmp324;

									end
								end

							endcase
						end

						9'h31: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_j_18 <= w_sys_tmp415;

									end
								end

							endcase
						end

						9'h37: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp476;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_run_j_18 <= w_sys_tmp492;

									end
								end

							endcase
						end

						9'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp565;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_run_j_18 <= w_sys_tmp581;

									end
								end

							endcase
						end

						9'h43: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp654;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_run_j_18 <= w_sys_tmp670;

									end
								end

							endcase
						end

						9'h4e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_j_18 <= w_sys_tmp761;

									end
								end

							endcase
						end

						9'h54: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp822;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_run_j_18 <= w_sys_tmp838;

									end
								end

							endcase
						end

						9'h5a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp911;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_run_j_18 <= w_sys_tmp927;

									end
								end

							endcase
						end

						9'h60: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp1000;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_run_j_18 <= w_sys_tmp1016;

									end
								end

							endcase
						end

						9'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_j_18 <= w_sys_tmp1107;

									end
								end

							endcase
						end

						9'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp1168;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_run_j_18 <= w_sys_tmp1184;

									end
								end

							endcase
						end

						9'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp1257;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_run_j_18 <= w_sys_tmp1273;

									end
								end

							endcase
						end

						9'h7d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp1346;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_run_j_18 <= w_sys_tmp1362;

									end
								end

							endcase
						end

						9'ha3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp1598;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h32)) begin
										r_run_j_18 <= w_sys_tmp1672;

									end
								end

							endcase
						end

						9'ha9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp2099;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e)) begin
										r_run_j_18 <= w_sys_tmp2167;

									end
								end

							endcase
						end

						9'haf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp2546;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e)) begin
										r_run_j_18 <= w_sys_tmp2614;

									end
								end

							endcase
						end

						9'hb5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp2993;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e)) begin
										r_run_j_18 <= w_sys_tmp3061;

									end
								end

							endcase
						end

						9'hc0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp3445;

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_j_18 <= w_sys_tmp3459;

									end
								end

							endcase
						end

						9'hc6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp3520;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_18 <= w_sys_tmp3537;

									end
								end

							endcase
						end

						9'hcc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp3616;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_18 <= w_sys_tmp3633;

									end
								end

							endcase
						end

						9'hd2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp3712;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_18 <= w_sys_tmp3729;

									end
								end

							endcase
						end

						9'hdd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp3813;

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_j_18 <= w_sys_tmp3827;

									end
								end

							endcase
						end

						9'he3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp3888;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_18 <= w_sys_tmp3905;

									end
								end

							endcase
						end

						9'he9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp3984;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_18 <= w_sys_tmp4001;

									end
								end

							endcase
						end

						9'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp4080;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_18 <= w_sys_tmp4097;

									end
								end

							endcase
						end

						9'hfa: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp4181;

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_j_18 <= w_sys_tmp4195;

									end
								end

							endcase
						end

						9'h100: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp4256;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_18 <= w_sys_tmp4273;

									end
								end

							endcase
						end

						9'h106: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp4352;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_18 <= w_sys_tmp4369;

									end
								end

							endcase
						end

						9'h10c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp4448;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_18 <= w_sys_tmp4465;

									end
								end

							endcase
						end

						9'h117: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp4549;

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_j_18 <= w_sys_tmp4563;

									end
								end

							endcase
						end

						9'h11d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp4624;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_18 <= w_sys_tmp4641;

									end
								end

							endcase
						end

						9'h123: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp4720;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_18 <= w_sys_tmp4737;

									end
								end

							endcase
						end

						9'h129: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_18 <= w_sys_tmp4816;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_18 <= w_sys_tmp4833;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h83: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_n_19 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h85: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_n_19 <= w_sys_tmp1437;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_mx_20 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_my_21 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_nlast_22 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_run_tmpj_23 <= w_sys_tmp135;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_run_tmpj_23 <= w_sys_tmp224;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_run_tmpj_23 <= w_sys_tmp313;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_run_tmpj_23 <= w_sys_tmp481;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_run_tmpj_23 <= w_sys_tmp570;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_run_tmpj_23 <= w_sys_tmp659;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_run_tmpj_23 <= w_sys_tmp827;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_run_tmpj_23 <= w_sys_tmp916;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_run_tmpj_23 <= w_sys_tmp1005;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_run_tmpj_23 <= w_sys_tmp1173;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_run_tmpj_23 <= w_sys_tmp1262;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_run_tmpj_23 <= w_sys_tmp1351;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e)) begin
										r_run_tmpj_23 <= w_sys_tmp2104;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e)) begin
										r_run_tmpj_23 <= w_sys_tmp2551;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e)) begin
										r_run_tmpj_23 <= w_sys_tmp2998;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_tmpj_23 <= w_sys_tmp3525;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_tmpj_23 <= w_sys_tmp3621;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_tmpj_23 <= w_sys_tmp3717;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_tmpj_23 <= w_sys_tmp3893;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_tmpj_23 <= w_sys_tmp3989;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_tmpj_23 <= w_sys_tmp4085;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_tmpj_23 <= w_sys_tmp4261;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_tmpj_23 <= w_sys_tmp4357;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_tmpj_23 <= w_sys_tmp4453;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_tmpj_23 <= w_sys_tmp4629;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_tmpj_23 <= w_sys_tmp4725;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_tmpj_23 <= w_sys_tmp4821;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_24 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_24 <= w_sys_tmp68;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_25 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_25 <= w_sys_tmp145;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h20: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_26 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_26 <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_27 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_27 <= w_sys_tmp323;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h31: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_28 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_28 <= w_sys_tmp414;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h37: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_29 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_29 <= w_sys_tmp491;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_30 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_30 <= w_sys_tmp580;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h43: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_31 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_31 <= w_sys_tmp669;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h4e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_32 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_32 <= w_sys_tmp760;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h54: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_33 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_33 <= w_sys_tmp837;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_34 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_34 <= w_sys_tmp926;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h60: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_35 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_35 <= w_sys_tmp1015;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_36 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_36 <= w_sys_tmp1106;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h71: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_37 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_37 <= w_sys_tmp1183;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h77: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_38 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_38 <= w_sys_tmp1272;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_39 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_39 <= w_sys_tmp1361;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_40 <= r_run_j_18;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hb) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h2b) || (r_sys_run_step==7'h33) || (r_sys_run_step==7'h3b)) begin
										r_run_copy0_j_40 <= w_sys_tmp1661;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_41 <= r_run_j_18;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h3d)) begin
										r_run_copy1_j_41 <= w_sys_tmp1662;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy2_j_42 <= r_run_j_18;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h36)) begin
										r_run_copy2_j_42 <= w_sys_tmp1663;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy3_j_43 <= r_run_j_18;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h3a)) begin
										r_run_copy3_j_43 <= w_sys_tmp1664;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy4_j_44 <= r_run_j_18;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h7) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h2f) || (r_sys_run_step==7'h37)) begin
										r_run_copy4_j_44 <= w_sys_tmp1665;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy5_j_45 <= r_run_j_18;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h39)) begin
										r_run_copy5_j_45 <= w_sys_tmp1666;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy6_j_46 <= r_run_j_18;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h34)) begin
										r_run_copy6_j_46 <= w_sys_tmp1667;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy7_j_47 <= r_run_j_18;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h36)) begin
										r_run_copy7_j_47 <= w_sys_tmp1668;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy8_j_48 <= r_run_j_18;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h2b) || (r_sys_run_step==7'h33)) begin
										r_run_copy8_j_48 <= w_sys_tmp1669;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy9_j_49 <= r_run_j_18;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h35)) begin
										r_run_copy9_j_49 <= w_sys_tmp1670;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy10_j_50 <= r_run_j_18;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h30)) begin
										r_run_copy10_j_50 <= w_sys_tmp1671;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hc0: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_51 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_51 <= w_sys_tmp3458;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hc6: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_52 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_52 <= w_sys_tmp3535;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hc6: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_53 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_53 <= w_sys_tmp3536;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hcc: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_54 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_54 <= w_sys_tmp3631;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hcc: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_55 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_55 <= w_sys_tmp3632;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd2: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_56 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_56 <= w_sys_tmp3727;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd2: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_57 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_57 <= w_sys_tmp3728;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hdd: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_58 <= r_run_j_18;

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_58 <= w_sys_tmp3826;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'he3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_59 <= r_run_j_18;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_59 <= w_sys_tmp3903;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'he3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_60 <= r_run_j_18;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_60 <= w_sys_tmp3904;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'he9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_61 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_61 <= w_sys_tmp3999;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'he9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_62 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_62 <= w_sys_tmp4000;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hef: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_63 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_63 <= w_sys_tmp4095;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hef: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_64 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_64 <= w_sys_tmp4096;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hfa: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_65 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_65 <= w_sys_tmp4194;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h100: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_66 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_66 <= w_sys_tmp4271;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h100: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_67 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_67 <= w_sys_tmp4272;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h106: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_68 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_68 <= w_sys_tmp4367;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h106: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_69 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_69 <= w_sys_tmp4368;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h10c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_70 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_70 <= w_sys_tmp4463;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h10c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_71 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_71 <= w_sys_tmp4464;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h117: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_72 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_72 <= w_sys_tmp4562;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h11d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_73 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_73 <= w_sys_tmp4639;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h11d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_74 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_74 <= w_sys_tmp4640;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h123: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_75 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_75 <= w_sys_tmp4735;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h123: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_76 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_76 <= w_sys_tmp4736;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h129: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_77 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_77 <= w_sys_tmp4831;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h129: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_78 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_78 <= w_sys_tmp4832;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h7: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub09_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub09_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp830[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub09_u_datain <= w_sys_tmp833;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub09_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub09_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp1524[12:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp1527[12:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp1530[12:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp1536[12:0] );

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h57)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp2138[12:0] );

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp2132[12:0] );

									end
									else
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h3e) || (r_sys_run_step==7'h4b) || (r_sys_run_step==7'h58)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp2148[12:0] );

									end
									else
									if((r_sys_run_step==7'hb) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h3f) || (r_sys_run_step==7'h4c) || (r_sys_run_step==7'h59)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp2158[12:0] );

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4268[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sub09_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub09_result_datain <= w_sys_tmp1532;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h3e) || (r_sys_run_step==7'h4b) || (r_sys_run_step==7'h58)) begin
										r_sub09_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h57)) begin
										r_sub09_result_datain <= w_sys_tmp2111;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h7)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h6)) begin
										r_sub09_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h3f) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4c) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h59)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h3e) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h4b) || (r_sys_run_step==7'h57) || (r_sys_run_step==7'h58)) begin
										r_sub09_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub09_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub08_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub08_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp753[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub08_u_datain <= w_sys_tmp756;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub08_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub08_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1524[12:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1533[12:0] );

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h3a)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1643[12:0] );

									end
									else
									if((r_sys_run_step==7'hb) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h2b) || (r_sys_run_step==7'h33) || (r_sys_run_step==7'h3b)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1657[12:0] );

									end
									else
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h39)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1633[12:0] );

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h34)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1628[12:0] );

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4191[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub08_result_datain <= w_sys_tmp1526;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h3a)) begin
										r_sub08_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h39)) begin
										r_sub08_result_datain <= w_sys_tmp1608;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub08_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h2b) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h33) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h3b)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h3a)) begin
										r_sub08_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub08_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h10: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub12_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub12_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp1099[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub12_u_datain <= w_sys_tmp1102;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub12_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub12_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp1564[12:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp1573[12:0] );

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h36)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp1647[12:0] );

									end
									else
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h3d)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp1652[12:0] );

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp4559[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub12_result_datain <= w_sys_tmp1566;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h3d)) begin
										r_sub12_result_datain <= w_sys_tmp1656;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub12_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h36)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h3d)) begin
										r_sub12_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub12_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h3: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp316[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub03_u_datain <= w_sys_tmp319;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub03_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub03_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1450[12:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1447[12:0] );

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h50)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp3001[12:0] );

									end
									else
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h51)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp3012[12:0] );

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp3724[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sub03_result_datain <= w_sys_tmp1474;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h50)) begin
										r_sub03_result_datain <= w_sys_tmp3005;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_sub03_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h51)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h50)) begin
										r_sub03_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub03_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h2: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp227[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub02_u_datain <= w_sys_tmp230;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub02_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub02_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hb)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1444[12:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1456[12:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1450[12:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1447[12:0] );

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h50)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2554[12:0] );

									end
									else
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h51)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2565[12:0] );

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3628[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sub02_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub02_result_datain <= w_sys_tmp1446;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h50)) begin
										r_sub02_result_datain <= w_sys_tmp2558;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hb)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'ha)) begin
										r_sub02_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h51)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h50)) begin
										r_sub02_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub02_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h9: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub11_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub11_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1008[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub11_u_datain <= w_sys_tmp1011;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub11_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub11_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp1527[12:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp1530[12:0] );

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hb) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h3f) || (r_sys_run_step==7'h4c) || (r_sys_run_step==7'h59)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp3052[12:0] );

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp3026[12:0] );

									end
									else
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h57)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp3032[12:0] );

									end
									else
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h3e) || (r_sys_run_step==7'h4b) || (r_sys_run_step==7'h58)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp3042[12:0] );

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp4460[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sub11_result_datain <= w_sys_tmp1554;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h3e) || (r_sys_run_step==7'h4b) || (r_sys_run_step==7'h58)) begin
										r_sub11_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h57)) begin
										r_sub11_result_datain <= w_sys_tmp3005;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_sub11_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h3f) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4c) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h59)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h3e) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h4b) || (r_sys_run_step==7'h57) || (r_sys_run_step==7'h58)) begin
										r_sub11_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub11_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'hb: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub14_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub14_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp1265[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub14_u_datain <= w_sys_tmp1268;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub14_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub14_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp1576[12:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp1595[12:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp1567[12:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp1570[12:0] );

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h5b)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp2605[12:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp2599[12:0] );

									end
									else
									if((r_sys_run_step==7'he) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h42) || (r_sys_run_step==7'h4f)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp2595[12:0] );

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp4732[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sub14_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub14_result_datain <= w_sys_tmp1566;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h5b)) begin
										r_sub14_result_datain <= w_sys_tmp2609;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hb)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'ha)) begin
										r_sub14_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h42) || (r_sys_run_step==7'h4f)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h5b)) begin
										r_sub14_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub14_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp138[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub01_u_datain <= w_sys_tmp141;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub01_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub01_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1444[12:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1456[12:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1450[12:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1447[12:0] );

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h50)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2107[12:0] );

									end
									else
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h51)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2118[12:0] );

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3532[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sub01_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub01_result_datain <= w_sys_tmp1452;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h50)) begin
										r_sub01_result_datain <= w_sys_tmp2111;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h7)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h6)) begin
										r_sub01_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h51)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h50)) begin
										r_sub01_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'ha: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub13_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub13_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp1176[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub13_u_datain <= w_sys_tmp1179;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub13_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub13_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp1576[12:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp1567[12:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp1564[12:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp1570[12:0] );

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'he) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h42) || (r_sys_run_step==7'h4f)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp2148[12:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp2152[12:0] );

									end
									else
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h5b)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp2158[12:0] );

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp4636[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sub13_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub13_result_datain <= w_sys_tmp1572;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h5b)) begin
										r_sub13_result_datain <= w_sys_tmp2162;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h7)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h6)) begin
										r_sub13_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h42) || (r_sys_run_step==7'h4f)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h5b)) begin
										r_sub13_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub13_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp61[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub00_u_datain <= w_sys_tmp64;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub00_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub00_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1444[12:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1453[12:0] );

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h2b) || (r_sys_run_step==7'h33)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1619[12:0] );

									end
									else
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h32)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1604[12:0] );

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3455[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub00_result_datain <= w_sys_tmp1446;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h32)) begin
										r_sub00_result_datain <= w_sys_tmp1608;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub00_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h2b) || (r_sys_run_step==7'h33)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h32)) begin
										r_sub00_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h6: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub07_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub07_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp662[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub07_u_datain <= w_sys_tmp665;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub07_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub07_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1490[12:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1487[12:0] );

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h46) || (r_sys_run_step==7'h53)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp3012[12:0] );

									end
									else
									if((r_sys_run_step==7'h7) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h3b) || (r_sys_run_step==7'h48) || (r_sys_run_step==7'h55)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp3032[12:0] );

									end
									else
									if((r_sys_run_step==7'h6) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h47) || (r_sys_run_step==7'h54)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp3022[12:0] );

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp3006[12:0] );

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4092[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sub07_result_datain <= w_sys_tmp1514;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h46) || (r_sys_run_step==7'h53)) begin
										r_sub07_result_datain <= w_sys_tmp3016;

									end
									else
									if((r_sys_run_step==7'h6) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h47) || (r_sys_run_step==7'h54)) begin
										r_sub07_result_datain <= r_sys_tmp0_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_sub07_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h3b) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h48) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h55)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h46) || (r_sys_run_step==7'h47) || (r_sys_run_step==7'h53) || (r_sys_run_step==7'h54)) begin
										r_sub07_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub07_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h5: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub06_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub06_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp573[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub06_u_datain <= w_sys_tmp576;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub06_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub06_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1490[12:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1487[12:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1484[12:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1496[12:0] );

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2559[12:0] );

									end
									else
									if((r_sys_run_step==7'h6) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h47) || (r_sys_run_step==7'h54)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2575[12:0] );

									end
									else
									if((r_sys_run_step==7'h7) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h3b) || (r_sys_run_step==7'h48) || (r_sys_run_step==7'h55)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2585[12:0] );

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h46) || (r_sys_run_step==7'h53)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2565[12:0] );

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp3996[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sub06_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub06_result_datain <= w_sys_tmp1486;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h46) || (r_sys_run_step==7'h53)) begin
										r_sub06_result_datain <= w_sys_tmp2569;

									end
									else
									if((r_sys_run_step==7'h6) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h47) || (r_sys_run_step==7'h54)) begin
										r_sub06_result_datain <= r_sys_tmp0_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hb)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'ha)) begin
										r_sub06_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h3b) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h48) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h55)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h46) || (r_sys_run_step==7'h47) || (r_sys_run_step==7'h53) || (r_sys_run_step==7'h54)) begin
										r_sub06_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub06_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'hc: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub15_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub15_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp1354[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub15_u_datain <= w_sys_tmp1357;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub15_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub15_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp1567[12:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp1570[12:0] );

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h5b)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp3052[12:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp3046[12:0] );

									end
									else
									if((r_sys_run_step==7'he) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h42) || (r_sys_run_step==7'h4f)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp3042[12:0] );

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp4828[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sub15_result_datain <= w_sys_tmp1594;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h5b)) begin
										r_sub15_result_datain <= w_sys_tmp3056;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_sub15_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h42) || (r_sys_run_step==7'h4f)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h5b)) begin
										r_sub15_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub15_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h4: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub05_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub05_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp484[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub05_u_datain <= w_sys_tmp487;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub05_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub05_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1490[12:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1487[12:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1484[12:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1496[12:0] );

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2112[12:0] );

									end
									else
									if((r_sys_run_step==7'h7) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h3b) || (r_sys_run_step==7'h48) || (r_sys_run_step==7'h55)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2138[12:0] );

									end
									else
									if((r_sys_run_step==7'h6) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h47) || (r_sys_run_step==7'h54)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2128[12:0] );

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h46) || (r_sys_run_step==7'h53)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2118[12:0] );

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp3900[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sub05_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub05_result_datain <= w_sys_tmp1492;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h47) || (r_sys_run_step==7'h54)) begin
										r_sub05_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h46) || (r_sys_run_step==7'h53)) begin
										r_sub05_result_datain <= w_sys_tmp2122;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h7)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h6)) begin
										r_sub05_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h3b) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h48) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h55)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h46) || (r_sys_run_step==7'h47) || (r_sys_run_step==7'h53) || (r_sys_run_step==7'h54)) begin
										r_sub05_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub05_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'he: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub04_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub04_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp407[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub04_u_datain <= w_sys_tmp410;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub04_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub04_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1493[12:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1484[12:0] );

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h7) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h2f) || (r_sys_run_step==7'h37)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1638[12:0] );

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h35)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1614[12:0] );

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h30)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1609[12:0] );

									end
									else
									if((r_sys_run_step==7'h6) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h36)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1624[12:0] );

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp3823[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub04_result_datain <= w_sys_tmp1486;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sub04_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h35)) begin
										r_sub04_result_datain <= w_sys_tmp1618;

									end
									else
									if((r_sys_run_step==7'he) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h36)) begin
										r_sub04_result_datain <= w_sys_tmp1656;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub04_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h2f) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h37)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h36)) begin
										r_sub04_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub04_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub10_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub10_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp919[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub10_u_datain <= w_sys_tmp922;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub10_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub10_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hb)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp1524[12:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp1527[12:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp1530[12:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp1536[12:0] );

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hb) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h3f) || (r_sys_run_step==7'h4c) || (r_sys_run_step==7'h59)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp2605[12:0] );

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp2579[12:0] );

									end
									else
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h3e) || (r_sys_run_step==7'h4b) || (r_sys_run_step==7'h58)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp2595[12:0] );

									end
									else
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h57)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp2585[12:0] );

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp4364[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sub10_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub10_result_datain <= w_sys_tmp1526;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h3e) || (r_sys_run_step==7'h4b) || (r_sys_run_step==7'h58)) begin
										r_sub10_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h57)) begin
										r_sub10_result_datain <= w_sys_tmp2558;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hb)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'ha)) begin
										r_sub10_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h3f) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4c) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h59)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h3e) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h4b) || (r_sys_run_step==7'h57) || (r_sys_run_step==7'h58)) begin
										r_sub10_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub10_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp0_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp0_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp0_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp0_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp0_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h50)) begin
										r_sys_tmp0_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h50)) begin
										r_sys_tmp0_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h50)) begin
										r_sys_tmp0_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp1_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp1_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp1_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp1_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h38)) begin
										r_sys_tmp1_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h51)) begin
										r_sys_tmp1_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h51)) begin
										r_sys_tmp1_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h51)) begin
										r_sys_tmp1_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
