/*
TimeStamp:	2017/1/23		13:27
*/


module c1(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy,	
	output signed  [31:0] o_run_return,

	
	//subup
	input                 w_sub00_run_busy,
	output                r_sub00_run_req,
    output  signed [31:0] w_sub00_u_addr,
    output         [31:0] w_sub00_u_datain,
    input          [31:0] w_sub00_u_dataout,
    output                w_sub00_u_r_w,
    output  signed [31:0] w_sub00_result_addr,
    output         [31:0] w_sub00_result_datain,
    input          [31:0] w_sub00_result_dataout,
    output                w_sub00_result_r_w,
     
    
    //subunder
    input                 w_sub01_run_busy,
    output                r_sub01_run_req,
    output  signed [31:0] w_sub01_u_addr,
    output         [31:0] w_sub01_u_datain,
    input          [31:0] w_sub01_u_dataout,
    output                w_sub01_u_r_w,
    output  signed [31:0] w_sub01_result_addr,
    output         [31:0] w_sub01_result_datain,
    input          [31:0] w_sub01_result_dataout,
output w_sub01_result_r_w	
);

	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [31:0] r_sys_run_return;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 6:0] r_sys_run_phase;
	reg         [ 1:0] r_sys_run_stage;
	reg         [ 3:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 1:0] w_sys_run_stage_p1;
	wire        [ 3:0] w_sys_run_step_p1;
	wire signed [14:0] w_fld_u_0_addr_0;
	wire        [31:0] w_fld_u_0_datain_0;
	wire        [31:0] w_fld_u_0_dataout_0;
	wire               w_fld_u_0_r_w_0;
	wire               w_fld_u_0_ce_0;
	reg  signed [14:0] r_fld_u_0_addr_1;
	reg         [31:0] r_fld_u_0_datain_1;
	wire        [31:0] w_fld_u_0_dataout_1;
	reg                r_fld_u_0_r_w_1;
	wire               w_fld_u_0_ce_1;
	reg  signed [31:0] r_run_k_3;
	reg  signed [31:0] r_run_j_4;
	reg  signed [31:0] r_run_n_5;
	reg  signed [31:0] r_run_mx_6;
	reg  signed [31:0] r_run_my_7;
	reg  signed [31:0] r_run_nlast_8;
	reg         [31:0] r_run_dx_9;
	reg         [31:0] r_run_dy_10;
	reg         [31:0] r_run_r1_11;
	reg         [31:0] r_run_r2_12;
	reg         [31:0] r_run_dt_13;
	reg  signed [31:0] r_run_copy0_j_14;
	reg  signed [31:0] r_run_copy0_j_15;
	reg  signed [31:0] r_run_copy0_j_16;
	reg  signed [31:0] r_run_copy0_j_17;
	reg  signed [31:0] r_run_copy0_j_18;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [13:0] w_sub01_u_addr;
	reg  signed [13:0] r_sub01_u_addr;
	wire        [31:0] w_sub01_u_datain;
	reg         [31:0] r_sub01_u_datain;
	wire        [31:0] w_sub01_u_dataout;
	wire               w_sub01_u_r_w;
	reg                r_sub01_u_r_w;
	wire signed [13:0] w_sub01_result_addr;
	reg  signed [13:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [13:0] w_sub00_u_addr;
	reg  signed [13:0] r_sub00_u_addr;
	wire        [31:0] w_sub00_u_datain;
	reg         [31:0] r_sub00_u_datain;
	wire        [31:0] w_sub00_u_dataout;
	wire               w_sub00_u_r_w;
	reg                r_sub00_u_r_w;
	wire signed [13:0] w_sub00_result_addr;
	reg  signed [13:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	reg  signed [31:0] r_sys_tmp0_int;
	reg  signed [31:0] r_sys_tmp1_int;
	reg  signed [31:0] r_sys_tmp2_int;
	reg  signed [31:0] r_sys_tmp3_int;
	reg  signed [31:0] r_sys_tmp4_int;
	reg  signed [31:0] r_sys_tmp5_int;
	reg  signed [31:0] r_sys_tmp6_int;
	reg  signed [31:0] r_sys_tmp7_int;
	reg         [31:0] r_sys_tmp0_float;
	wire signed [31:0] w_sys_tmp1;
	wire        [31:0] w_sys_tmp3;
	wire        [31:0] w_sys_tmp5;
	wire        [31:0] w_sys_tmp6;
	wire               w_sys_tmp8;
	wire               w_sys_tmp9;
	wire signed [31:0] w_sys_tmp10;
	wire               w_sys_tmp11;
	wire               w_sys_tmp12;
	wire signed [31:0] w_sys_tmp15;
	wire signed [31:0] w_sys_tmp16;
	wire signed [31:0] w_sys_tmp17;
	wire        [31:0] w_sys_tmp18;
	wire signed [31:0] w_sys_tmp19;
	wire signed [31:0] w_sys_tmp21;
	wire signed [31:0] w_sys_tmp22;
	wire               w_sys_tmp56;
	wire               w_sys_tmp57;
	wire signed [31:0] w_sys_tmp58;
	wire signed [31:0] w_sys_tmp61;
	wire signed [31:0] w_sys_tmp62;
	wire        [31:0] w_sys_tmp63;
	wire signed [31:0] w_sys_tmp65;
	wire        [31:0] w_sys_tmp66;
	wire signed [31:0] w_sys_tmp67;
	wire               w_sys_tmp68;
	wire               w_sys_tmp69;
	wire signed [31:0] w_sys_tmp70;
	wire signed [31:0] w_sys_tmp73;
	wire signed [31:0] w_sys_tmp74;
	wire signed [31:0] w_sys_tmp75;
	wire        [31:0] w_sys_tmp76;
	wire signed [31:0] w_sys_tmp78;
	wire        [31:0] w_sys_tmp81;
	wire signed [31:0] w_sys_tmp82;
	wire signed [31:0] w_sys_tmp83;
	wire signed [31:0] w_sys_tmp85;
	wire signed [31:0] w_sys_tmp86;
	wire signed [31:0] w_sys_tmp90;
	wire signed [31:0] w_sys_tmp91;
	wire               w_sys_tmp162;
	wire               w_sys_tmp163;
	wire signed [31:0] w_sys_tmp164;
	wire signed [31:0] w_sys_tmp165;
	wire               w_sys_tmp166;
	wire               w_sys_tmp167;
	wire signed [31:0] w_sys_tmp168;
	wire signed [31:0] w_sys_tmp171;
	wire signed [31:0] w_sys_tmp172;
	wire        [31:0] w_sys_tmp173;
	wire signed [31:0] w_sys_tmp174;
	wire signed [31:0] w_sys_tmp175;
	wire signed [31:0] w_sys_tmp177;
	wire signed [31:0] w_sys_tmp178;
	wire signed [31:0] w_sys_tmp180;
	wire signed [31:0] w_sys_tmp181;
	wire signed [31:0] w_sys_tmp184;
	wire signed [31:0] w_sys_tmp185;
	wire signed [31:0] w_sys_tmp239;
	wire               w_sys_tmp240;
	wire               w_sys_tmp241;
	wire signed [31:0] w_sys_tmp242;
	wire signed [31:0] w_sys_tmp245;
	wire signed [31:0] w_sys_tmp246;
	wire signed [31:0] w_sys_tmp247;
	wire signed [31:0] w_sys_tmp248;
	wire        [31:0] w_sys_tmp249;
	wire signed [31:0] w_sys_tmp250;
	wire signed [31:0] w_sys_tmp251;
	wire signed [31:0] w_sys_tmp253;
	wire signed [31:0] w_sys_tmp254;
	wire signed [31:0] w_sys_tmp256;
	wire signed [31:0] w_sys_tmp257;
	wire signed [31:0] w_sys_tmp258;
	wire signed [31:0] w_sys_tmp262;
	wire signed [31:0] w_sys_tmp263;
	wire               w_sys_tmp327;
	wire               w_sys_tmp328;
	wire signed [31:0] w_sys_tmp329;
	wire signed [31:0] w_sys_tmp330;
	wire               w_sys_tmp331;
	wire               w_sys_tmp332;
	wire signed [31:0] w_sys_tmp333;
	wire signed [31:0] w_sys_tmp334;
	wire signed [31:0] w_sys_tmp335;
	wire               w_sys_tmp336;
	wire               w_sys_tmp337;
	wire signed [31:0] w_sys_tmp338;
	wire signed [31:0] w_sys_tmp341;
	wire signed [31:0] w_sys_tmp342;
	wire        [31:0] w_sys_tmp343;
	wire signed [31:0] w_sys_tmp344;
	wire signed [31:0] w_sys_tmp345;
	wire signed [31:0] w_sys_tmp347;
	wire signed [31:0] w_sys_tmp348;
	wire signed [31:0] w_sys_tmp350;
	wire signed [31:0] w_sys_tmp351;
	wire signed [31:0] w_sys_tmp354;
	wire signed [31:0] w_sys_tmp355;
	wire signed [31:0] w_sys_tmp409;
	wire               w_sys_tmp410;
	wire               w_sys_tmp411;
	wire signed [31:0] w_sys_tmp412;
	wire signed [31:0] w_sys_tmp415;
	wire signed [31:0] w_sys_tmp416;
	wire        [31:0] w_sys_tmp417;
	wire signed [31:0] w_sys_tmp418;
	wire signed [31:0] w_sys_tmp419;
	wire signed [31:0] w_sys_tmp420;
	wire signed [31:0] w_sys_tmp421;
	wire signed [31:0] w_sys_tmp423;
	wire signed [31:0] w_sys_tmp424;
	wire signed [31:0] w_sys_tmp426;
	wire signed [31:0] w_sys_tmp427;
	wire signed [31:0] w_sys_tmp430;
	wire signed [31:0] w_sys_tmp431;
	wire signed [31:0] w_sys_tmp432;
	wire        [31:0] w_sys_tmp497;
	wire signed [31:0] w_sys_tmp498;
	wire signed [31:0] w_sys_tmp499;
	wire signed [31:0] w_sys_tmp505;
	wire signed [31:0] w_sys_tmp506;
	wire signed [31:0] w_sys_tmp507;
	wire signed [31:0] w_sys_tmp508;
	wire signed [31:0] w_sys_tmp519;
	wire signed [31:0] w_sys_tmp520;
	wire signed [31:0] w_sys_tmp521;
	wire signed [31:0] w_sys_tmp532;
	wire signed [31:0] w_sys_tmp533;
	wire signed [31:0] w_sys_tmp534;
	wire signed [31:0] w_sys_tmp545;
	wire signed [31:0] w_sys_tmp546;
	wire signed [31:0] w_sys_tmp547;
	wire signed [31:0] w_sys_tmp558;
	wire signed [31:0] w_sys_tmp559;
	wire signed [31:0] w_sys_tmp560;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign o_run_return = r_sys_run_return;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 2'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 4'h1);
	assign w_fld_u_0_addr_0 = 15'sh0;
	assign w_fld_u_0_datain_0 = 32'h0;
	assign w_fld_u_0_r_w_0 = 1'h0;
	assign w_fld_u_0_ce_0 = w_sys_ce;
	assign w_fld_u_0_ce_1 = w_sys_ce;
	assign w_sub01_u_addr = ( (|r_sys_processing_methodID) ? r_sub01_u_addr : 14'sh0 ) ;
	assign w_sub01_u_datain = ( (|r_sys_processing_methodID) ? r_sub01_u_datain : 32'h0 ) ;
	assign w_sub01_u_r_w = ( (|r_sys_processing_methodID) ? r_sub01_u_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 14'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub00_u_addr = ( (|r_sys_processing_methodID) ? r_sub00_u_addr : 14'sh0 ) ;
	assign w_sub00_u_datain = ( (|r_sys_processing_methodID) ? r_sub00_u_datain : 32'h0 ) ;
	assign w_sub00_u_r_w = ( (|r_sys_processing_methodID) ? r_sub00_u_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 14'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh00000081;
	assign w_sys_tmp3 = 32'h3c000000;
	assign w_sys_tmp5 = 32'h3ba3d70a;
	assign w_sys_tmp6 = 32'h42a3d70a;
	assign w_sys_tmp8 = ( !w_sys_tmp9 );
	assign w_sys_tmp9 = (r_run_my_7 < r_run_k_3);
	assign w_sys_tmp10 = (r_run_k_3 + w_sys_intOne);
	assign w_sys_tmp11 = ( !w_sys_tmp12 );
	assign w_sys_tmp12 = (r_run_mx_6 < r_run_j_4);
	assign w_sys_tmp15 = (w_sys_tmp16 + r_run_k_3);
	assign w_sys_tmp16 = (r_run_j_4 * w_sys_tmp17);
	assign w_sys_tmp17 = 32'sh00000081;
	assign w_sys_tmp18 = 32'h0;
	assign w_sys_tmp19 = (r_run_j_4 + w_sys_intOne);
	assign w_sys_tmp21 = (w_sys_tmp22 * w_sys_tmp17);
	assign w_sys_tmp22 = w_sys_tmp19;
	assign w_sys_tmp56 = ( !w_sys_tmp57 );
	assign w_sys_tmp57 = (w_sys_tmp58 < r_run_k_3);
	assign w_sys_tmp58 = 32'sh00000081;
	assign w_sys_tmp61 = (w_sys_tmp62 + r_run_k_3);
	assign w_sys_tmp62 = 32'sh00000081;
	assign w_sys_tmp63 = 32'h3f000000;
	assign w_sys_tmp65 = 32'sh00004101;
	assign w_sys_tmp66 = 32'h0;
	assign w_sys_tmp67 = (r_run_k_3 + w_sys_intOne);
	assign w_sys_tmp68 = ( !w_sys_tmp69 );
	assign w_sys_tmp69 = (w_sys_tmp70 < r_run_j_4);
	assign w_sys_tmp70 = 32'sh00000081;
	assign w_sys_tmp73 = (w_sys_tmp74 + w_sys_intOne);
	assign w_sys_tmp74 = (r_run_j_4 * w_sys_tmp75);
	assign w_sys_tmp75 = 32'sh00000081;
	assign w_sys_tmp76 = 32'h3f800000;
	assign w_sys_tmp78 = (r_run_copy0_j_14 * w_sys_tmp75);
	assign w_sys_tmp81 = 32'h0;
	assign w_sys_tmp82 = (r_run_copy0_j_14 + w_sys_intOne);
	assign w_sys_tmp83 = (r_run_j_4 + w_sys_intOne);
	assign w_sys_tmp85 = (w_sys_tmp86 * w_sys_tmp75);
	assign w_sys_tmp86 = w_sys_tmp83;
	assign w_sys_tmp90 = (w_sys_tmp91 * w_sys_tmp75);
	assign w_sys_tmp91 = w_sys_tmp82;
	assign w_sys_tmp162 = ( !w_sys_tmp163 );
	assign w_sys_tmp163 = (w_sys_tmp164 < r_run_k_3);
	assign w_sys_tmp164 = 32'sh00000081;
	assign w_sys_tmp165 = (r_run_k_3 + w_sys_intOne);
	assign w_sys_tmp166 = ( !w_sys_tmp167 );
	assign w_sys_tmp167 = (w_sys_tmp168 < r_run_j_4);
	assign w_sys_tmp168 = 32'sh00000041;
	assign w_sys_tmp171 = (r_run_j_4 * w_sys_tmp172);
	assign w_sys_tmp172 = 32'sh00000081;
	assign w_sys_tmp173 = w_fld_u_0_dataout_1;
	assign w_sys_tmp174 = (w_sys_tmp175 + r_run_k_3);
	assign w_sys_tmp175 = (r_run_copy0_j_15 * w_sys_tmp172);
	assign w_sys_tmp177 = (r_run_copy0_j_15 + w_sys_intOne);
	assign w_sys_tmp178 = (r_run_j_4 + w_sys_intOne);
	assign w_sys_tmp180 = (w_sys_tmp181 * w_sys_tmp172);
	assign w_sys_tmp181 = w_sys_tmp178;
	assign w_sys_tmp184 = (w_sys_tmp185 * w_sys_tmp172);
	assign w_sys_tmp185 = w_sys_tmp177;
	assign w_sys_tmp239 = 32'sh00000040;
	assign w_sys_tmp240 = ( !w_sys_tmp241 );
	assign w_sys_tmp241 = (w_sys_tmp242 < r_run_j_4);
	assign w_sys_tmp242 = 32'sh00000081;
	assign w_sys_tmp245 = (w_sys_tmp246 * w_sys_tmp248);
	assign w_sys_tmp246 = (r_run_j_4 - w_sys_tmp247);
	assign w_sys_tmp247 = 32'sh0000003f;
	assign w_sys_tmp248 = 32'sh00000081;
	assign w_sys_tmp249 = w_fld_u_0_dataout_1;
	assign w_sys_tmp250 = (w_sys_tmp251 + r_run_k_3);
	assign w_sys_tmp251 = (r_run_copy0_j_16 * w_sys_tmp248);
	assign w_sys_tmp253 = (r_run_copy0_j_16 + w_sys_intOne);
	assign w_sys_tmp254 = (r_run_j_4 + w_sys_intOne);
	assign w_sys_tmp256 = (w_sys_tmp257 * w_sys_tmp248);
	assign w_sys_tmp257 = (w_sys_tmp258 - w_sys_tmp247);
	assign w_sys_tmp258 = w_sys_tmp254;
	assign w_sys_tmp262 = (w_sys_tmp263 * w_sys_tmp248);
	assign w_sys_tmp263 = w_sys_tmp253;
	assign w_sys_tmp327 = ( !w_sys_tmp328 );
	assign w_sys_tmp328 = (r_run_nlast_8 < r_run_n_5);
	assign w_sys_tmp329 = (r_run_n_5 + w_sys_intOne);
	assign w_sys_tmp330 = 32'sh00000002;
	assign w_sys_tmp331 = ( !w_sys_tmp332 );
	assign w_sys_tmp332 = (w_sys_tmp333 < r_run_k_3);
	assign w_sys_tmp333 = 32'sh00000080;
	assign w_sys_tmp334 = (r_run_k_3 + w_sys_intOne);
	assign w_sys_tmp335 = 32'sh00000002;
	assign w_sys_tmp336 = ( !w_sys_tmp337 );
	assign w_sys_tmp337 = (w_sys_tmp338 < r_run_j_4);
	assign w_sys_tmp338 = 32'sh00000040;
	assign w_sys_tmp341 = (r_run_j_4 * w_sys_tmp342);
	assign w_sys_tmp342 = 32'sh00000081;
	assign w_sys_tmp343 = w_sub00_result_dataout;
	assign w_sys_tmp344 = (w_sys_tmp345 + r_run_k_3);
	assign w_sys_tmp345 = (r_run_copy0_j_17 * w_sys_tmp342);
	assign w_sys_tmp347 = (r_run_copy0_j_17 + w_sys_intOne);
	assign w_sys_tmp348 = (r_run_j_4 + w_sys_intOne);
	assign w_sys_tmp350 = (w_sys_tmp351 * w_sys_tmp342);
	assign w_sys_tmp351 = w_sys_tmp348;
	assign w_sys_tmp354 = (w_sys_tmp355 * w_sys_tmp342);
	assign w_sys_tmp355 = w_sys_tmp347;
	assign w_sys_tmp409 = 32'sh00000041;
	assign w_sys_tmp410 = ( !w_sys_tmp411 );
	assign w_sys_tmp411 = (w_sys_tmp412 < r_run_j_4);
	assign w_sys_tmp412 = 32'sh00000080;
	assign w_sys_tmp415 = (r_run_j_4 * w_sys_tmp416);
	assign w_sys_tmp416 = 32'sh00000081;
	assign w_sys_tmp417 = w_sub01_result_dataout;
	assign w_sys_tmp418 = (w_sys_tmp419 + r_run_k_3);
	assign w_sys_tmp419 = (w_sys_tmp420 * w_sys_tmp416);
	assign w_sys_tmp420 = (r_run_copy0_j_18 - w_sys_tmp421);
	assign w_sys_tmp421 = 32'sh0000003f;
	assign w_sys_tmp423 = (r_run_copy0_j_18 + w_sys_intOne);
	assign w_sys_tmp424 = (r_run_j_4 + w_sys_intOne);
	assign w_sys_tmp426 = (w_sys_tmp427 * w_sys_tmp416);
	assign w_sys_tmp427 = w_sys_tmp424;
	assign w_sys_tmp430 = (w_sys_tmp431 * w_sys_tmp416);
	assign w_sys_tmp431 = (w_sys_tmp432 - w_sys_tmp421);
	assign w_sys_tmp432 = w_sys_tmp423;
	assign w_sys_tmp497 = w_fld_u_0_dataout_1;
	assign w_sys_tmp498 = 32'sh00000104;
	assign w_sys_tmp499 = (w_sys_tmp21 + r_run_k_3);
	assign w_sys_tmp505 = (w_sys_tmp65 + r_run_k_3);
	assign w_sys_tmp506 = (w_sys_tmp78 + w_sys_tmp75);
	assign w_sys_tmp507 = (w_sys_tmp85 + w_sys_intOne);
	assign w_sys_tmp508 = (w_sys_tmp90 + w_sys_tmp75);
	assign w_sys_tmp519 = (w_sys_tmp171 + r_run_k_3);
	assign w_sys_tmp520 = (w_sys_tmp180 + r_run_k_3);
	assign w_sys_tmp521 = (w_sys_tmp184 + r_run_k_3);
	assign w_sys_tmp532 = (w_sys_tmp245 + r_run_k_3);
	assign w_sys_tmp533 = (w_sys_tmp256 + r_run_k_3);
	assign w_sys_tmp534 = (w_sys_tmp262 + r_run_k_3);
	assign w_sys_tmp545 = (w_sys_tmp341 + r_run_k_3);
	assign w_sys_tmp546 = (w_sys_tmp350 + r_run_k_3);
	assign w_sys_tmp547 = (w_sys_tmp354 + r_run_k_3);
	assign w_sys_tmp558 = (w_sys_tmp415 + r_run_k_3);
	assign w_sys_tmp559 = (w_sys_tmp426 + r_run_k_3);
	assign w_sys_tmp560 = (w_sys_tmp430 + r_run_k_3);

/*
	subunder
		sub01_inst(
			.i_fld_result_1_addr_0 (w_sub01_result_addr),
			.i_fld_result_1_datain_0 (w_sub01_result_datain),
			.o_fld_result_1_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub01_result_r_w),
			.i_fld_u_0_addr_0 (w_sub01_u_addr),
			.i_fld_u_0_datain_0 (w_sub01_u_datain),
			.o_fld_u_0_dataout_0 (w_sub01_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub01_u_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	subup
		sub00_inst(
			.i_fld_result_1_addr_0 (w_sub00_result_addr),
			.i_fld_result_1_datain_0 (w_sub00_result_datain),
			.o_fld_result_1_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub00_result_r_w),
			.i_fld_u_0_addr_0 (w_sub00_u_addr),
			.i_fld_u_0_datain_0 (w_sub00_u_datain),
			.o_fld_u_0_dataout_0 (w_sub00_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub00_u_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);
*/
	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_u_0(
			.clk (clock),
			.ce_0 (w_fld_u_0_ce_0),
			.addr_0 (w_fld_u_0_addr_0),
			.datain_0 (w_fld_u_0_datain_0),
			.dataout_0 (w_fld_u_0_dataout_0),
			.r_w_0 (w_fld_u_0_r_w_0),
			.ce_1 (w_fld_u_0_ce_1),
			.addr_1 (r_fld_u_0_addr_1),
			.datain_1 (r_fld_u_0_datain_1),
			.dataout_1 (w_fld_u_0_dataout_1),
			.r_w_1 (r_fld_u_0_r_w_1)
		);

	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						7'h47: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_return <= 32'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h44: begin
							r_sys_run_return <= r_sys_tmp0_float;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 7'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h0: begin
							r_sys_run_phase <= 7'h2;
						end

						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h4;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h5;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp8) ? 7'h9 : 7'hf);

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h5;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'ha;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp11) ? 7'hd : 7'h6);

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h6)) begin
										r_sys_run_phase <= 7'ha;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h10;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp56) ? 7'h13 : 7'h15);

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h1)) begin
										r_sys_run_phase <= 7'h10;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h16;

									end
								end

							endcase
						end

						7'h16: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp68) ? 7'h19 : 7'h1b);

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'hd)) begin
										r_sys_run_phase <= 7'h16;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h1c;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp162) ? 7'h20 : 7'h2c);

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h1c;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h21;

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp166) ? 7'h24 : 7'h26);

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h8)) begin
										r_sys_run_phase <= 7'h21;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h27;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp240) ? 7'h2a : 7'h1d);

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h8)) begin
										r_sys_run_phase <= 7'h27;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h2d;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp327) ? 7'h30 : 7'h34);

									end
								end

							endcase
						end

						7'h2e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h2d;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==4'h1)) begin
										r_sys_run_phase <= 7'h32;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==4'h1)) begin
										r_sys_run_phase <= 7'h2e;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h35;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp331) ? 7'h39 : 7'h45);

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h35;

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h3a;

									end
								end

							endcase
						end

						7'h3a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp336) ? 7'h3d : 7'h3f);

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h8)) begin
										r_sys_run_phase <= 7'h3a;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h40;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp410) ? 7'h43 : 7'h36);

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h8)) begin
										r_sys_run_phase <= 7'h40;

									end
								end

							endcase
						end

						7'h44: begin
							r_sys_run_phase <= 7'h47;
						end

						7'h45: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h2)) begin
										r_sys_run_phase <= 7'h44;

									end
								end

							endcase
						end

						7'h47: begin
							r_sys_run_phase <= 7'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h6)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h1)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h16: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'hd)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h8)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h8)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h2e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h1)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h1)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h3a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h8)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h8)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h2)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 4'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h5)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==4'h6)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==4'h1)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h16: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'hc)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==4'hd)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==4'h8)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==4'h8)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h2e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==4'h1)) begin
										r_sys_run_step <= 4'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==4'h1)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= ((w_sub00_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==4'h1)) begin
										r_sys_run_step <= 4'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= ((w_sub01_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==4'h1)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h3a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==4'h8)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==4'h8)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0) || (r_sys_run_step==4'h1)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==4'h2)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						7'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						7'h47: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h1<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp0_int[14:0] );

									end
									else
									if((r_sys_run_step==4'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp15[14:0] );

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h1)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp0_int[14:0] );

									end
									else
									if((r_sys_run_step==4'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp61[14:0] );

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'hb)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp1_int[14:0] );

									end
									else
									if((r_sys_run_step==4'h8)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp2_int[14:0] );

									end
									else
									if((r_sys_run_step==4'hc)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp0_int[14:0] );

									end
									else
									if((r_sys_run_step==4'h2) || (r_sys_run_step==4'h6)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp5_int[14:0] );

									end
									else
									if((r_sys_run_step==4'h3) || (r_sys_run_step==4'h9)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp6_int[14:0] );

									end
									else
									if((r_sys_run_step==4'h1) || (r_sys_run_step==4'h5) || (r_sys_run_step==4'hd)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp7_int[14:0] );

									end
									else
									if((r_sys_run_step==4'h4) || (r_sys_run_step==4'ha)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp4_int[14:0] );

									end
									else
									if((r_sys_run_step==4'h7)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp3_int[14:0] );

									end
									else
									if((r_sys_run_step==4'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp73[14:0] );

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp174[14:0] );

									end
									else
									if((4'h1<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp4_int[14:0] );

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h1<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp2_int[14:0] );

									end
									else
									if((r_sys_run_step==4'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp250[14:0] );

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h2) || (r_sys_run_step==4'h5) || (r_sys_run_step==4'h8)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp5_int[14:0] );

									end
									else
									if((r_sys_run_step==4'h4) || (r_sys_run_step==4'h7)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp7_int[14:0] );

									end
									else
									if((r_sys_run_step==4'h3) || (r_sys_run_step==4'h6)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp3_int[14:0] );

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h3) || (r_sys_run_step==4'h6)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp1_int[14:0] );

									end
									else
									if((r_sys_run_step==4'h4) || (r_sys_run_step==4'h7)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp7_int[14:0] );

									end
									else
									if((r_sys_run_step==4'h2) || (r_sys_run_step==4'h5) || (r_sys_run_step==4'h8)) begin
										r_fld_u_0_addr_1 <= $signed( r_sys_tmp3_int[14:0] );

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp498[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp18;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp63;

									end
									else
									if((r_sys_run_step==4'h1)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp66;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h1) || (r_sys_run_step==4'h3) || (r_sys_run_step==4'h5) || (r_sys_run_step==4'h7) || (r_sys_run_step==4'h9) || (r_sys_run_step==4'hb) || (r_sys_run_step==4'hd)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp81;

									end
									else
									if((r_sys_run_step==4'h0) || (r_sys_run_step==4'h2) || (r_sys_run_step==4'h4) || (r_sys_run_step==4'h6) || (r_sys_run_step==4'h8) || (r_sys_run_step==4'ha) || (r_sys_run_step==4'hc)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp76;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h2<=r_sys_run_step && r_sys_run_step<=4'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp343;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h2<=r_sys_run_step && r_sys_run_step<=4'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp417;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0) || (r_sys_run_step==4'h1)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'hd)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h2<=r_sys_run_step && r_sys_run_step<=4'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h2<=r_sys_run_step && r_sys_run_step<=4'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h47: begin
							r_fld_u_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_k_3 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_k_3 <= w_sys_tmp10;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_k_3 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_k_3 <= w_sys_tmp67;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_k_3 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_k_3 <= w_sys_tmp165;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_k_3 <= w_sys_tmp330;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_k_3 <= w_sys_tmp334;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_j_4 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_run_j_4 <= w_sys_tmp19;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_j_4 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_run_j_4 <= w_sys_tmp83;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_j_4 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_run_j_4 <= w_sys_tmp178;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_j_4 <= w_sys_tmp239;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_run_j_4 <= w_sys_tmp254;

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_j_4 <= w_sys_tmp335;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_run_j_4 <= w_sys_tmp348;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_j_4 <= w_sys_tmp409;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_run_j_4 <= w_sys_tmp424;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_n_5 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h2e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_n_5 <= w_sys_tmp329;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_mx_6 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_my_7 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_nlast_8 <= w_sys_intOne;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_dx_9 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_dy_10 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_r1_11 <= w_sys_tmp6;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_r2_12 <= w_sys_tmp6;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_dt_13 <= w_sys_tmp5;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h15: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_copy0_j_14 <= r_run_j_4;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_run_copy0_j_14 <= w_sys_tmp82;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h20: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_copy0_j_15 <= r_run_j_4;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_run_copy0_j_15 <= w_sys_tmp177;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h26: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_copy0_j_16 <= r_run_j_4;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_run_copy0_j_16 <= w_sys_tmp253;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h39: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_copy0_j_17 <= r_run_j_4;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_run_copy0_j_17 <= w_sys_tmp347;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3f: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_copy0_j_18 <= r_run_j_4;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_run_copy0_j_18 <= w_sys_tmp423;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h30: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==4'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h2) || (r_sys_run_step==4'h5) || (r_sys_run_step==4'h8)) begin
										r_sub01_u_addr <= $signed( r_sys_tmp1_int[13:0] );

									end
									else
									if((r_sys_run_step==4'h4) || (r_sys_run_step==4'h7)) begin
										r_sub01_u_addr <= $signed( r_sys_tmp5_int[13:0] );

									end
									else
									if((r_sys_run_step==4'h3) || (r_sys_run_step==4'h6)) begin
										r_sub01_u_addr <= $signed( r_sys_tmp6_int[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h2<=r_sys_run_step && r_sys_run_step<=4'h8)) begin
										r_sub01_u_datain <= w_sys_tmp249;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h2<=r_sys_run_step && r_sys_run_step<=4'h8)) begin
										r_sub01_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h47: begin
							r_sub01_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h43: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp418[13:0] );

									end
									else
									if((4'h1<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_sub01_result_addr <= $signed( r_sys_tmp5_int[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h30: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h47: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h30: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==4'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h4) || (r_sys_run_step==4'h7)) begin
										r_sub00_u_addr <= $signed( r_sys_tmp1_int[13:0] );

									end
									else
									if((r_sys_run_step==4'h3) || (r_sys_run_step==4'h6)) begin
										r_sub00_u_addr <= $signed( r_sys_tmp2_int[13:0] );

									end
									else
									if((r_sys_run_step==4'h2) || (r_sys_run_step==4'h5) || (r_sys_run_step==4'h8)) begin
										r_sub00_u_addr <= $signed( r_sys_tmp3_int[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h2<=r_sys_run_step && r_sys_run_step<=4'h8)) begin
										r_sub00_u_datain <= w_sys_tmp173;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h2<=r_sys_run_step && r_sys_run_step<=4'h8)) begin
										r_sub00_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h47: begin
							r_sub00_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h1<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_sub00_result_addr <= $signed( r_sys_tmp6_int[13:0] );

									end
									else
									if((r_sys_run_step==4'h0)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp344[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h30: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h47: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h5)) begin
										r_sys_tmp0_int <= w_sys_tmp499;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_tmp0_int <= w_sys_tmp505;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h5)) begin
										r_sys_tmp0_int <= w_sys_tmp507;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h4)) begin
										r_sys_tmp1_int <= w_sys_tmp508;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h1) || (r_sys_run_step==4'h4)) begin
										r_sys_tmp1_int <= w_sys_tmp520;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_tmp1_int <= w_sys_tmp532;

									end
									else
									if((r_sys_run_step==4'h2) || (r_sys_run_step==4'h5)) begin
										r_sys_tmp1_int <= w_sys_tmp533;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0) || (r_sys_run_step==4'h3)) begin
										r_sys_tmp1_int <= w_sys_tmp559;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h3)) begin
										r_sys_tmp2_int <= w_sys_tmp507;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0) || (r_sys_run_step==4'h3)) begin
										r_sys_tmp2_int <= w_sys_tmp520;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h5)) begin
										r_sys_tmp2_int <= w_sys_tmp534;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h2)) begin
										r_sys_tmp3_int <= w_sys_tmp508;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_tmp3_int <= w_sys_tmp519;

									end
									else
									if((r_sys_run_step==4'h2) || (r_sys_run_step==4'h5)) begin
										r_sys_tmp3_int <= w_sys_tmp520;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0) || (r_sys_run_step==4'h3)) begin
										r_sys_tmp3_int <= w_sys_tmp546;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h2) || (r_sys_run_step==4'h5)) begin
										r_sys_tmp3_int <= w_sys_tmp559;

									end
									else
									if((r_sys_run_step==4'h0)) begin
										r_sys_tmp3_int <= w_sys_tmp558;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h1) || (r_sys_run_step==4'h4)) begin
										r_sys_tmp4_int <= w_sys_tmp507;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h5)) begin
										r_sys_tmp4_int <= w_sys_tmp521;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0) || (r_sys_run_step==4'h2)) begin
										r_sys_tmp5_int <= w_sys_tmp507;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h1) || (r_sys_run_step==4'h4)) begin
										r_sys_tmp5_int <= w_sys_tmp533;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h2) || (r_sys_run_step==4'h5)) begin
										r_sys_tmp5_int <= w_sys_tmp546;

									end
									else
									if((r_sys_run_step==4'h0)) begin
										r_sys_tmp5_int <= w_sys_tmp545;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h5)) begin
										r_sys_tmp5_int <= w_sys_tmp560;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0) || (r_sys_run_step==4'h3)) begin
										r_sys_tmp6_int <= w_sys_tmp508;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0) || (r_sys_run_step==4'h3)) begin
										r_sys_tmp6_int <= w_sys_tmp533;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h5)) begin
										r_sys_tmp6_int <= w_sys_tmp547;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h1) || (r_sys_run_step==4'h5)) begin
										r_sys_tmp7_int <= w_sys_tmp508;

									end
									else
									if((r_sys_run_step==4'h0)) begin
										r_sys_tmp7_int <= w_sys_tmp506;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h1) || (r_sys_run_step==4'h4)) begin
										r_sys_tmp7_int <= w_sys_tmp546;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h1) || (r_sys_run_step==4'h4)) begin
										r_sys_tmp7_int <= w_sys_tmp559;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h2)) begin
										r_sys_tmp0_float <= w_sys_tmp497;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
