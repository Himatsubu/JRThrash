/*
TimeStamp:	2016/4/26		14:59
*/


module c1(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy	
);

	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 5:0] r_sys_run_phase;
	reg         [ 2:0] r_sys_run_stage;
	reg         [ 8:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 2:0] w_sys_run_stage_p1;
	wire        [ 8:0] w_sys_run_step_p1;
	wire signed [ 8:0] w_fld_u_0_addr_0;
	wire        [31:0] w_fld_u_0_datain_0;
	wire        [31:0] w_fld_u_0_dataout_0;
	wire               w_fld_u_0_r_w_0;
	wire               w_fld_u_0_ce_0;
	reg  signed [ 8:0] r_fld_u_0_addr_1;
	reg         [31:0] r_fld_u_0_datain_1;
	wire        [31:0] w_fld_u_0_dataout_1;
	reg                r_fld_u_0_r_w_1;
	wire               w_fld_u_0_ce_1;
	wire signed [ 8:0] w_fld_uu_1_addr_0;
	wire        [31:0] w_fld_uu_1_datain_0;
	wire        [31:0] w_fld_uu_1_dataout_0;
	wire               w_fld_uu_1_r_w_0;
	wire               w_fld_uu_1_ce_0;
	reg  signed [ 8:0] r_fld_uu_1_addr_1;
	reg         [31:0] r_fld_uu_1_datain_1;
	wire        [31:0] w_fld_uu_1_dataout_1;
	reg                r_fld_uu_1_r_w_1;
	wire               w_fld_uu_1_ce_1;
	reg  signed [31:0] r_run_k_6;
	reg  signed [31:0] r_run_j_7;
	reg  signed [31:0] r_run_n_8;
	reg  signed [31:0] r_run_mx_9;
	reg  signed [31:0] r_run_my_10;
	reg  signed [31:0] r_run_nlast_11;
	reg         [31:0] r_run_dx_12;
	reg         [31:0] r_run_dy_13;
	reg  signed [31:0] r_run_copy0_j_14;
	reg  signed [31:0] r_run_copy0_j_15;
	reg  signed [31:0] r_run_copy1_j_16;
	reg  signed [31:0] r_run_copy2_j_17;
	reg                r_sub03_run_req;
	wire               w_sub03_run_busy;
	wire signed [ 8:0] w_sub03_u_addr;
	reg  signed [ 8:0] r_sub03_u_addr;
	wire        [31:0] w_sub03_u_datain;
	reg         [31:0] r_sub03_u_datain;
	wire        [31:0] w_sub03_u_dataout;
	wire               w_sub03_u_r_w;
	reg                r_sub03_u_r_w;
	wire signed [ 8:0] w_sub03_result_addr;
	reg  signed [ 8:0] r_sub03_result_addr;
	wire        [31:0] w_sub03_result_datain;
	reg         [31:0] r_sub03_result_datain;
	wire        [31:0] w_sub03_result_dataout;
	wire               w_sub03_result_r_w;
	reg                r_sub03_result_r_w;
	reg                r_sub02_run_req;
	wire               w_sub02_run_busy;
	wire signed [ 8:0] w_sub02_u_addr;
	reg  signed [ 8:0] r_sub02_u_addr;
	wire        [31:0] w_sub02_u_datain;
	reg         [31:0] r_sub02_u_datain;
	wire        [31:0] w_sub02_u_dataout;
	wire               w_sub02_u_r_w;
	reg                r_sub02_u_r_w;
	wire signed [ 8:0] w_sub02_result_addr;
	reg  signed [ 8:0] r_sub02_result_addr;
	wire        [31:0] w_sub02_result_datain;
	reg         [31:0] r_sub02_result_datain;
	wire        [31:0] w_sub02_result_dataout;
	wire               w_sub02_result_r_w;
	reg                r_sub02_result_r_w;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [ 8:0] w_sub01_u_addr;
	reg  signed [ 8:0] r_sub01_u_addr;
	wire        [31:0] w_sub01_u_datain;
	reg         [31:0] r_sub01_u_datain;
	wire        [31:0] w_sub01_u_dataout;
	wire               w_sub01_u_r_w;
	reg                r_sub01_u_r_w;
	wire signed [ 8:0] w_sub01_result_addr;
	reg  signed [ 8:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [ 8:0] w_sub00_u_addr;
	reg  signed [ 8:0] r_sub00_u_addr;
	wire        [31:0] w_sub00_u_datain;
	reg         [31:0] r_sub00_u_datain;
	wire        [31:0] w_sub00_u_dataout;
	wire               w_sub00_u_r_w;
	reg                r_sub00_u_r_w;
	wire signed [ 8:0] w_sub00_result_addr;
	reg  signed [ 8:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg         [31:0] r_sys_tmp4_float;
	reg         [31:0] r_sys_tmp5_float;
	reg         [31:0] r_sys_tmp6_float;
	reg         [31:0] r_sys_tmp7_float;
	reg         [31:0] r_sys_tmp8_float;
	wire signed [31:0] w_sys_tmp1;
	wire        [31:0] w_sys_tmp3;
	wire signed [31:0] w_sys_tmp5;
	wire               w_sys_tmp6;
	wire               w_sys_tmp7;
	wire signed [31:0] w_sys_tmp8;
	wire               w_sys_tmp9;
	wire               w_sys_tmp10;
	wire signed [31:0] w_sys_tmp13;
	wire signed [31:0] w_sys_tmp14;
	wire signed [31:0] w_sys_tmp15;
	wire        [31:0] w_sys_tmp16;
	wire signed [31:0] w_sys_tmp18;
	wire signed [31:0] w_sys_tmp19;
	wire signed [31:0] w_sys_tmp22;
	wire signed [31:0] w_sys_tmp23;
	wire               w_sys_tmp780;
	wire               w_sys_tmp781;
	wire signed [31:0] w_sys_tmp782;
	wire               w_sys_tmp783;
	wire               w_sys_tmp784;
	wire signed [31:0] w_sys_tmp787;
	wire signed [31:0] w_sys_tmp788;
	wire        [31:0] w_sys_tmp789;
	wire signed [31:0] w_sys_tmp791;
	wire signed [31:0] w_sys_tmp792;
	wire        [31:0] w_sys_tmp794;
	wire signed [31:0] w_sys_tmp796;
	wire signed [31:0] w_sys_tmp797;
	wire        [31:0] w_sys_tmp799;
	wire signed [31:0] w_sys_tmp801;
	wire signed [31:0] w_sys_tmp802;
	wire signed [31:0] w_sys_tmp805;
	wire signed [31:0] w_sys_tmp806;
	wire signed [31:0] w_sys_tmp807;
	wire signed [31:0] w_sys_tmp808;
	wire signed [31:0] w_sys_tmp2258;
	wire               w_sys_tmp2259;
	wire               w_sys_tmp2260;
	wire signed [31:0] w_sys_tmp2263;
	wire signed [31:0] w_sys_tmp2264;
	wire        [31:0] w_sys_tmp2265;
	wire signed [31:0] w_sys_tmp2269;
	wire signed [31:0] w_sys_tmp2270;
	wire signed [31:0] w_sys_tmp2275;
	wire signed [31:0] w_sys_tmp2276;
	wire signed [31:0] w_sys_tmp2281;
	wire signed [31:0] w_sys_tmp2282;
	wire signed [31:0] w_sys_tmp2287;
	wire signed [31:0] w_sys_tmp2288;
	wire signed [31:0] w_sys_tmp2293;
	wire signed [31:0] w_sys_tmp2294;
	wire signed [31:0] w_sys_tmp2299;
	wire signed [31:0] w_sys_tmp2300;
	wire signed [31:0] w_sys_tmp2305;
	wire signed [31:0] w_sys_tmp2306;
	wire signed [31:0] w_sys_tmp2311;
	wire signed [31:0] w_sys_tmp2312;
	wire signed [31:0] w_sys_tmp2317;
	wire signed [31:0] w_sys_tmp2318;
	wire signed [31:0] w_sys_tmp2323;
	wire signed [31:0] w_sys_tmp2324;
	wire signed [31:0] w_sys_tmp2329;
	wire signed [31:0] w_sys_tmp2330;
	wire signed [31:0] w_sys_tmp2335;
	wire signed [31:0] w_sys_tmp2336;
	wire signed [31:0] w_sys_tmp2341;
	wire signed [31:0] w_sys_tmp2342;
	wire signed [31:0] w_sys_tmp2347;
	wire signed [31:0] w_sys_tmp2348;
	wire signed [31:0] w_sys_tmp2353;
	wire signed [31:0] w_sys_tmp2354;
	wire signed [31:0] w_sys_tmp2359;
	wire signed [31:0] w_sys_tmp2360;
	wire signed [31:0] w_sys_tmp2365;
	wire signed [31:0] w_sys_tmp2366;
	wire signed [31:0] w_sys_tmp2371;
	wire signed [31:0] w_sys_tmp2372;
	wire signed [31:0] w_sys_tmp2377;
	wire signed [31:0] w_sys_tmp2378;
	wire signed [31:0] w_sys_tmp2383;
	wire signed [31:0] w_sys_tmp2384;
	wire signed [31:0] w_sys_tmp2400;
	wire               w_sys_tmp2401;
	wire               w_sys_tmp2402;
	wire signed [31:0] w_sys_tmp2403;
	wire signed [31:0] w_sys_tmp2406;
	wire signed [31:0] w_sys_tmp2407;
	wire        [31:0] w_sys_tmp2408;
	wire signed [31:0] w_sys_tmp2412;
	wire signed [31:0] w_sys_tmp2413;
	wire signed [31:0] w_sys_tmp2418;
	wire signed [31:0] w_sys_tmp2419;
	wire signed [31:0] w_sys_tmp2424;
	wire signed [31:0] w_sys_tmp2425;
	wire signed [31:0] w_sys_tmp2430;
	wire signed [31:0] w_sys_tmp2431;
	wire signed [31:0] w_sys_tmp2436;
	wire signed [31:0] w_sys_tmp2437;
	wire signed [31:0] w_sys_tmp2442;
	wire signed [31:0] w_sys_tmp2443;
	wire signed [31:0] w_sys_tmp2448;
	wire signed [31:0] w_sys_tmp2449;
	wire signed [31:0] w_sys_tmp2454;
	wire signed [31:0] w_sys_tmp2455;
	wire signed [31:0] w_sys_tmp2460;
	wire signed [31:0] w_sys_tmp2461;
	wire signed [31:0] w_sys_tmp2466;
	wire signed [31:0] w_sys_tmp2467;
	wire signed [31:0] w_sys_tmp2472;
	wire signed [31:0] w_sys_tmp2473;
	wire signed [31:0] w_sys_tmp2478;
	wire signed [31:0] w_sys_tmp2479;
	wire signed [31:0] w_sys_tmp2484;
	wire signed [31:0] w_sys_tmp2485;
	wire signed [31:0] w_sys_tmp2490;
	wire signed [31:0] w_sys_tmp2491;
	wire signed [31:0] w_sys_tmp2496;
	wire signed [31:0] w_sys_tmp2497;
	wire signed [31:0] w_sys_tmp2502;
	wire signed [31:0] w_sys_tmp2503;
	wire signed [31:0] w_sys_tmp2508;
	wire signed [31:0] w_sys_tmp2509;
	wire signed [31:0] w_sys_tmp2514;
	wire signed [31:0] w_sys_tmp2515;
	wire signed [31:0] w_sys_tmp2520;
	wire signed [31:0] w_sys_tmp2521;
	wire signed [31:0] w_sys_tmp2526;
	wire signed [31:0] w_sys_tmp2527;
	wire signed [31:0] w_sys_tmp2543;
	wire signed [31:0] w_sys_tmp2544;
	wire               w_sys_tmp2545;
	wire               w_sys_tmp2546;
	wire signed [31:0] w_sys_tmp2547;
	wire signed [31:0] w_sys_tmp2550;
	wire signed [31:0] w_sys_tmp2551;
	wire        [31:0] w_sys_tmp2552;
	wire signed [31:0] w_sys_tmp2553;
	wire signed [31:0] w_sys_tmp2554;
	wire signed [31:0] w_sys_tmp2555;
	wire signed [31:0] w_sys_tmp2557;
	wire signed [31:0] w_sys_tmp2558;
	wire signed [31:0] w_sys_tmp2564;
	wire signed [31:0] w_sys_tmp2565;
	wire signed [31:0] w_sys_tmp2571;
	wire signed [31:0] w_sys_tmp2572;
	wire signed [31:0] w_sys_tmp2578;
	wire signed [31:0] w_sys_tmp2579;
	wire signed [31:0] w_sys_tmp2585;
	wire signed [31:0] w_sys_tmp2586;
	wire signed [31:0] w_sys_tmp2592;
	wire signed [31:0] w_sys_tmp2593;
	wire signed [31:0] w_sys_tmp2599;
	wire signed [31:0] w_sys_tmp2600;
	wire signed [31:0] w_sys_tmp2606;
	wire signed [31:0] w_sys_tmp2607;
	wire signed [31:0] w_sys_tmp2613;
	wire signed [31:0] w_sys_tmp2614;
	wire signed [31:0] w_sys_tmp2618;
	wire signed [31:0] w_sys_tmp2619;
	wire signed [31:0] w_sys_tmp2623;
	wire signed [31:0] w_sys_tmp2624;
	wire signed [31:0] w_sys_tmp2628;
	wire signed [31:0] w_sys_tmp2629;
	wire signed [31:0] w_sys_tmp2633;
	wire signed [31:0] w_sys_tmp2634;
	wire signed [31:0] w_sys_tmp2638;
	wire signed [31:0] w_sys_tmp2639;
	wire signed [31:0] w_sys_tmp2643;
	wire signed [31:0] w_sys_tmp2644;
	wire signed [31:0] w_sys_tmp2648;
	wire signed [31:0] w_sys_tmp2649;
	wire signed [31:0] w_sys_tmp2653;
	wire signed [31:0] w_sys_tmp2654;
	wire signed [31:0] w_sys_tmp2658;
	wire signed [31:0] w_sys_tmp2659;
	wire signed [31:0] w_sys_tmp2662;
	wire signed [31:0] w_sys_tmp2663;
	wire               w_sys_tmp2664;
	wire               w_sys_tmp2665;
	wire signed [31:0] w_sys_tmp2666;
	wire signed [31:0] w_sys_tmp2669;
	wire signed [31:0] w_sys_tmp2670;
	wire        [31:0] w_sys_tmp2671;
	wire signed [31:0] w_sys_tmp2672;
	wire signed [31:0] w_sys_tmp2673;
	wire signed [31:0] w_sys_tmp2674;
	wire signed [31:0] w_sys_tmp2676;
	wire signed [31:0] w_sys_tmp2677;
	wire signed [31:0] w_sys_tmp2683;
	wire signed [31:0] w_sys_tmp2684;
	wire signed [31:0] w_sys_tmp2690;
	wire signed [31:0] w_sys_tmp2691;
	wire signed [31:0] w_sys_tmp2697;
	wire signed [31:0] w_sys_tmp2698;
	wire signed [31:0] w_sys_tmp2704;
	wire signed [31:0] w_sys_tmp2705;
	wire signed [31:0] w_sys_tmp2711;
	wire signed [31:0] w_sys_tmp2712;
	wire signed [31:0] w_sys_tmp2718;
	wire signed [31:0] w_sys_tmp2719;
	wire signed [31:0] w_sys_tmp2725;
	wire signed [31:0] w_sys_tmp2726;
	wire signed [31:0] w_sys_tmp2732;
	wire signed [31:0] w_sys_tmp2733;
	wire signed [31:0] w_sys_tmp2737;
	wire signed [31:0] w_sys_tmp2738;
	wire signed [31:0] w_sys_tmp2742;
	wire signed [31:0] w_sys_tmp2743;
	wire signed [31:0] w_sys_tmp2747;
	wire signed [31:0] w_sys_tmp2748;
	wire signed [31:0] w_sys_tmp2752;
	wire signed [31:0] w_sys_tmp2753;
	wire signed [31:0] w_sys_tmp2757;
	wire signed [31:0] w_sys_tmp2758;
	wire signed [31:0] w_sys_tmp2762;
	wire signed [31:0] w_sys_tmp2763;
	wire signed [31:0] w_sys_tmp2767;
	wire signed [31:0] w_sys_tmp2768;
	wire signed [31:0] w_sys_tmp2772;
	wire signed [31:0] w_sys_tmp2773;
	wire signed [31:0] w_sys_tmp2777;
	wire signed [31:0] w_sys_tmp2778;
	wire signed [31:0] w_sys_tmp2781;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 3'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 9'h1);
	assign w_fld_u_0_addr_0 = 9'sh0;
	assign w_fld_u_0_datain_0 = 32'h0;
	assign w_fld_u_0_r_w_0 = 1'h0;
	assign w_fld_u_0_ce_0 = w_sys_ce;
	assign w_fld_u_0_ce_1 = w_sys_ce;
	assign w_fld_uu_1_addr_0 = 9'sh0;
	assign w_fld_uu_1_datain_0 = 32'h0;
	assign w_fld_uu_1_r_w_0 = 1'h0;
	assign w_fld_uu_1_ce_0 = w_sys_ce;
	assign w_fld_uu_1_ce_1 = w_sys_ce;
	assign w_sub03_u_addr = ( (|r_sys_processing_methodID) ? r_sub03_u_addr : 9'sh0 ) ;
	assign w_sub03_u_datain = ( (|r_sys_processing_methodID) ? r_sub03_u_datain : 32'h0 ) ;
	assign w_sub03_u_r_w = ( (|r_sys_processing_methodID) ? r_sub03_u_r_w : 1'h0 ) ;
	assign w_sub03_result_addr = ( (|r_sys_processing_methodID) ? r_sub03_result_addr : 9'sh0 ) ;
	assign w_sub03_result_datain = ( (|r_sys_processing_methodID) ? r_sub03_result_datain : 32'h0 ) ;
	assign w_sub03_result_r_w = ( (|r_sys_processing_methodID) ? r_sub03_result_r_w : 1'h0 ) ;
	assign w_sub02_u_addr = ( (|r_sys_processing_methodID) ? r_sub02_u_addr : 9'sh0 ) ;
	assign w_sub02_u_datain = ( (|r_sys_processing_methodID) ? r_sub02_u_datain : 32'h0 ) ;
	assign w_sub02_u_r_w = ( (|r_sys_processing_methodID) ? r_sub02_u_r_w : 1'h0 ) ;
	assign w_sub02_result_addr = ( (|r_sys_processing_methodID) ? r_sub02_result_addr : 9'sh0 ) ;
	assign w_sub02_result_datain = ( (|r_sys_processing_methodID) ? r_sub02_result_datain : 32'h0 ) ;
	assign w_sub02_result_r_w = ( (|r_sys_processing_methodID) ? r_sub02_result_r_w : 1'h0 ) ;
	assign w_sub01_u_addr = ( (|r_sys_processing_methodID) ? r_sub01_u_addr : 9'sh0 ) ;
	assign w_sub01_u_datain = ( (|r_sys_processing_methodID) ? r_sub01_u_datain : 32'h0 ) ;
	assign w_sub01_u_r_w = ( (|r_sys_processing_methodID) ? r_sub01_u_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 9'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub00_u_addr = ( (|r_sys_processing_methodID) ? r_sub00_u_addr : 9'sh0 ) ;
	assign w_sub00_u_datain = ( (|r_sys_processing_methodID) ? r_sub00_u_datain : 32'h0 ) ;
	assign w_sub00_u_r_w = ( (|r_sys_processing_methodID) ? r_sub00_u_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 9'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh00000015;
	assign w_sys_tmp3 = 32'h3d4ccccd;
	assign w_sys_tmp5 = 32'sh00000002;
	assign w_sys_tmp6 = ( !w_sys_tmp7 );
	assign w_sys_tmp7 = (r_run_my_10 < r_run_k_6);
	assign w_sys_tmp8 = (r_run_k_6 + w_sys_intOne);
	assign w_sys_tmp9 = ( !w_sys_tmp10 );
	assign w_sys_tmp10 = (r_run_mx_9 < r_run_j_7);
	assign w_sys_tmp13 = (w_sys_tmp14 + r_run_k_6);
	assign w_sys_tmp14 = (r_run_j_7 * w_sys_tmp15);
	assign w_sys_tmp15 = 32'sh00000015;
	assign w_sys_tmp16 = 32'h0;
	assign w_sys_tmp18 = (w_sys_tmp19 + r_run_k_6);
	assign w_sys_tmp19 = (r_run_copy0_j_14 * w_sys_tmp15);
	assign w_sys_tmp22 = (r_run_copy0_j_14 + w_sys_intOne);
	assign w_sys_tmp23 = (r_run_j_7 + w_sys_intOne);
	assign w_sys_tmp780 = ( !w_sys_tmp781 );
	assign w_sys_tmp781 = (r_run_nlast_11 < r_run_n_8);
	assign w_sys_tmp782 = (r_run_n_8 + w_sys_intOne);
	assign w_sys_tmp783 = ( !w_sys_tmp784 );
	assign w_sys_tmp784 = (r_run_my_10 < r_run_j_7);
	assign w_sys_tmp787 = (w_sys_tmp788 + r_run_j_7);
	assign w_sys_tmp788 = 32'sh00000015;
	assign w_sys_tmp789 = 32'h3f000000;
	assign w_sys_tmp791 = (w_sys_tmp792 + r_run_copy2_j_17);
	assign w_sys_tmp792 = (r_run_mx_9 * w_sys_tmp788);
	assign w_sys_tmp794 = 32'h0;
	assign w_sys_tmp796 = (w_sys_tmp797 + w_sys_intOne);
	assign w_sys_tmp797 = (r_run_copy1_j_16 * w_sys_tmp788);
	assign w_sys_tmp799 = 32'h3f800000;
	assign w_sys_tmp801 = (w_sys_tmp802 + r_run_my_10);
	assign w_sys_tmp802 = (r_run_copy0_j_15 * w_sys_tmp788);
	assign w_sys_tmp805 = (r_run_copy0_j_15 + w_sys_intOne);
	assign w_sys_tmp806 = (r_run_copy1_j_16 + w_sys_intOne);
	assign w_sys_tmp807 = (r_run_copy2_j_17 + w_sys_intOne);
	assign w_sys_tmp808 = (r_run_j_7 + w_sys_intOne);
	assign w_sys_tmp2258 = 32'sh0000000a;
	assign w_sys_tmp2259 = ( !w_sys_tmp2260 );
	assign w_sys_tmp2260 = (r_run_my_10 < r_run_k_6);
	assign w_sys_tmp2263 = (w_sys_tmp2264 + r_run_k_6);
	assign w_sys_tmp2264 = 32'sh000000d2;
	assign w_sys_tmp2265 = w_fld_u_0_dataout_1;
	assign w_sys_tmp2269 = (w_sys_tmp2270 + r_run_k_6);
	assign w_sys_tmp2270 = 32'sh000000e7;
	assign w_sys_tmp2275 = (w_sys_tmp2276 + r_run_k_6);
	assign w_sys_tmp2276 = 32'sh000000fc;
	assign w_sys_tmp2281 = (w_sys_tmp2282 + r_run_k_6);
	assign w_sys_tmp2282 = 32'sh00000111;
	assign w_sys_tmp2287 = (w_sys_tmp2288 + r_run_k_6);
	assign w_sys_tmp2288 = 32'sh00000126;
	assign w_sys_tmp2293 = (w_sys_tmp2294 + r_run_k_6);
	assign w_sys_tmp2294 = 32'sh0000013b;
	assign w_sys_tmp2299 = (w_sys_tmp2300 + r_run_k_6);
	assign w_sys_tmp2300 = 32'sh00000150;
	assign w_sys_tmp2305 = (w_sys_tmp2306 + r_run_k_6);
	assign w_sys_tmp2306 = 32'sh00000165;
	assign w_sys_tmp2311 = (w_sys_tmp2312 + r_run_k_6);
	assign w_sys_tmp2312 = 32'sh0000017a;
	assign w_sys_tmp2317 = (w_sys_tmp2318 + r_run_k_6);
	assign w_sys_tmp2318 = 32'sh0000018f;
	assign w_sys_tmp2323 = (w_sys_tmp2324 + r_run_k_6);
	assign w_sys_tmp2324 = 32'sh000001a4;
	assign w_sys_tmp2329 = (w_sys_tmp2330 + r_run_k_6);
	assign w_sys_tmp2330 = 32'sh000001b9;
	assign w_sys_tmp2335 = (w_sys_tmp2336 + r_run_k_6);
	assign w_sys_tmp2336 = 32'sh00000015;
	assign w_sys_tmp2341 = (w_sys_tmp2342 + r_run_k_6);
	assign w_sys_tmp2342 = 32'sh0000002a;
	assign w_sys_tmp2347 = (w_sys_tmp2348 + r_run_k_6);
	assign w_sys_tmp2348 = 32'sh0000003f;
	assign w_sys_tmp2353 = (w_sys_tmp2354 + r_run_k_6);
	assign w_sys_tmp2354 = 32'sh00000054;
	assign w_sys_tmp2359 = (w_sys_tmp2360 + r_run_k_6);
	assign w_sys_tmp2360 = 32'sh00000069;
	assign w_sys_tmp2365 = (w_sys_tmp2366 + r_run_k_6);
	assign w_sys_tmp2366 = 32'sh0000007e;
	assign w_sys_tmp2371 = (w_sys_tmp2372 + r_run_k_6);
	assign w_sys_tmp2372 = 32'sh00000093;
	assign w_sys_tmp2377 = (w_sys_tmp2378 + r_run_k_6);
	assign w_sys_tmp2378 = 32'sh000000a8;
	assign w_sys_tmp2383 = (w_sys_tmp2384 + r_run_k_6);
	assign w_sys_tmp2384 = 32'sh000000bd;
	assign w_sys_tmp2400 = (r_run_k_6 + w_sys_intOne);
	assign w_sys_tmp2401 = ( !w_sys_tmp2402 );
	assign w_sys_tmp2402 = (w_sys_tmp2403 < r_run_k_6);
	assign w_sys_tmp2403 = 32'sh0000000b;
	assign w_sys_tmp2406 = (w_sys_tmp2407 + r_run_k_6);
	assign w_sys_tmp2407 = 32'sh000000d2;
	assign w_sys_tmp2408 = w_fld_u_0_dataout_1;
	assign w_sys_tmp2412 = (w_sys_tmp2413 + r_run_k_6);
	assign w_sys_tmp2413 = 32'sh000000e7;
	assign w_sys_tmp2418 = (w_sys_tmp2419 + r_run_k_6);
	assign w_sys_tmp2419 = 32'sh000000fc;
	assign w_sys_tmp2424 = (w_sys_tmp2425 + r_run_k_6);
	assign w_sys_tmp2425 = 32'sh00000111;
	assign w_sys_tmp2430 = (w_sys_tmp2431 + r_run_k_6);
	assign w_sys_tmp2431 = 32'sh00000126;
	assign w_sys_tmp2436 = (w_sys_tmp2437 + r_run_k_6);
	assign w_sys_tmp2437 = 32'sh0000013b;
	assign w_sys_tmp2442 = (w_sys_tmp2443 + r_run_k_6);
	assign w_sys_tmp2443 = 32'sh00000150;
	assign w_sys_tmp2448 = (w_sys_tmp2449 + r_run_k_6);
	assign w_sys_tmp2449 = 32'sh00000165;
	assign w_sys_tmp2454 = (w_sys_tmp2455 + r_run_k_6);
	assign w_sys_tmp2455 = 32'sh0000017a;
	assign w_sys_tmp2460 = (w_sys_tmp2461 + r_run_k_6);
	assign w_sys_tmp2461 = 32'sh0000018f;
	assign w_sys_tmp2466 = (w_sys_tmp2467 + r_run_k_6);
	assign w_sys_tmp2467 = 32'sh000001a4;
	assign w_sys_tmp2472 = (w_sys_tmp2473 + r_run_k_6);
	assign w_sys_tmp2473 = 32'sh000001b9;
	assign w_sys_tmp2478 = (w_sys_tmp2479 + r_run_k_6);
	assign w_sys_tmp2479 = 32'sh00000015;
	assign w_sys_tmp2484 = (w_sys_tmp2485 + r_run_k_6);
	assign w_sys_tmp2485 = 32'sh0000002a;
	assign w_sys_tmp2490 = (w_sys_tmp2491 + r_run_k_6);
	assign w_sys_tmp2491 = 32'sh0000003f;
	assign w_sys_tmp2496 = (w_sys_tmp2497 + r_run_k_6);
	assign w_sys_tmp2497 = 32'sh00000054;
	assign w_sys_tmp2502 = (w_sys_tmp2503 + r_run_k_6);
	assign w_sys_tmp2503 = 32'sh00000069;
	assign w_sys_tmp2508 = (w_sys_tmp2509 + r_run_k_6);
	assign w_sys_tmp2509 = 32'sh0000007e;
	assign w_sys_tmp2514 = (w_sys_tmp2515 + r_run_k_6);
	assign w_sys_tmp2515 = 32'sh00000093;
	assign w_sys_tmp2520 = (w_sys_tmp2521 + r_run_k_6);
	assign w_sys_tmp2521 = 32'sh000000a8;
	assign w_sys_tmp2526 = (w_sys_tmp2527 + r_run_k_6);
	assign w_sys_tmp2527 = 32'sh000000bd;
	assign w_sys_tmp2543 = (r_run_k_6 + w_sys_intOne);
	assign w_sys_tmp2544 = 32'sh00000002;
	assign w_sys_tmp2545 = ( !w_sys_tmp2546 );
	assign w_sys_tmp2546 = (w_sys_tmp2547 < r_run_k_6);
	assign w_sys_tmp2547 = 32'sh0000000a;
	assign w_sys_tmp2550 = (w_sys_tmp2551 + r_run_k_6);
	assign w_sys_tmp2551 = 32'sh0000002a;
	assign w_sys_tmp2552 = w_sub00_result_dataout;
	assign w_sys_tmp2553 = (w_sys_tmp2554 + r_run_k_6);
	assign w_sys_tmp2554 = (r_run_j_7 * w_sys_tmp2555);
	assign w_sys_tmp2555 = 32'sh00000015;
	assign w_sys_tmp2557 = (w_sys_tmp2558 + r_run_k_6);
	assign w_sys_tmp2558 = 32'sh0000003f;
	assign w_sys_tmp2564 = (w_sys_tmp2565 + r_run_k_6);
	assign w_sys_tmp2565 = 32'sh00000054;
	assign w_sys_tmp2571 = (w_sys_tmp2572 + r_run_k_6);
	assign w_sys_tmp2572 = 32'sh00000069;
	assign w_sys_tmp2578 = (w_sys_tmp2579 + r_run_k_6);
	assign w_sys_tmp2579 = 32'sh0000007e;
	assign w_sys_tmp2585 = (w_sys_tmp2586 + r_run_k_6);
	assign w_sys_tmp2586 = 32'sh00000093;
	assign w_sys_tmp2592 = (w_sys_tmp2593 + r_run_k_6);
	assign w_sys_tmp2593 = 32'sh000000a8;
	assign w_sys_tmp2599 = (w_sys_tmp2600 + r_run_k_6);
	assign w_sys_tmp2600 = 32'sh000000bd;
	assign w_sys_tmp2606 = (w_sys_tmp2607 + r_run_k_6);
	assign w_sys_tmp2607 = 32'sh000000d2;
	assign w_sys_tmp2613 = (w_sys_tmp2614 + r_run_k_6);
	assign w_sys_tmp2614 = 32'sh000000e7;
	assign w_sys_tmp2618 = (w_sys_tmp2619 + r_run_k_6);
	assign w_sys_tmp2619 = 32'sh000000fc;
	assign w_sys_tmp2623 = (w_sys_tmp2624 + r_run_k_6);
	assign w_sys_tmp2624 = 32'sh00000111;
	assign w_sys_tmp2628 = (w_sys_tmp2629 + r_run_k_6);
	assign w_sys_tmp2629 = 32'sh00000126;
	assign w_sys_tmp2633 = (w_sys_tmp2634 + r_run_k_6);
	assign w_sys_tmp2634 = 32'sh0000013b;
	assign w_sys_tmp2638 = (w_sys_tmp2639 + r_run_k_6);
	assign w_sys_tmp2639 = 32'sh00000150;
	assign w_sys_tmp2643 = (w_sys_tmp2644 + r_run_k_6);
	assign w_sys_tmp2644 = 32'sh00000165;
	assign w_sys_tmp2648 = (w_sys_tmp2649 + r_run_k_6);
	assign w_sys_tmp2649 = 32'sh0000017a;
	assign w_sys_tmp2653 = (w_sys_tmp2654 + r_run_k_6);
	assign w_sys_tmp2654 = 32'sh0000018f;
	assign w_sys_tmp2658 = (w_sys_tmp2659 + r_run_k_6);
	assign w_sys_tmp2659 = 32'sh000001a4;
	assign w_sys_tmp2662 = (r_run_k_6 + w_sys_intOne);
	assign w_sys_tmp2663 = 32'sh0000000b;
	assign w_sys_tmp2664 = ( !w_sys_tmp2665 );
	assign w_sys_tmp2665 = (w_sys_tmp2666 < r_run_k_6);
	assign w_sys_tmp2666 = 32'sh00000014;
	assign w_sys_tmp2669 = (w_sys_tmp2670 + r_run_k_6);
	assign w_sys_tmp2670 = 32'sh0000002a;
	assign w_sys_tmp2671 = w_sub02_result_dataout;
	assign w_sys_tmp2672 = (w_sys_tmp2673 + r_run_k_6);
	assign w_sys_tmp2673 = (r_run_j_7 * w_sys_tmp2674);
	assign w_sys_tmp2674 = 32'sh00000015;
	assign w_sys_tmp2676 = (w_sys_tmp2677 + r_run_k_6);
	assign w_sys_tmp2677 = 32'sh0000003f;
	assign w_sys_tmp2683 = (w_sys_tmp2684 + r_run_k_6);
	assign w_sys_tmp2684 = 32'sh00000054;
	assign w_sys_tmp2690 = (w_sys_tmp2691 + r_run_k_6);
	assign w_sys_tmp2691 = 32'sh00000069;
	assign w_sys_tmp2697 = (w_sys_tmp2698 + r_run_k_6);
	assign w_sys_tmp2698 = 32'sh0000007e;
	assign w_sys_tmp2704 = (w_sys_tmp2705 + r_run_k_6);
	assign w_sys_tmp2705 = 32'sh00000093;
	assign w_sys_tmp2711 = (w_sys_tmp2712 + r_run_k_6);
	assign w_sys_tmp2712 = 32'sh000000a8;
	assign w_sys_tmp2718 = (w_sys_tmp2719 + r_run_k_6);
	assign w_sys_tmp2719 = 32'sh000000bd;
	assign w_sys_tmp2725 = (w_sys_tmp2726 + r_run_k_6);
	assign w_sys_tmp2726 = 32'sh000000d2;
	assign w_sys_tmp2732 = (w_sys_tmp2733 + r_run_k_6);
	assign w_sys_tmp2733 = 32'sh000000e7;
	assign w_sys_tmp2737 = (w_sys_tmp2738 + r_run_k_6);
	assign w_sys_tmp2738 = 32'sh000000fc;
	assign w_sys_tmp2742 = (w_sys_tmp2743 + r_run_k_6);
	assign w_sys_tmp2743 = 32'sh00000111;
	assign w_sys_tmp2747 = (w_sys_tmp2748 + r_run_k_6);
	assign w_sys_tmp2748 = 32'sh00000126;
	assign w_sys_tmp2752 = (w_sys_tmp2753 + r_run_k_6);
	assign w_sys_tmp2753 = 32'sh0000013b;
	assign w_sys_tmp2757 = (w_sys_tmp2758 + r_run_k_6);
	assign w_sys_tmp2758 = 32'sh00000150;
	assign w_sys_tmp2762 = (w_sys_tmp2763 + r_run_k_6);
	assign w_sys_tmp2763 = 32'sh00000165;
	assign w_sys_tmp2767 = (w_sys_tmp2768 + r_run_k_6);
	assign w_sys_tmp2768 = 32'sh0000017a;
	assign w_sys_tmp2772 = (w_sys_tmp2773 + r_run_k_6);
	assign w_sys_tmp2773 = 32'sh0000018f;
	assign w_sys_tmp2777 = (w_sys_tmp2778 + r_run_k_6);
	assign w_sys_tmp2778 = 32'sh000001a4;
	assign w_sys_tmp2781 = (r_run_k_6 + w_sys_intOne);


	sub03
		sub03_inst(
			.i_fld_result_1_addr_0 (w_sub03_result_addr),
			.i_fld_result_1_datain_0 (w_sub03_result_datain),
			.o_fld_result_1_dataout_0 (w_sub03_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub03_result_r_w),
			.i_fld_u_0_addr_0 (w_sub03_u_addr),
			.i_fld_u_0_datain_0 (w_sub03_u_datain),
			.o_fld_u_0_dataout_0 (w_sub03_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub03_u_r_w),
			.o_run_busy (w_sub03_run_busy),
			.i_run_req (r_sub03_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub02
		sub02_inst(
			.i_fld_result_1_addr_0 (w_sub02_result_addr),
			.i_fld_result_1_datain_0 (w_sub02_result_datain),
			.o_fld_result_1_dataout_0 (w_sub02_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub02_result_r_w),
			.i_fld_u_0_addr_0 (w_sub02_u_addr),
			.i_fld_u_0_datain_0 (w_sub02_u_datain),
			.o_fld_u_0_dataout_0 (w_sub02_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub02_u_r_w),
			.o_run_busy (w_sub02_run_busy),
			.i_run_req (r_sub02_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub01
		sub01_inst(
			.i_fld_result_1_addr_0 (w_sub01_result_addr),
			.i_fld_result_1_datain_0 (w_sub01_result_datain),
			.o_fld_result_1_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub01_result_r_w),
			.i_fld_u_0_addr_0 (w_sub01_u_addr),
			.i_fld_u_0_datain_0 (w_sub01_u_datain),
			.o_fld_u_0_dataout_0 (w_sub01_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub01_u_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub00
		sub00_inst(
			.i_fld_result_1_addr_0 (w_sub00_result_addr),
			.i_fld_result_1_datain_0 (w_sub00_result_datain),
			.o_fld_result_1_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub00_result_r_w),
			.i_fld_u_0_addr_0 (w_sub00_u_addr),
			.i_fld_u_0_datain_0 (w_sub00_u_datain),
			.o_fld_u_0_dataout_0 (w_sub00_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub00_u_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(9), .WORDS(484) )
		dpram_u_0(
			.clk (clock),
			.ce_0 (w_fld_u_0_ce_0),
			.addr_0 (w_fld_u_0_addr_0),
			.datain_0 (w_fld_u_0_datain_0),
			.dataout_0 (w_fld_u_0_dataout_0),
			.r_w_0 (w_fld_u_0_r_w_0),
			.ce_1 (w_fld_u_0_ce_1),
			.addr_1 (r_fld_u_0_addr_1),
			.datain_1 (r_fld_u_0_datain_1),
			.dataout_1 (w_fld_u_0_dataout_1),
			.r_w_1 (r_fld_u_0_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(9), .WORDS(484) )
		dpram_uu_1(
			.clk (clock),
			.ce_0 (w_fld_uu_1_ce_0),
			.addr_0 (w_fld_uu_1_addr_0),
			.datain_0 (w_fld_uu_1_datain_0),
			.dataout_0 (w_fld_uu_1_dataout_0),
			.r_w_0 (w_fld_uu_1_r_w_0),
			.ce_1 (w_fld_uu_1_ce_1),
			.addr_1 (r_fld_uu_1_addr_1),
			.datain_1 (r_fld_uu_1_datain_1),
			.dataout_1 (w_fld_uu_1_dataout_1),
			.r_w_1 (r_fld_uu_1_r_w_1)
		);

	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h36: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 6'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_phase <= 6'h2;
						end

						6'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'h4;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6) ? 6'h9 : 6'hf);

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'ha;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp9) ? 6'hd : 6'h6);

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h3f)) begin
										r_sys_run_phase <= 6'ha;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'h10;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp780) ? 6'h14 : 6'h36);

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'h10;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'h15;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp783) ? 6'h18 : 6'h1a);

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'hff)) begin
										r_sys_run_phase <= 6'h15;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'h1b;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2259) ? 6'h1e : 6'h1f);

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_run_phase <= 6'h1b;

									end
								end

							endcase
						end

						6'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_phase <= 6'h21;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'h22;

									end
								end

							endcase
						end

						6'h22: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2401) ? 6'h25 : 6'h26);

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_run_phase <= 6'h22;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_phase <= 6'h28;

									end
								end

							endcase
						end

						6'h28: begin

							case(r_sys_run_stage) 
								3'h3: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_phase <= 6'h2a;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'h2b;

									end
								end

							endcase
						end

						6'h2b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2545) ? 6'h2e : 6'h30);

									end
								end

							endcase
						end

						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_run_phase <= 6'h2b;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'h31;

									end
								end

							endcase
						end

						6'h31: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2664) ? 6'h34 : 6'h11);

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_run_phase <= 6'h31;

									end
								end

							endcase
						end

						6'h36: begin
							r_sys_run_phase <= 6'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 3'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h3f)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'hff)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h22: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h28: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h2: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h3: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h2b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h31: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 9'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h3f)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h3e)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'hfe)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==9'hff)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h17)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h22: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h17)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h28: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub00_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								3'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub01_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								3'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub02_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								3'h3: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub03_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h2b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h31: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						6'h36: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_addr_1 <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h3f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp13[8:0] );

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h2) || (r_sys_run_step==9'h6) || (r_sys_run_step==9'ha) || (r_sys_run_step==9'he) || (r_sys_run_step==9'h12) || (r_sys_run_step==9'h16) || (r_sys_run_step==9'h1a) || (r_sys_run_step==9'h1e) || (r_sys_run_step==9'h22) || (r_sys_run_step==9'h26) || (r_sys_run_step==9'h2a) || (r_sys_run_step==9'h2e) || (r_sys_run_step==9'h32) || (r_sys_run_step==9'h36) || (r_sys_run_step==9'h3a) || (r_sys_run_step==9'h3e) || (r_sys_run_step==9'h42) || (r_sys_run_step==9'h46) || (r_sys_run_step==9'h4a) || (r_sys_run_step==9'h4e) || (r_sys_run_step==9'h52) || (r_sys_run_step==9'h56) || (r_sys_run_step==9'h5a) || (r_sys_run_step==9'h5e) || (r_sys_run_step==9'h62) || (r_sys_run_step==9'h66) || (r_sys_run_step==9'h6a) || (r_sys_run_step==9'h6e) || (r_sys_run_step==9'h72) || (r_sys_run_step==9'h76) || (r_sys_run_step==9'h7a) || (r_sys_run_step==9'h7e) || (r_sys_run_step==9'h82) || (r_sys_run_step==9'h86) || (r_sys_run_step==9'h8a) || (r_sys_run_step==9'h8e) || (r_sys_run_step==9'h92) || (r_sys_run_step==9'h96) || (r_sys_run_step==9'h9a) || (r_sys_run_step==9'h9e) || (r_sys_run_step==9'ha2) || (r_sys_run_step==9'ha6) || (r_sys_run_step==9'haa) || (r_sys_run_step==9'hae) || (r_sys_run_step==9'hb2) || (r_sys_run_step==9'hb6) || (r_sys_run_step==9'hba) || (r_sys_run_step==9'hbe) || (r_sys_run_step==9'hc2) || (r_sys_run_step==9'hc6) || (r_sys_run_step==9'hca) || (r_sys_run_step==9'hce) || (r_sys_run_step==9'hd2) || (r_sys_run_step==9'hd6) || (r_sys_run_step==9'hda) || (r_sys_run_step==9'hde) || (r_sys_run_step==9'he2) || (r_sys_run_step==9'he6) || (r_sys_run_step==9'hea) || (r_sys_run_step==9'hee) || (r_sys_run_step==9'hf2) || (r_sys_run_step==9'hf6) || (r_sys_run_step==9'hfa) || (r_sys_run_step==9'hfe)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp796[8:0] );

									end
									else
									if((r_sys_run_step==9'h0) || (r_sys_run_step==9'h4) || (r_sys_run_step==9'h8) || (r_sys_run_step==9'hc) || (r_sys_run_step==9'h10) || (r_sys_run_step==9'h14) || (r_sys_run_step==9'h18) || (r_sys_run_step==9'h1c) || (r_sys_run_step==9'h20) || (r_sys_run_step==9'h24) || (r_sys_run_step==9'h28) || (r_sys_run_step==9'h2c) || (r_sys_run_step==9'h30) || (r_sys_run_step==9'h34) || (r_sys_run_step==9'h38) || (r_sys_run_step==9'h3c) || (r_sys_run_step==9'h40) || (r_sys_run_step==9'h44) || (r_sys_run_step==9'h48) || (r_sys_run_step==9'h4c) || (r_sys_run_step==9'h50) || (r_sys_run_step==9'h54) || (r_sys_run_step==9'h58) || (r_sys_run_step==9'h5c) || (r_sys_run_step==9'h60) || (r_sys_run_step==9'h64) || (r_sys_run_step==9'h68) || (r_sys_run_step==9'h6c) || (r_sys_run_step==9'h70) || (r_sys_run_step==9'h74) || (r_sys_run_step==9'h78) || (r_sys_run_step==9'h7c) || (r_sys_run_step==9'h80) || (r_sys_run_step==9'h84) || (r_sys_run_step==9'h88) || (r_sys_run_step==9'h8c) || (r_sys_run_step==9'h90) || (r_sys_run_step==9'h94) || (r_sys_run_step==9'h98) || (r_sys_run_step==9'h9c) || (r_sys_run_step==9'ha0) || (r_sys_run_step==9'ha4) || (r_sys_run_step==9'ha8) || (r_sys_run_step==9'hac) || (r_sys_run_step==9'hb0) || (r_sys_run_step==9'hb4) || (r_sys_run_step==9'hb8) || (r_sys_run_step==9'hbc) || (r_sys_run_step==9'hc0) || (r_sys_run_step==9'hc4) || (r_sys_run_step==9'hc8) || (r_sys_run_step==9'hcc) || (r_sys_run_step==9'hd0) || (r_sys_run_step==9'hd4) || (r_sys_run_step==9'hd8) || (r_sys_run_step==9'hdc) || (r_sys_run_step==9'he0) || (r_sys_run_step==9'he4) || (r_sys_run_step==9'he8) || (r_sys_run_step==9'hec) || (r_sys_run_step==9'hf0) || (r_sys_run_step==9'hf4) || (r_sys_run_step==9'hf8) || (r_sys_run_step==9'hfc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp787[8:0] );

									end
									else
									if((r_sys_run_step==9'h3) || (r_sys_run_step==9'h7) || (r_sys_run_step==9'hb) || (r_sys_run_step==9'hf) || (r_sys_run_step==9'h13) || (r_sys_run_step==9'h17) || (r_sys_run_step==9'h1b) || (r_sys_run_step==9'h1f) || (r_sys_run_step==9'h23) || (r_sys_run_step==9'h27) || (r_sys_run_step==9'h2b) || (r_sys_run_step==9'h2f) || (r_sys_run_step==9'h33) || (r_sys_run_step==9'h37) || (r_sys_run_step==9'h3b) || (r_sys_run_step==9'h3f) || (r_sys_run_step==9'h43) || (r_sys_run_step==9'h47) || (r_sys_run_step==9'h4b) || (r_sys_run_step==9'h4f) || (r_sys_run_step==9'h53) || (r_sys_run_step==9'h57) || (r_sys_run_step==9'h5b) || (r_sys_run_step==9'h5f) || (r_sys_run_step==9'h63) || (r_sys_run_step==9'h67) || (r_sys_run_step==9'h6b) || (r_sys_run_step==9'h6f) || (r_sys_run_step==9'h73) || (r_sys_run_step==9'h77) || (r_sys_run_step==9'h7b) || (r_sys_run_step==9'h7f) || (r_sys_run_step==9'h83) || (r_sys_run_step==9'h87) || (r_sys_run_step==9'h8b) || (r_sys_run_step==9'h8f) || (r_sys_run_step==9'h93) || (r_sys_run_step==9'h97) || (r_sys_run_step==9'h9b) || (r_sys_run_step==9'h9f) || (r_sys_run_step==9'ha3) || (r_sys_run_step==9'ha7) || (r_sys_run_step==9'hab) || (r_sys_run_step==9'haf) || (r_sys_run_step==9'hb3) || (r_sys_run_step==9'hb7) || (r_sys_run_step==9'hbb) || (r_sys_run_step==9'hbf) || (r_sys_run_step==9'hc3) || (r_sys_run_step==9'hc7) || (r_sys_run_step==9'hcb) || (r_sys_run_step==9'hcf) || (r_sys_run_step==9'hd3) || (r_sys_run_step==9'hd7) || (r_sys_run_step==9'hdb) || (r_sys_run_step==9'hdf) || (r_sys_run_step==9'he3) || (r_sys_run_step==9'he7) || (r_sys_run_step==9'heb) || (r_sys_run_step==9'hef) || (r_sys_run_step==9'hf3) || (r_sys_run_step==9'hf7) || (r_sys_run_step==9'hfb) || (r_sys_run_step==9'hff)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp801[8:0] );

									end
									else
									if((r_sys_run_step==9'h1) || (r_sys_run_step==9'h5) || (r_sys_run_step==9'h9) || (r_sys_run_step==9'hd) || (r_sys_run_step==9'h11) || (r_sys_run_step==9'h15) || (r_sys_run_step==9'h19) || (r_sys_run_step==9'h1d) || (r_sys_run_step==9'h21) || (r_sys_run_step==9'h25) || (r_sys_run_step==9'h29) || (r_sys_run_step==9'h2d) || (r_sys_run_step==9'h31) || (r_sys_run_step==9'h35) || (r_sys_run_step==9'h39) || (r_sys_run_step==9'h3d) || (r_sys_run_step==9'h41) || (r_sys_run_step==9'h45) || (r_sys_run_step==9'h49) || (r_sys_run_step==9'h4d) || (r_sys_run_step==9'h51) || (r_sys_run_step==9'h55) || (r_sys_run_step==9'h59) || (r_sys_run_step==9'h5d) || (r_sys_run_step==9'h61) || (r_sys_run_step==9'h65) || (r_sys_run_step==9'h69) || (r_sys_run_step==9'h6d) || (r_sys_run_step==9'h71) || (r_sys_run_step==9'h75) || (r_sys_run_step==9'h79) || (r_sys_run_step==9'h7d) || (r_sys_run_step==9'h81) || (r_sys_run_step==9'h85) || (r_sys_run_step==9'h89) || (r_sys_run_step==9'h8d) || (r_sys_run_step==9'h91) || (r_sys_run_step==9'h95) || (r_sys_run_step==9'h99) || (r_sys_run_step==9'h9d) || (r_sys_run_step==9'ha1) || (r_sys_run_step==9'ha5) || (r_sys_run_step==9'ha9) || (r_sys_run_step==9'had) || (r_sys_run_step==9'hb1) || (r_sys_run_step==9'hb5) || (r_sys_run_step==9'hb9) || (r_sys_run_step==9'hbd) || (r_sys_run_step==9'hc1) || (r_sys_run_step==9'hc5) || (r_sys_run_step==9'hc9) || (r_sys_run_step==9'hcd) || (r_sys_run_step==9'hd1) || (r_sys_run_step==9'hd5) || (r_sys_run_step==9'hd9) || (r_sys_run_step==9'hdd) || (r_sys_run_step==9'he1) || (r_sys_run_step==9'he5) || (r_sys_run_step==9'he9) || (r_sys_run_step==9'hed) || (r_sys_run_step==9'hf1) || (r_sys_run_step==9'hf5) || (r_sys_run_step==9'hf9) || (r_sys_run_step==9'hfd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp791[8:0] );

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2365[8:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2299[8:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2377[8:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2341[8:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2275[8:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2287[8:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2323[8:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2293[8:0] );

									end
									else
									if((r_sys_run_step==9'h1) || (r_sys_run_step==9'h16)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2269[8:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2305[8:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2383[8:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2347[8:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2371[8:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2281[8:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2335[8:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2353[8:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2317[8:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2311[8:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2359[8:0] );

									end
									else
									if((r_sys_run_step==9'h0) || (r_sys_run_step==9'h15)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2263[8:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2329[8:0] );

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2436[8:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2448[8:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2418[8:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2466[8:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2520[8:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2424[8:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2430[8:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2490[8:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2460[8:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2508[8:0] );

									end
									else
									if((r_sys_run_step==9'h0) || (r_sys_run_step==9'h15)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2406[8:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2496[8:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2514[8:0] );

									end
									else
									if((r_sys_run_step==9'h1) || (r_sys_run_step==9'h16)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2412[8:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2442[8:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2454[8:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2526[8:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2478[8:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2502[8:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2472[8:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2484[8:0] );

									end
								end

							endcase
						end

						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2578[8:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2599[8:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2606[8:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2571[8:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2653[8:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2623[8:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2633[8:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2550[8:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2643[8:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2585[8:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2618[8:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2658[8:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2648[8:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2628[8:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2557[8:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2613[8:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2592[8:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2638[8:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2564[8:0] );

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2737[8:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2747[8:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2767[8:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2676[8:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2772[8:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2697[8:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2732[8:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2718[8:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2669[8:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2683[8:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2742[8:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2711[8:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2704[8:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2725[8:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2757[8:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2762[8:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2777[8:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2690[8:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2752[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h3f)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp16;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h2) || (r_sys_run_step==9'h6) || (r_sys_run_step==9'ha) || (r_sys_run_step==9'he) || (r_sys_run_step==9'h12) || (r_sys_run_step==9'h16) || (r_sys_run_step==9'h1a) || (r_sys_run_step==9'h1e) || (r_sys_run_step==9'h22) || (r_sys_run_step==9'h26) || (r_sys_run_step==9'h2a) || (r_sys_run_step==9'h2e) || (r_sys_run_step==9'h32) || (r_sys_run_step==9'h36) || (r_sys_run_step==9'h3a) || (r_sys_run_step==9'h3e) || (r_sys_run_step==9'h42) || (r_sys_run_step==9'h46) || (r_sys_run_step==9'h4a) || (r_sys_run_step==9'h4e) || (r_sys_run_step==9'h52) || (r_sys_run_step==9'h56) || (r_sys_run_step==9'h5a) || (r_sys_run_step==9'h5e) || (r_sys_run_step==9'h62) || (r_sys_run_step==9'h66) || (r_sys_run_step==9'h6a) || (r_sys_run_step==9'h6e) || (r_sys_run_step==9'h72) || (r_sys_run_step==9'h76) || (r_sys_run_step==9'h7a) || (r_sys_run_step==9'h7e) || (r_sys_run_step==9'h82) || (r_sys_run_step==9'h86) || (r_sys_run_step==9'h8a) || (r_sys_run_step==9'h8e) || (r_sys_run_step==9'h92) || (r_sys_run_step==9'h96) || (r_sys_run_step==9'h9a) || (r_sys_run_step==9'h9e) || (r_sys_run_step==9'ha2) || (r_sys_run_step==9'ha6) || (r_sys_run_step==9'haa) || (r_sys_run_step==9'hae) || (r_sys_run_step==9'hb2) || (r_sys_run_step==9'hb6) || (r_sys_run_step==9'hba) || (r_sys_run_step==9'hbe) || (r_sys_run_step==9'hc2) || (r_sys_run_step==9'hc6) || (r_sys_run_step==9'hca) || (r_sys_run_step==9'hce) || (r_sys_run_step==9'hd2) || (r_sys_run_step==9'hd6) || (r_sys_run_step==9'hda) || (r_sys_run_step==9'hde) || (r_sys_run_step==9'he2) || (r_sys_run_step==9'he6) || (r_sys_run_step==9'hea) || (r_sys_run_step==9'hee) || (r_sys_run_step==9'hf2) || (r_sys_run_step==9'hf6) || (r_sys_run_step==9'hfa) || (r_sys_run_step==9'hfe)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp799;

									end
									else
									if((r_sys_run_step==9'h1) || (r_sys_run_step==9'h3) || (r_sys_run_step==9'h5) || (r_sys_run_step==9'h7) || (r_sys_run_step==9'h9) || (r_sys_run_step==9'hb) || (r_sys_run_step==9'hd) || (r_sys_run_step==9'hf) || (r_sys_run_step==9'h11) || (r_sys_run_step==9'h13) || (r_sys_run_step==9'h15) || (r_sys_run_step==9'h17) || (r_sys_run_step==9'h19) || (r_sys_run_step==9'h1b) || (r_sys_run_step==9'h1d) || (r_sys_run_step==9'h1f) || (r_sys_run_step==9'h21) || (r_sys_run_step==9'h23) || (r_sys_run_step==9'h25) || (r_sys_run_step==9'h27) || (r_sys_run_step==9'h29) || (r_sys_run_step==9'h2b) || (r_sys_run_step==9'h2d) || (r_sys_run_step==9'h2f) || (r_sys_run_step==9'h31) || (r_sys_run_step==9'h33) || (r_sys_run_step==9'h35) || (r_sys_run_step==9'h37) || (r_sys_run_step==9'h39) || (r_sys_run_step==9'h3b) || (r_sys_run_step==9'h3d) || (r_sys_run_step==9'h3f) || (r_sys_run_step==9'h41) || (r_sys_run_step==9'h43) || (r_sys_run_step==9'h45) || (r_sys_run_step==9'h47) || (r_sys_run_step==9'h49) || (r_sys_run_step==9'h4b) || (r_sys_run_step==9'h4d) || (r_sys_run_step==9'h4f) || (r_sys_run_step==9'h51) || (r_sys_run_step==9'h53) || (r_sys_run_step==9'h55) || (r_sys_run_step==9'h57) || (r_sys_run_step==9'h59) || (r_sys_run_step==9'h5b) || (r_sys_run_step==9'h5d) || (r_sys_run_step==9'h5f) || (r_sys_run_step==9'h61) || (r_sys_run_step==9'h63) || (r_sys_run_step==9'h65) || (r_sys_run_step==9'h67) || (r_sys_run_step==9'h69) || (r_sys_run_step==9'h6b) || (r_sys_run_step==9'h6d) || (r_sys_run_step==9'h6f) || (r_sys_run_step==9'h71) || (r_sys_run_step==9'h73) || (r_sys_run_step==9'h75) || (r_sys_run_step==9'h77) || (r_sys_run_step==9'h79) || (r_sys_run_step==9'h7b) || (r_sys_run_step==9'h7d) || (r_sys_run_step==9'h7f) || (r_sys_run_step==9'h81) || (r_sys_run_step==9'h83) || (r_sys_run_step==9'h85) || (r_sys_run_step==9'h87) || (r_sys_run_step==9'h89) || (r_sys_run_step==9'h8b) || (r_sys_run_step==9'h8d) || (r_sys_run_step==9'h8f) || (r_sys_run_step==9'h91) || (r_sys_run_step==9'h93) || (r_sys_run_step==9'h95) || (r_sys_run_step==9'h97) || (r_sys_run_step==9'h99) || (r_sys_run_step==9'h9b) || (r_sys_run_step==9'h9d) || (r_sys_run_step==9'h9f) || (r_sys_run_step==9'ha1) || (r_sys_run_step==9'ha3) || (r_sys_run_step==9'ha5) || (r_sys_run_step==9'ha7) || (r_sys_run_step==9'ha9) || (r_sys_run_step==9'hab) || (r_sys_run_step==9'had) || (r_sys_run_step==9'haf) || (r_sys_run_step==9'hb1) || (r_sys_run_step==9'hb3) || (r_sys_run_step==9'hb5) || (r_sys_run_step==9'hb7) || (r_sys_run_step==9'hb9) || (r_sys_run_step==9'hbb) || (r_sys_run_step==9'hbd) || (r_sys_run_step==9'hbf) || (r_sys_run_step==9'hc1) || (r_sys_run_step==9'hc3) || (r_sys_run_step==9'hc5) || (r_sys_run_step==9'hc7) || (r_sys_run_step==9'hc9) || (r_sys_run_step==9'hcb) || (r_sys_run_step==9'hcd) || (r_sys_run_step==9'hcf) || (r_sys_run_step==9'hd1) || (r_sys_run_step==9'hd3) || (r_sys_run_step==9'hd5) || (r_sys_run_step==9'hd7) || (r_sys_run_step==9'hd9) || (r_sys_run_step==9'hdb) || (r_sys_run_step==9'hdd) || (r_sys_run_step==9'hdf) || (r_sys_run_step==9'he1) || (r_sys_run_step==9'he3) || (r_sys_run_step==9'he5) || (r_sys_run_step==9'he7) || (r_sys_run_step==9'he9) || (r_sys_run_step==9'heb) || (r_sys_run_step==9'hed) || (r_sys_run_step==9'hef) || (r_sys_run_step==9'hf1) || (r_sys_run_step==9'hf3) || (r_sys_run_step==9'hf5) || (r_sys_run_step==9'hf7) || (r_sys_run_step==9'hf9) || (r_sys_run_step==9'hfb) || (r_sys_run_step==9'hfd) || (r_sys_run_step==9'hff)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp794;

									end
									else
									if((r_sys_run_step==9'h0) || (r_sys_run_step==9'h4) || (r_sys_run_step==9'h8) || (r_sys_run_step==9'hc) || (r_sys_run_step==9'h10) || (r_sys_run_step==9'h14) || (r_sys_run_step==9'h18) || (r_sys_run_step==9'h1c) || (r_sys_run_step==9'h20) || (r_sys_run_step==9'h24) || (r_sys_run_step==9'h28) || (r_sys_run_step==9'h2c) || (r_sys_run_step==9'h30) || (r_sys_run_step==9'h34) || (r_sys_run_step==9'h38) || (r_sys_run_step==9'h3c) || (r_sys_run_step==9'h40) || (r_sys_run_step==9'h44) || (r_sys_run_step==9'h48) || (r_sys_run_step==9'h4c) || (r_sys_run_step==9'h50) || (r_sys_run_step==9'h54) || (r_sys_run_step==9'h58) || (r_sys_run_step==9'h5c) || (r_sys_run_step==9'h60) || (r_sys_run_step==9'h64) || (r_sys_run_step==9'h68) || (r_sys_run_step==9'h6c) || (r_sys_run_step==9'h70) || (r_sys_run_step==9'h74) || (r_sys_run_step==9'h78) || (r_sys_run_step==9'h7c) || (r_sys_run_step==9'h80) || (r_sys_run_step==9'h84) || (r_sys_run_step==9'h88) || (r_sys_run_step==9'h8c) || (r_sys_run_step==9'h90) || (r_sys_run_step==9'h94) || (r_sys_run_step==9'h98) || (r_sys_run_step==9'h9c) || (r_sys_run_step==9'ha0) || (r_sys_run_step==9'ha4) || (r_sys_run_step==9'ha8) || (r_sys_run_step==9'hac) || (r_sys_run_step==9'hb0) || (r_sys_run_step==9'hb4) || (r_sys_run_step==9'hb8) || (r_sys_run_step==9'hbc) || (r_sys_run_step==9'hc0) || (r_sys_run_step==9'hc4) || (r_sys_run_step==9'hc8) || (r_sys_run_step==9'hcc) || (r_sys_run_step==9'hd0) || (r_sys_run_step==9'hd4) || (r_sys_run_step==9'hd8) || (r_sys_run_step==9'hdc) || (r_sys_run_step==9'he0) || (r_sys_run_step==9'he4) || (r_sys_run_step==9'he8) || (r_sys_run_step==9'hec) || (r_sys_run_step==9'hf0) || (r_sys_run_step==9'hf4) || (r_sys_run_step==9'hf8) || (r_sys_run_step==9'hfc)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp789;

									end
								end

							endcase
						end

						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==9'hb) || (r_sys_run_step==9'h14)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp7_float;

									end
									else
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'ha)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp2552;

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp0_float;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==9'hb) || (r_sys_run_step==9'h14)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp8_float;

									end
									else
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'ha)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp2671;

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp0_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h3f)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'hff)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h16)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h16)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h14)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h14)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h36: begin
							r_fld_u_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_uu_1_addr_1 <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h3f)) begin
										r_fld_uu_1_addr_1 <= $signed( w_sys_tmp18[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h3f)) begin
										r_fld_uu_1_datain_1 <= w_sys_tmp16;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_uu_1_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h3f)) begin
										r_fld_uu_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h36: begin
							r_fld_uu_1_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h4: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_6 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_6 <= w_sys_tmp8;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_6 <= w_sys_tmp2258;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_run_k_6 <= w_sys_tmp2400;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_6 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_run_k_6 <= w_sys_tmp2543;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_6 <= w_sys_tmp2544;

									end
								end

							endcase
						end

						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_run_k_6 <= w_sys_tmp2662;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_6 <= w_sys_tmp2663;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_run_k_6 <= w_sys_tmp2781;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_j_7 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h3f)) begin
										r_run_j_7 <= w_sys_tmp23;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_j_7 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0) || (r_sys_run_step==9'h4) || (r_sys_run_step==9'h8) || (r_sys_run_step==9'hc) || (r_sys_run_step==9'h10) || (r_sys_run_step==9'h14) || (r_sys_run_step==9'h18) || (r_sys_run_step==9'h1c) || (r_sys_run_step==9'h20) || (r_sys_run_step==9'h24) || (r_sys_run_step==9'h28) || (r_sys_run_step==9'h2c) || (r_sys_run_step==9'h30) || (r_sys_run_step==9'h34) || (r_sys_run_step==9'h38) || (r_sys_run_step==9'h3c) || (r_sys_run_step==9'h40) || (r_sys_run_step==9'h44) || (r_sys_run_step==9'h48) || (r_sys_run_step==9'h4c) || (r_sys_run_step==9'h50) || (r_sys_run_step==9'h54) || (r_sys_run_step==9'h58) || (r_sys_run_step==9'h5c) || (r_sys_run_step==9'h60) || (r_sys_run_step==9'h64) || (r_sys_run_step==9'h68) || (r_sys_run_step==9'h6c) || (r_sys_run_step==9'h70) || (r_sys_run_step==9'h74) || (r_sys_run_step==9'h78) || (r_sys_run_step==9'h7c) || (r_sys_run_step==9'h80) || (r_sys_run_step==9'h84) || (r_sys_run_step==9'h88) || (r_sys_run_step==9'h8c) || (r_sys_run_step==9'h90) || (r_sys_run_step==9'h94) || (r_sys_run_step==9'h98) || (r_sys_run_step==9'h9c) || (r_sys_run_step==9'ha0) || (r_sys_run_step==9'ha4) || (r_sys_run_step==9'ha8) || (r_sys_run_step==9'hac) || (r_sys_run_step==9'hb0) || (r_sys_run_step==9'hb4) || (r_sys_run_step==9'hb8) || (r_sys_run_step==9'hbc) || (r_sys_run_step==9'hc0) || (r_sys_run_step==9'hc4) || (r_sys_run_step==9'hc8) || (r_sys_run_step==9'hcc) || (r_sys_run_step==9'hd0) || (r_sys_run_step==9'hd4) || (r_sys_run_step==9'hd8) || (r_sys_run_step==9'hdc) || (r_sys_run_step==9'he0) || (r_sys_run_step==9'he4) || (r_sys_run_step==9'he8) || (r_sys_run_step==9'hec) || (r_sys_run_step==9'hf0) || (r_sys_run_step==9'hf4) || (r_sys_run_step==9'hf8) || (r_sys_run_step==9'hfc)) begin
										r_run_j_7 <= w_sys_tmp808;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_n_8 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_n_8 <= w_sys_tmp782;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_mx_9 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_my_10 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_nlast_11 <= w_sys_tmp5;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_dx_12 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_dy_13 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy0_j_14 <= r_run_j_7;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h3f)) begin
										r_run_copy0_j_14 <= w_sys_tmp22;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy0_j_15 <= r_run_j_7;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h3) || (r_sys_run_step==9'h7) || (r_sys_run_step==9'hb) || (r_sys_run_step==9'hf) || (r_sys_run_step==9'h13) || (r_sys_run_step==9'h17) || (r_sys_run_step==9'h1b) || (r_sys_run_step==9'h1f) || (r_sys_run_step==9'h23) || (r_sys_run_step==9'h27) || (r_sys_run_step==9'h2b) || (r_sys_run_step==9'h2f) || (r_sys_run_step==9'h33) || (r_sys_run_step==9'h37) || (r_sys_run_step==9'h3b) || (r_sys_run_step==9'h3f) || (r_sys_run_step==9'h43) || (r_sys_run_step==9'h47) || (r_sys_run_step==9'h4b) || (r_sys_run_step==9'h4f) || (r_sys_run_step==9'h53) || (r_sys_run_step==9'h57) || (r_sys_run_step==9'h5b) || (r_sys_run_step==9'h5f) || (r_sys_run_step==9'h63) || (r_sys_run_step==9'h67) || (r_sys_run_step==9'h6b) || (r_sys_run_step==9'h6f) || (r_sys_run_step==9'h73) || (r_sys_run_step==9'h77) || (r_sys_run_step==9'h7b) || (r_sys_run_step==9'h7f) || (r_sys_run_step==9'h83) || (r_sys_run_step==9'h87) || (r_sys_run_step==9'h8b) || (r_sys_run_step==9'h8f) || (r_sys_run_step==9'h93) || (r_sys_run_step==9'h97) || (r_sys_run_step==9'h9b) || (r_sys_run_step==9'h9f) || (r_sys_run_step==9'ha3) || (r_sys_run_step==9'ha7) || (r_sys_run_step==9'hab) || (r_sys_run_step==9'haf) || (r_sys_run_step==9'hb3) || (r_sys_run_step==9'hb7) || (r_sys_run_step==9'hbb) || (r_sys_run_step==9'hbf) || (r_sys_run_step==9'hc3) || (r_sys_run_step==9'hc7) || (r_sys_run_step==9'hcb) || (r_sys_run_step==9'hcf) || (r_sys_run_step==9'hd3) || (r_sys_run_step==9'hd7) || (r_sys_run_step==9'hdb) || (r_sys_run_step==9'hdf) || (r_sys_run_step==9'he3) || (r_sys_run_step==9'he7) || (r_sys_run_step==9'heb) || (r_sys_run_step==9'hef) || (r_sys_run_step==9'hf3) || (r_sys_run_step==9'hf7) || (r_sys_run_step==9'hfb) || (r_sys_run_step==9'hff)) begin
										r_run_copy0_j_15 <= w_sys_tmp805;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy1_j_16 <= r_run_j_7;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h2) || (r_sys_run_step==9'h6) || (r_sys_run_step==9'ha) || (r_sys_run_step==9'he) || (r_sys_run_step==9'h12) || (r_sys_run_step==9'h16) || (r_sys_run_step==9'h1a) || (r_sys_run_step==9'h1e) || (r_sys_run_step==9'h22) || (r_sys_run_step==9'h26) || (r_sys_run_step==9'h2a) || (r_sys_run_step==9'h2e) || (r_sys_run_step==9'h32) || (r_sys_run_step==9'h36) || (r_sys_run_step==9'h3a) || (r_sys_run_step==9'h3e) || (r_sys_run_step==9'h42) || (r_sys_run_step==9'h46) || (r_sys_run_step==9'h4a) || (r_sys_run_step==9'h4e) || (r_sys_run_step==9'h52) || (r_sys_run_step==9'h56) || (r_sys_run_step==9'h5a) || (r_sys_run_step==9'h5e) || (r_sys_run_step==9'h62) || (r_sys_run_step==9'h66) || (r_sys_run_step==9'h6a) || (r_sys_run_step==9'h6e) || (r_sys_run_step==9'h72) || (r_sys_run_step==9'h76) || (r_sys_run_step==9'h7a) || (r_sys_run_step==9'h7e) || (r_sys_run_step==9'h82) || (r_sys_run_step==9'h86) || (r_sys_run_step==9'h8a) || (r_sys_run_step==9'h8e) || (r_sys_run_step==9'h92) || (r_sys_run_step==9'h96) || (r_sys_run_step==9'h9a) || (r_sys_run_step==9'h9e) || (r_sys_run_step==9'ha2) || (r_sys_run_step==9'ha6) || (r_sys_run_step==9'haa) || (r_sys_run_step==9'hae) || (r_sys_run_step==9'hb2) || (r_sys_run_step==9'hb6) || (r_sys_run_step==9'hba) || (r_sys_run_step==9'hbe) || (r_sys_run_step==9'hc2) || (r_sys_run_step==9'hc6) || (r_sys_run_step==9'hca) || (r_sys_run_step==9'hce) || (r_sys_run_step==9'hd2) || (r_sys_run_step==9'hd6) || (r_sys_run_step==9'hda) || (r_sys_run_step==9'hde) || (r_sys_run_step==9'he2) || (r_sys_run_step==9'he6) || (r_sys_run_step==9'hea) || (r_sys_run_step==9'hee) || (r_sys_run_step==9'hf2) || (r_sys_run_step==9'hf6) || (r_sys_run_step==9'hfa) || (r_sys_run_step==9'hfe)) begin
										r_run_copy1_j_16 <= w_sys_tmp806;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy2_j_17 <= r_run_j_7;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h1) || (r_sys_run_step==9'h5) || (r_sys_run_step==9'h9) || (r_sys_run_step==9'hd) || (r_sys_run_step==9'h11) || (r_sys_run_step==9'h15) || (r_sys_run_step==9'h19) || (r_sys_run_step==9'h1d) || (r_sys_run_step==9'h21) || (r_sys_run_step==9'h25) || (r_sys_run_step==9'h29) || (r_sys_run_step==9'h2d) || (r_sys_run_step==9'h31) || (r_sys_run_step==9'h35) || (r_sys_run_step==9'h39) || (r_sys_run_step==9'h3d) || (r_sys_run_step==9'h41) || (r_sys_run_step==9'h45) || (r_sys_run_step==9'h49) || (r_sys_run_step==9'h4d) || (r_sys_run_step==9'h51) || (r_sys_run_step==9'h55) || (r_sys_run_step==9'h59) || (r_sys_run_step==9'h5d) || (r_sys_run_step==9'h61) || (r_sys_run_step==9'h65) || (r_sys_run_step==9'h69) || (r_sys_run_step==9'h6d) || (r_sys_run_step==9'h71) || (r_sys_run_step==9'h75) || (r_sys_run_step==9'h79) || (r_sys_run_step==9'h7d) || (r_sys_run_step==9'h81) || (r_sys_run_step==9'h85) || (r_sys_run_step==9'h89) || (r_sys_run_step==9'h8d) || (r_sys_run_step==9'h91) || (r_sys_run_step==9'h95) || (r_sys_run_step==9'h99) || (r_sys_run_step==9'h9d) || (r_sys_run_step==9'ha1) || (r_sys_run_step==9'ha5) || (r_sys_run_step==9'ha9) || (r_sys_run_step==9'had) || (r_sys_run_step==9'hb1) || (r_sys_run_step==9'hb5) || (r_sys_run_step==9'hb9) || (r_sys_run_step==9'hbd) || (r_sys_run_step==9'hc1) || (r_sys_run_step==9'hc5) || (r_sys_run_step==9'hc9) || (r_sys_run_step==9'hcd) || (r_sys_run_step==9'hd1) || (r_sys_run_step==9'hd5) || (r_sys_run_step==9'hd9) || (r_sys_run_step==9'hdd) || (r_sys_run_step==9'he1) || (r_sys_run_step==9'he5) || (r_sys_run_step==9'he9) || (r_sys_run_step==9'hed) || (r_sys_run_step==9'hf1) || (r_sys_run_step==9'hf5) || (r_sys_run_step==9'hf9) || (r_sys_run_step==9'hfd)) begin
										r_run_copy2_j_17 <= w_sys_tmp807;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp2299[8:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp2275[8:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp2281[8:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp2323[8:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp2287[8:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp2317[8:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp2311[8:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp2293[8:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp2329[8:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp2269[8:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp2263[8:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp2305[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'hd)) begin
										r_sub03_u_datain <= w_sys_tmp2265;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'hd)) begin
										r_sub03_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h36: begin
							r_sub03_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2737[8:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2742[8:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2747[8:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2767[8:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2757[8:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2772[8:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2732[8:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2762[8:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2777[8:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2752[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h9)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h36: begin
							r_sub03_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h16)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp2383[8:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp2365[8:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp2377[8:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp2347[8:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp2341[8:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp2371[8:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp2335[8:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp2353[8:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp2269[8:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp2263[8:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp2359[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'he<=r_sys_run_step && r_sys_run_step<=9'h18)) begin
										r_sub02_u_datain <= w_sys_tmp2265;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'he<=r_sys_run_step && r_sys_run_step<=9'h18)) begin
										r_sub02_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h36: begin
							r_sub02_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2672[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h36: begin
							r_sub02_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h26: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp2448[8:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp2436[8:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp2418[8:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp2466[8:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp2442[8:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp2424[8:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp2412[8:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp2454[8:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp2430[8:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp2460[8:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp2472[8:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp2406[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'hd)) begin
										r_sub01_u_datain <= w_sys_tmp2408;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'hd)) begin
										r_sub01_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h36: begin
							r_sub01_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2618[8:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2658[8:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2648[8:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2628[8:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2613[8:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2653[8:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2623[8:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2633[8:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2638[8:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2643[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h9)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h36: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h26: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp2496[8:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp2520[8:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp2514[8:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp2412[8:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp2526[8:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp2490[8:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp2478[8:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp2406[8:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp2508[8:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp2502[8:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp2484[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'he<=r_sys_run_step && r_sys_run_step<=9'h18)) begin
										r_sub00_u_datain <= w_sys_tmp2408;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'he<=r_sys_run_step && r_sys_run_step<=9'h18)) begin
										r_sub00_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h36: begin
							r_sub00_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp2553[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h8)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h36: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp0_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp0_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp1_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp1_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp2_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp2_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp3_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp3_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp4_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp4_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp5_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp5_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp6_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp6_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp7_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp7_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h2) || (r_sys_run_step==9'hb)) begin
										r_sys_tmp8_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==9'h2) || (r_sys_run_step==9'hb)) begin
										r_sys_tmp8_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
