/*
TimeStamp:	2016/9/15		15:58
*/


module c1_test(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy	
);

	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 5:0] r_sys_run_phase;
	reg         [ 1:0] r_sys_run_stage;
	reg         [ 6:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 1:0] w_sys_run_stage_p1;
	wire        [ 6:0] w_sys_run_step_p1;
	wire signed [ 8:0] w_fld_u_0_addr_0;
	wire        [31:0] w_fld_u_0_datain_0;
	wire        [31:0] w_fld_u_0_dataout_0;
	wire               w_fld_u_0_r_w_0;
	wire               w_fld_u_0_ce_0;
	reg  signed [ 8:0] r_fld_u_0_addr_1;
	reg         [31:0] r_fld_u_0_datain_1;
	wire        [31:0] w_fld_u_0_dataout_1;
	reg                r_fld_u_0_r_w_1;
	wire               w_fld_u_0_ce_1;
	wire signed [ 8:0] w_fld_uu_1_addr_0;
	wire        [31:0] w_fld_uu_1_datain_0;
	wire        [31:0] w_fld_uu_1_dataout_0;
	wire               w_fld_uu_1_r_w_0;
	wire               w_fld_uu_1_ce_0;
	reg  signed [ 8:0] r_fld_uu_1_addr_1;
	reg         [31:0] r_fld_uu_1_datain_1;
	wire        [31:0] w_fld_uu_1_dataout_1;
	reg                r_fld_uu_1_r_w_1;
	wire               w_fld_uu_1_ce_1;
	wire signed [ 8:0] w_fld_q_2_addr_0;
	wire        [31:0] w_fld_q_2_datain_0;
	wire        [31:0] w_fld_q_2_dataout_0;
	wire               w_fld_q_2_r_w_0;
	wire               w_fld_q_2_ce_0;
	reg  signed [ 8:0] r_fld_q_2_addr_1;
	reg         [31:0] r_fld_q_2_datain_1;
	wire        [31:0] w_fld_q_2_dataout_1;
	reg                r_fld_q_2_r_w_1;
	wire               w_fld_q_2_ce_1;
	reg  signed [31:0] r_run_k_5;
	reg  signed [31:0] r_run_j_6;
	reg  signed [31:0] r_run_n_7;
	reg  signed [31:0] r_run_mx_8;
	reg  signed [31:0] r_run_my_9;
	reg  signed [31:0] r_run_nlast_10;
	reg         [31:0] r_run_dx_11;
	reg         [31:0] r_run_dy_12;
	reg  signed [31:0] r_run_copy0_j_13;
	reg  signed [31:0] r_run_copy0_j_14;
	reg  signed [31:0] r_run_copy1_j_15;
	reg  signed [31:0] r_run_copy2_j_16;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [ 8:0] w_sub01_u_addr;
	reg  signed [ 8:0] r_sub01_u_addr;
	wire        [31:0] w_sub01_u_datain;
	reg         [31:0] r_sub01_u_datain;
	wire        [31:0] w_sub01_u_dataout;
	wire               w_sub01_u_r_w;
	reg                r_sub01_u_r_w;
	wire signed [ 8:0] w_sub01_q_addr;
	reg  signed [ 8:0] r_sub01_q_addr;
	wire        [31:0] w_sub01_q_datain;
	reg         [31:0] r_sub01_q_datain;
	wire        [31:0] w_sub01_q_dataout;
	wire               w_sub01_q_r_w;
	reg                r_sub01_q_r_w;
	wire signed [ 8:0] w_sub01_result_addr;
	reg  signed [ 8:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [ 8:0] w_sub00_u_addr;
	reg  signed [ 8:0] r_sub00_u_addr;
	wire        [31:0] w_sub00_u_datain;
	reg         [31:0] r_sub00_u_datain;
	wire        [31:0] w_sub00_u_dataout;
	wire               w_sub00_u_r_w;
	reg                r_sub00_u_r_w;
	wire signed [ 8:0] w_sub00_q_addr;
	reg  signed [ 8:0] r_sub00_q_addr;
	wire        [31:0] w_sub00_q_datain;
	reg         [31:0] r_sub00_q_datain;
	wire        [31:0] w_sub00_q_dataout;
	wire               w_sub00_q_r_w;
	reg                r_sub00_q_r_w;
	wire signed [ 8:0] w_sub00_result_addr;
	reg  signed [ 8:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	wire signed [31:0] w_sys_tmp1;
	wire        [31:0] w_sys_tmp3;
	wire signed [31:0] w_sys_tmp5;
	wire               w_sys_tmp6;
	wire               w_sys_tmp7;
	wire signed [31:0] w_sys_tmp8;
	wire               w_sys_tmp9;
	wire               w_sys_tmp10;
	wire signed [31:0] w_sys_tmp13;
	wire signed [31:0] w_sys_tmp14;
	wire signed [31:0] w_sys_tmp15;
	wire        [31:0] w_sys_tmp16;
	wire signed [31:0] w_sys_tmp18;
	wire signed [31:0] w_sys_tmp19;
	wire signed [31:0] w_sys_tmp22;
	wire signed [31:0] w_sys_tmp23;
	wire               w_sys_tmp252;
	wire               w_sys_tmp253;
	wire signed [31:0] w_sys_tmp254;
	wire               w_sys_tmp255;
	wire               w_sys_tmp256;
	wire signed [31:0] w_sys_tmp259;
	wire signed [31:0] w_sys_tmp260;
	wire        [31:0] w_sys_tmp261;
	wire signed [31:0] w_sys_tmp263;
	wire signed [31:0] w_sys_tmp264;
	wire        [31:0] w_sys_tmp266;
	wire signed [31:0] w_sys_tmp268;
	wire signed [31:0] w_sys_tmp269;
	wire        [31:0] w_sys_tmp271;
	wire signed [31:0] w_sys_tmp273;
	wire signed [31:0] w_sys_tmp274;
	wire signed [31:0] w_sys_tmp277;
	wire signed [31:0] w_sys_tmp278;
	wire signed [31:0] w_sys_tmp279;
	wire signed [31:0] w_sys_tmp280;
	wire               w_sys_tmp718;
	wire               w_sys_tmp719;
	wire signed [31:0] w_sys_tmp720;
	wire signed [31:0] w_sys_tmp723;
	wire signed [31:0] w_sys_tmp724;
	wire        [31:0] w_sys_tmp725;
	wire signed [31:0] w_sys_tmp729;
	wire signed [31:0] w_sys_tmp730;
	wire signed [31:0] w_sys_tmp735;
	wire signed [31:0] w_sys_tmp736;
	wire signed [31:0] w_sys_tmp741;
	wire signed [31:0] w_sys_tmp742;
	wire signed [31:0] w_sys_tmp747;
	wire signed [31:0] w_sys_tmp748;
	wire signed [31:0] w_sys_tmp753;
	wire signed [31:0] w_sys_tmp754;
	wire signed [31:0] w_sys_tmp759;
	wire signed [31:0] w_sys_tmp760;
	wire signed [31:0] w_sys_tmp765;
	wire signed [31:0] w_sys_tmp766;
	wire signed [31:0] w_sys_tmp771;
	wire signed [31:0] w_sys_tmp772;
	wire signed [31:0] w_sys_tmp777;
	wire signed [31:0] w_sys_tmp778;
	wire signed [31:0] w_sys_tmp783;
	wire signed [31:0] w_sys_tmp784;
	wire signed [31:0] w_sys_tmp789;
	wire signed [31:0] w_sys_tmp790;
	wire signed [31:0] w_sys_tmp795;
	wire signed [31:0] w_sys_tmp796;
	wire signed [31:0] w_sys_tmp801;
	wire signed [31:0] w_sys_tmp802;
	wire signed [31:0] w_sys_tmp807;
	wire signed [31:0] w_sys_tmp808;
	wire signed [31:0] w_sys_tmp813;
	wire signed [31:0] w_sys_tmp814;
	wire signed [31:0] w_sys_tmp819;
	wire signed [31:0] w_sys_tmp820;
	wire signed [31:0] w_sys_tmp825;
	wire signed [31:0] w_sys_tmp826;
	wire signed [31:0] w_sys_tmp831;
	wire signed [31:0] w_sys_tmp832;
	wire signed [31:0] w_sys_tmp837;
	wire signed [31:0] w_sys_tmp838;
	wire signed [31:0] w_sys_tmp843;
	wire signed [31:0] w_sys_tmp844;
	wire signed [31:0] w_sys_tmp848;
	wire signed [31:0] w_sys_tmp849;
	wire               w_sys_tmp850;
	wire               w_sys_tmp851;
	wire signed [31:0] w_sys_tmp854;
	wire signed [31:0] w_sys_tmp855;
	wire        [31:0] w_sys_tmp856;
	wire signed [31:0] w_sys_tmp860;
	wire signed [31:0] w_sys_tmp861;
	wire signed [31:0] w_sys_tmp866;
	wire signed [31:0] w_sys_tmp867;
	wire signed [31:0] w_sys_tmp872;
	wire signed [31:0] w_sys_tmp873;
	wire signed [31:0] w_sys_tmp878;
	wire signed [31:0] w_sys_tmp879;
	wire signed [31:0] w_sys_tmp884;
	wire signed [31:0] w_sys_tmp885;
	wire signed [31:0] w_sys_tmp890;
	wire signed [31:0] w_sys_tmp891;
	wire signed [31:0] w_sys_tmp896;
	wire signed [31:0] w_sys_tmp897;
	wire signed [31:0] w_sys_tmp902;
	wire signed [31:0] w_sys_tmp903;
	wire signed [31:0] w_sys_tmp908;
	wire signed [31:0] w_sys_tmp909;
	wire signed [31:0] w_sys_tmp914;
	wire signed [31:0] w_sys_tmp915;
	wire signed [31:0] w_sys_tmp920;
	wire signed [31:0] w_sys_tmp921;
	wire signed [31:0] w_sys_tmp926;
	wire signed [31:0] w_sys_tmp927;
	wire signed [31:0] w_sys_tmp932;
	wire signed [31:0] w_sys_tmp933;
	wire signed [31:0] w_sys_tmp938;
	wire signed [31:0] w_sys_tmp939;
	wire signed [31:0] w_sys_tmp944;
	wire signed [31:0] w_sys_tmp945;
	wire signed [31:0] w_sys_tmp950;
	wire signed [31:0] w_sys_tmp951;
	wire signed [31:0] w_sys_tmp956;
	wire signed [31:0] w_sys_tmp957;
	wire signed [31:0] w_sys_tmp962;
	wire signed [31:0] w_sys_tmp963;
	wire signed [31:0] w_sys_tmp968;
	wire signed [31:0] w_sys_tmp969;
	wire signed [31:0] w_sys_tmp974;
	wire signed [31:0] w_sys_tmp975;
	wire signed [31:0] w_sys_tmp979;
	wire signed [31:0] w_sys_tmp980;
	wire               w_sys_tmp981;
	wire               w_sys_tmp982;
	wire signed [31:0] w_sys_tmp983;
	wire signed [31:0] w_sys_tmp986;
	wire signed [31:0] w_sys_tmp987;
	wire        [31:0] w_sys_tmp988;
	wire signed [31:0] w_sys_tmp992;
	wire signed [31:0] w_sys_tmp993;
	wire signed [31:0] w_sys_tmp998;
	wire signed [31:0] w_sys_tmp999;
	wire signed [31:0] w_sys_tmp1004;
	wire signed [31:0] w_sys_tmp1005;
	wire signed [31:0] w_sys_tmp1010;
	wire signed [31:0] w_sys_tmp1011;
	wire signed [31:0] w_sys_tmp1016;
	wire signed [31:0] w_sys_tmp1017;
	wire signed [31:0] w_sys_tmp1022;
	wire signed [31:0] w_sys_tmp1023;
	wire signed [31:0] w_sys_tmp1028;
	wire signed [31:0] w_sys_tmp1029;
	wire signed [31:0] w_sys_tmp1034;
	wire signed [31:0] w_sys_tmp1035;
	wire signed [31:0] w_sys_tmp1040;
	wire signed [31:0] w_sys_tmp1041;
	wire signed [31:0] w_sys_tmp1046;
	wire signed [31:0] w_sys_tmp1047;
	wire signed [31:0] w_sys_tmp1052;
	wire signed [31:0] w_sys_tmp1053;
	wire signed [31:0] w_sys_tmp1058;
	wire signed [31:0] w_sys_tmp1059;
	wire signed [31:0] w_sys_tmp1064;
	wire signed [31:0] w_sys_tmp1065;
	wire signed [31:0] w_sys_tmp1070;
	wire signed [31:0] w_sys_tmp1071;
	wire signed [31:0] w_sys_tmp1076;
	wire signed [31:0] w_sys_tmp1077;
	wire signed [31:0] w_sys_tmp1082;
	wire signed [31:0] w_sys_tmp1083;
	wire signed [31:0] w_sys_tmp1088;
	wire signed [31:0] w_sys_tmp1089;
	wire signed [31:0] w_sys_tmp1094;
	wire signed [31:0] w_sys_tmp1095;
	wire signed [31:0] w_sys_tmp1099;
	wire signed [31:0] w_sys_tmp1100;
	wire               w_sys_tmp1101;
	wire               w_sys_tmp1102;
	wire signed [31:0] w_sys_tmp1103;
	wire signed [31:0] w_sys_tmp1106;
	wire signed [31:0] w_sys_tmp1107;
	wire        [31:0] w_sys_tmp1108;
	wire signed [31:0] w_sys_tmp1112;
	wire signed [31:0] w_sys_tmp1113;
	wire signed [31:0] w_sys_tmp1118;
	wire signed [31:0] w_sys_tmp1119;
	wire signed [31:0] w_sys_tmp1124;
	wire signed [31:0] w_sys_tmp1125;
	wire signed [31:0] w_sys_tmp1130;
	wire signed [31:0] w_sys_tmp1131;
	wire signed [31:0] w_sys_tmp1136;
	wire signed [31:0] w_sys_tmp1137;
	wire signed [31:0] w_sys_tmp1142;
	wire signed [31:0] w_sys_tmp1143;
	wire signed [31:0] w_sys_tmp1148;
	wire signed [31:0] w_sys_tmp1149;
	wire signed [31:0] w_sys_tmp1154;
	wire signed [31:0] w_sys_tmp1155;
	wire signed [31:0] w_sys_tmp1160;
	wire signed [31:0] w_sys_tmp1161;
	wire signed [31:0] w_sys_tmp1166;
	wire signed [31:0] w_sys_tmp1167;
	wire signed [31:0] w_sys_tmp1172;
	wire signed [31:0] w_sys_tmp1173;
	wire signed [31:0] w_sys_tmp1178;
	wire signed [31:0] w_sys_tmp1179;
	wire signed [31:0] w_sys_tmp1184;
	wire signed [31:0] w_sys_tmp1185;
	wire signed [31:0] w_sys_tmp1190;
	wire signed [31:0] w_sys_tmp1191;
	wire signed [31:0] w_sys_tmp1196;
	wire signed [31:0] w_sys_tmp1197;
	wire signed [31:0] w_sys_tmp1202;
	wire signed [31:0] w_sys_tmp1203;
	wire signed [31:0] w_sys_tmp1208;
	wire signed [31:0] w_sys_tmp1209;
	wire signed [31:0] w_sys_tmp1214;
	wire signed [31:0] w_sys_tmp1215;
	wire signed [31:0] w_sys_tmp1219;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 2'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 7'h1);
	assign w_fld_u_0_addr_0 = 9'sh0;
	assign w_fld_u_0_datain_0 = 32'h0;
	assign w_fld_u_0_r_w_0 = 1'h0;
	assign w_fld_u_0_ce_0 = w_sys_ce;
	assign w_fld_u_0_ce_1 = w_sys_ce;
	assign w_fld_uu_1_addr_0 = 9'sh0;
	assign w_fld_uu_1_datain_0 = 32'h0;
	assign w_fld_uu_1_r_w_0 = 1'h0;
	assign w_fld_uu_1_ce_0 = w_sys_ce;
	assign w_fld_uu_1_ce_1 = w_sys_ce;
	assign w_fld_q_2_addr_0 = 9'sh0;
	assign w_fld_q_2_datain_0 = 32'h0;
	assign w_fld_q_2_r_w_0 = 1'h0;
	assign w_fld_q_2_ce_0 = w_sys_ce;
	assign w_fld_q_2_ce_1 = w_sys_ce;
	assign w_sub01_u_addr = ( (|r_sys_processing_methodID) ? r_sub01_u_addr : 9'sh0 ) ;
	assign w_sub01_u_datain = ( (|r_sys_processing_methodID) ? r_sub01_u_datain : 32'h0 ) ;
	assign w_sub01_u_r_w = ( (|r_sys_processing_methodID) ? r_sub01_u_r_w : 1'h0 ) ;
	assign w_sub01_q_addr = ( (|r_sys_processing_methodID) ? r_sub01_q_addr : 9'sh0 ) ;
	assign w_sub01_q_datain = ( (|r_sys_processing_methodID) ? r_sub01_q_datain : 32'h0 ) ;
	assign w_sub01_q_r_w = ( (|r_sys_processing_methodID) ? r_sub01_q_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 9'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub00_u_addr = ( (|r_sys_processing_methodID) ? r_sub00_u_addr : 9'sh0 ) ;
	assign w_sub00_u_datain = ( (|r_sys_processing_methodID) ? r_sub00_u_datain : 32'h0 ) ;
	assign w_sub00_u_r_w = ( (|r_sys_processing_methodID) ? r_sub00_u_r_w : 1'h0 ) ;
	assign w_sub00_q_addr = ( (|r_sys_processing_methodID) ? r_sub00_q_addr : 9'sh0 ) ;
	assign w_sub00_q_datain = ( (|r_sys_processing_methodID) ? r_sub00_q_datain : 32'h0 ) ;
	assign w_sub00_q_r_w = ( (|r_sys_processing_methodID) ? r_sub00_q_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 9'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh00000015;
	assign w_sys_tmp3 = 32'h3d4ccccd;
	assign w_sys_tmp5 = 32'sh00000190;
	assign w_sys_tmp6 = ( !w_sys_tmp7 );
	assign w_sys_tmp7 = (r_run_my_9 < r_run_k_5);
	assign w_sys_tmp8 = (r_run_k_5 + w_sys_intOne);
	assign w_sys_tmp9 = ( !w_sys_tmp10 );
	assign w_sys_tmp10 = (r_run_mx_8 < r_run_j_6);
	assign w_sys_tmp13 = (w_sys_tmp14 + r_run_k_5);
	assign w_sys_tmp14 = (r_run_j_6 * w_sys_tmp15);
	assign w_sys_tmp15 = 32'sh00000015;
	assign w_sys_tmp16 = 32'h0;
	assign w_sys_tmp18 = (w_sys_tmp19 + r_run_k_5);
	assign w_sys_tmp19 = (r_run_copy0_j_13 * w_sys_tmp15);
	assign w_sys_tmp22 = (r_run_copy0_j_13 + w_sys_intOne);
	assign w_sys_tmp23 = (r_run_j_6 + w_sys_intOne);
	assign w_sys_tmp252 = ( !w_sys_tmp253 );
	assign w_sys_tmp253 = (r_run_nlast_10 < r_run_n_7);
	assign w_sys_tmp254 = (r_run_n_7 + w_sys_intOne);
	assign w_sys_tmp255 = ( !w_sys_tmp256 );
	assign w_sys_tmp256 = (r_run_my_9 < r_run_j_6);
	assign w_sys_tmp259 = (w_sys_tmp260 + r_run_j_6);
	assign w_sys_tmp260 = 32'sh00000015;
	assign w_sys_tmp261 = 32'h3f000000;
	assign w_sys_tmp263 = (w_sys_tmp264 + r_run_copy2_j_16);
	assign w_sys_tmp264 = (r_run_mx_8 * w_sys_tmp260);
	assign w_sys_tmp266 = 32'h0;
	assign w_sys_tmp268 = (w_sys_tmp269 + w_sys_intOne);
	assign w_sys_tmp269 = (r_run_copy1_j_15 * w_sys_tmp260);
	assign w_sys_tmp271 = 32'h3f800000;
	assign w_sys_tmp273 = (w_sys_tmp274 + r_run_my_9);
	assign w_sys_tmp274 = (r_run_copy0_j_14 * w_sys_tmp260);
	assign w_sys_tmp277 = (r_run_copy0_j_14 + w_sys_intOne);
	assign w_sys_tmp278 = (r_run_copy1_j_15 + w_sys_intOne);
	assign w_sys_tmp279 = (r_run_copy2_j_16 + w_sys_intOne);
	assign w_sys_tmp280 = (r_run_j_6 + w_sys_intOne);
	assign w_sys_tmp718 = ( !w_sys_tmp719 );
	assign w_sys_tmp719 = (w_sys_tmp720 < r_run_k_5);
	assign w_sys_tmp720 = 32'sh0000000b;
	assign w_sys_tmp723 = (w_sys_tmp724 + r_run_k_5);
	assign w_sys_tmp724 = 32'sh00000015;
	assign w_sys_tmp725 = w_fld_u_0_dataout_1;
	assign w_sys_tmp729 = (w_sys_tmp730 + r_run_k_5);
	assign w_sys_tmp730 = 32'sh0000002a;
	assign w_sys_tmp735 = (w_sys_tmp736 + r_run_k_5);
	assign w_sys_tmp736 = 32'sh0000003f;
	assign w_sys_tmp741 = (w_sys_tmp742 + r_run_k_5);
	assign w_sys_tmp742 = 32'sh00000054;
	assign w_sys_tmp747 = (w_sys_tmp748 + r_run_k_5);
	assign w_sys_tmp748 = 32'sh00000069;
	assign w_sys_tmp753 = (w_sys_tmp754 + r_run_k_5);
	assign w_sys_tmp754 = 32'sh0000007e;
	assign w_sys_tmp759 = (w_sys_tmp760 + r_run_k_5);
	assign w_sys_tmp760 = 32'sh00000093;
	assign w_sys_tmp765 = (w_sys_tmp766 + r_run_k_5);
	assign w_sys_tmp766 = 32'sh000000a8;
	assign w_sys_tmp771 = (w_sys_tmp772 + r_run_k_5);
	assign w_sys_tmp772 = 32'sh000000bd;
	assign w_sys_tmp777 = (w_sys_tmp778 + r_run_k_5);
	assign w_sys_tmp778 = 32'sh000000d2;
	assign w_sys_tmp783 = (w_sys_tmp784 + r_run_k_5);
	assign w_sys_tmp784 = 32'sh000000e7;
	assign w_sys_tmp789 = (w_sys_tmp790 + r_run_k_5);
	assign w_sys_tmp790 = 32'sh000000fc;
	assign w_sys_tmp795 = (w_sys_tmp796 + r_run_k_5);
	assign w_sys_tmp796 = 32'sh00000111;
	assign w_sys_tmp801 = (w_sys_tmp802 + r_run_k_5);
	assign w_sys_tmp802 = 32'sh00000126;
	assign w_sys_tmp807 = (w_sys_tmp808 + r_run_k_5);
	assign w_sys_tmp808 = 32'sh0000013b;
	assign w_sys_tmp813 = (w_sys_tmp814 + r_run_k_5);
	assign w_sys_tmp814 = 32'sh00000150;
	assign w_sys_tmp819 = (w_sys_tmp820 + r_run_k_5);
	assign w_sys_tmp820 = 32'sh00000165;
	assign w_sys_tmp825 = (w_sys_tmp826 + r_run_k_5);
	assign w_sys_tmp826 = 32'sh0000017a;
	assign w_sys_tmp831 = (w_sys_tmp832 + r_run_k_5);
	assign w_sys_tmp832 = 32'sh0000018f;
	assign w_sys_tmp837 = (w_sys_tmp838 + r_run_k_5);
	assign w_sys_tmp838 = 32'sh000001a4;
	assign w_sys_tmp843 = (w_sys_tmp844 + r_run_k_5);
	assign w_sys_tmp844 = 32'sh000001b9;
	assign w_sys_tmp848 = (r_run_k_5 + w_sys_intOne);
	assign w_sys_tmp849 = 32'sh0000000a;
	assign w_sys_tmp850 = ( !w_sys_tmp851 );
	assign w_sys_tmp851 = (r_run_my_9 < r_run_k_5);
	assign w_sys_tmp854 = (w_sys_tmp855 + r_run_k_5);
	assign w_sys_tmp855 = 32'sh00000015;
	assign w_sys_tmp856 = w_fld_u_0_dataout_1;
	assign w_sys_tmp860 = (w_sys_tmp861 + r_run_k_5);
	assign w_sys_tmp861 = 32'sh0000002a;
	assign w_sys_tmp866 = (w_sys_tmp867 + r_run_k_5);
	assign w_sys_tmp867 = 32'sh0000003f;
	assign w_sys_tmp872 = (w_sys_tmp873 + r_run_k_5);
	assign w_sys_tmp873 = 32'sh00000054;
	assign w_sys_tmp878 = (w_sys_tmp879 + r_run_k_5);
	assign w_sys_tmp879 = 32'sh00000069;
	assign w_sys_tmp884 = (w_sys_tmp885 + r_run_k_5);
	assign w_sys_tmp885 = 32'sh0000007e;
	assign w_sys_tmp890 = (w_sys_tmp891 + r_run_k_5);
	assign w_sys_tmp891 = 32'sh00000093;
	assign w_sys_tmp896 = (w_sys_tmp897 + r_run_k_5);
	assign w_sys_tmp897 = 32'sh000000a8;
	assign w_sys_tmp902 = (w_sys_tmp903 + r_run_k_5);
	assign w_sys_tmp903 = 32'sh000000bd;
	assign w_sys_tmp908 = (w_sys_tmp909 + r_run_k_5);
	assign w_sys_tmp909 = 32'sh000000d2;
	assign w_sys_tmp914 = (w_sys_tmp915 + r_run_k_5);
	assign w_sys_tmp915 = 32'sh000000e7;
	assign w_sys_tmp920 = (w_sys_tmp921 + r_run_k_5);
	assign w_sys_tmp921 = 32'sh000000fc;
	assign w_sys_tmp926 = (w_sys_tmp927 + r_run_k_5);
	assign w_sys_tmp927 = 32'sh00000111;
	assign w_sys_tmp932 = (w_sys_tmp933 + r_run_k_5);
	assign w_sys_tmp933 = 32'sh00000126;
	assign w_sys_tmp938 = (w_sys_tmp939 + r_run_k_5);
	assign w_sys_tmp939 = 32'sh0000013b;
	assign w_sys_tmp944 = (w_sys_tmp945 + r_run_k_5);
	assign w_sys_tmp945 = 32'sh00000150;
	assign w_sys_tmp950 = (w_sys_tmp951 + r_run_k_5);
	assign w_sys_tmp951 = 32'sh00000165;
	assign w_sys_tmp956 = (w_sys_tmp957 + r_run_k_5);
	assign w_sys_tmp957 = 32'sh0000017a;
	assign w_sys_tmp962 = (w_sys_tmp963 + r_run_k_5);
	assign w_sys_tmp963 = 32'sh0000018f;
	assign w_sys_tmp968 = (w_sys_tmp969 + r_run_k_5);
	assign w_sys_tmp969 = 32'sh000001a4;
	assign w_sys_tmp974 = (w_sys_tmp975 + r_run_k_5);
	assign w_sys_tmp975 = 32'sh000001b9;
	assign w_sys_tmp979 = (r_run_k_5 + w_sys_intOne);
	assign w_sys_tmp980 = 32'sh00000002;
	assign w_sys_tmp981 = ( !w_sys_tmp982 );
	assign w_sys_tmp982 = (w_sys_tmp983 < r_run_k_5);
	assign w_sys_tmp983 = 32'sh0000000a;
	assign w_sys_tmp986 = (w_sys_tmp987 + r_run_k_5);
	assign w_sys_tmp987 = 32'sh0000002a;
	assign w_sys_tmp988 = w_sub00_result_dataout;
	assign w_sys_tmp992 = (w_sys_tmp993 + r_run_k_5);
	assign w_sys_tmp993 = 32'sh0000003f;
	assign w_sys_tmp998 = (w_sys_tmp999 + r_run_k_5);
	assign w_sys_tmp999 = 32'sh00000054;
	assign w_sys_tmp1004 = (w_sys_tmp1005 + r_run_k_5);
	assign w_sys_tmp1005 = 32'sh00000069;
	assign w_sys_tmp1010 = (w_sys_tmp1011 + r_run_k_5);
	assign w_sys_tmp1011 = 32'sh0000007e;
	assign w_sys_tmp1016 = (w_sys_tmp1017 + r_run_k_5);
	assign w_sys_tmp1017 = 32'sh00000093;
	assign w_sys_tmp1022 = (w_sys_tmp1023 + r_run_k_5);
	assign w_sys_tmp1023 = 32'sh000000a8;
	assign w_sys_tmp1028 = (w_sys_tmp1029 + r_run_k_5);
	assign w_sys_tmp1029 = 32'sh000000bd;
	assign w_sys_tmp1034 = (w_sys_tmp1035 + r_run_k_5);
	assign w_sys_tmp1035 = 32'sh000000d2;
	assign w_sys_tmp1040 = (w_sys_tmp1041 + r_run_k_5);
	assign w_sys_tmp1041 = 32'sh000000e7;
	assign w_sys_tmp1046 = (w_sys_tmp1047 + r_run_k_5);
	assign w_sys_tmp1047 = 32'sh000000fc;
	assign w_sys_tmp1052 = (w_sys_tmp1053 + r_run_k_5);
	assign w_sys_tmp1053 = 32'sh00000111;
	assign w_sys_tmp1058 = (w_sys_tmp1059 + r_run_k_5);
	assign w_sys_tmp1059 = 32'sh00000126;
	assign w_sys_tmp1064 = (w_sys_tmp1065 + r_run_k_5);
	assign w_sys_tmp1065 = 32'sh0000013b;
	assign w_sys_tmp1070 = (w_sys_tmp1071 + r_run_k_5);
	assign w_sys_tmp1071 = 32'sh00000150;
	assign w_sys_tmp1076 = (w_sys_tmp1077 + r_run_k_5);
	assign w_sys_tmp1077 = 32'sh00000165;
	assign w_sys_tmp1082 = (w_sys_tmp1083 + r_run_k_5);
	assign w_sys_tmp1083 = 32'sh0000017a;
	assign w_sys_tmp1088 = (w_sys_tmp1089 + r_run_k_5);
	assign w_sys_tmp1089 = 32'sh0000018f;
	assign w_sys_tmp1094 = (w_sys_tmp1095 + r_run_k_5);
	assign w_sys_tmp1095 = 32'sh000001a4;
	assign w_sys_tmp1099 = (r_run_k_5 + w_sys_intOne);
	assign w_sys_tmp1100 = 32'sh0000000b;
	assign w_sys_tmp1101 = ( !w_sys_tmp1102 );
	assign w_sys_tmp1102 = (w_sys_tmp1103 < r_run_k_5);
	assign w_sys_tmp1103 = 32'sh00000014;
	assign w_sys_tmp1106 = (w_sys_tmp1107 + r_run_k_5);
	assign w_sys_tmp1107 = 32'sh0000002a;
	assign w_sys_tmp1108 = w_sub01_result_dataout;
	assign w_sys_tmp1112 = (w_sys_tmp1113 + r_run_k_5);
	assign w_sys_tmp1113 = 32'sh0000003f;
	assign w_sys_tmp1118 = (w_sys_tmp1119 + r_run_k_5);
	assign w_sys_tmp1119 = 32'sh00000054;
	assign w_sys_tmp1124 = (w_sys_tmp1125 + r_run_k_5);
	assign w_sys_tmp1125 = 32'sh00000069;
	assign w_sys_tmp1130 = (w_sys_tmp1131 + r_run_k_5);
	assign w_sys_tmp1131 = 32'sh0000007e;
	assign w_sys_tmp1136 = (w_sys_tmp1137 + r_run_k_5);
	assign w_sys_tmp1137 = 32'sh00000093;
	assign w_sys_tmp1142 = (w_sys_tmp1143 + r_run_k_5);
	assign w_sys_tmp1143 = 32'sh000000a8;
	assign w_sys_tmp1148 = (w_sys_tmp1149 + r_run_k_5);
	assign w_sys_tmp1149 = 32'sh000000bd;
	assign w_sys_tmp1154 = (w_sys_tmp1155 + r_run_k_5);
	assign w_sys_tmp1155 = 32'sh000000d2;
	assign w_sys_tmp1160 = (w_sys_tmp1161 + r_run_k_5);
	assign w_sys_tmp1161 = 32'sh000000e7;
	assign w_sys_tmp1166 = (w_sys_tmp1167 + r_run_k_5);
	assign w_sys_tmp1167 = 32'sh000000fc;
	assign w_sys_tmp1172 = (w_sys_tmp1173 + r_run_k_5);
	assign w_sys_tmp1173 = 32'sh00000111;
	assign w_sys_tmp1178 = (w_sys_tmp1179 + r_run_k_5);
	assign w_sys_tmp1179 = 32'sh00000126;
	assign w_sys_tmp1184 = (w_sys_tmp1185 + r_run_k_5);
	assign w_sys_tmp1185 = 32'sh0000013b;
	assign w_sys_tmp1190 = (w_sys_tmp1191 + r_run_k_5);
	assign w_sys_tmp1191 = 32'sh00000150;
	assign w_sys_tmp1196 = (w_sys_tmp1197 + r_run_k_5);
	assign w_sys_tmp1197 = 32'sh00000165;
	assign w_sys_tmp1202 = (w_sys_tmp1203 + r_run_k_5);
	assign w_sys_tmp1203 = 32'sh0000017a;
	assign w_sys_tmp1208 = (w_sys_tmp1209 + r_run_k_5);
	assign w_sys_tmp1209 = 32'sh0000018f;
	assign w_sys_tmp1214 = (w_sys_tmp1215 + r_run_k_5);
	assign w_sys_tmp1215 = 32'sh000001a4;
	assign w_sys_tmp1219 = (r_run_k_5 + w_sys_intOne);


	subunder
		sub01_inst(
			.i_fld_q_1_addr_0 (w_sub01_q_addr),
			.i_fld_q_1_datain_0 (w_sub01_q_datain),
			.o_fld_q_1_dataout_0 (w_sub01_q_dataout),
			.i_fld_q_1_r_w_0 (w_sub01_q_r_w),
			.i_fld_result_2_addr_0 (w_sub01_result_addr),
			.i_fld_result_2_datain_0 (w_sub01_result_datain),
			.o_fld_result_2_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub01_result_r_w),
			.i_fld_u_0_addr_0 (w_sub01_u_addr),
			.i_fld_u_0_datain_0 (w_sub01_u_datain),
			.o_fld_u_0_dataout_0 (w_sub01_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub01_u_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	subup
		sub00_inst(
			.i_fld_q_1_addr_0 (w_sub00_q_addr),
			.i_fld_q_1_datain_0 (w_sub00_q_datain),
			.o_fld_q_1_dataout_0 (w_sub00_q_dataout),
			.i_fld_q_1_r_w_0 (w_sub00_q_r_w),
			.i_fld_result_2_addr_0 (w_sub00_result_addr),
			.i_fld_result_2_datain_0 (w_sub00_result_datain),
			.o_fld_result_2_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub00_result_r_w),
			.i_fld_u_0_addr_0 (w_sub00_u_addr),
			.i_fld_u_0_datain_0 (w_sub00_u_datain),
			.o_fld_u_0_dataout_0 (w_sub00_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub00_u_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(9), .WORDS(484) )
		dpram_u_0(
			.clk (clock),
			.ce_0 (w_fld_u_0_ce_0),
			.addr_0 (w_fld_u_0_addr_0),
			.datain_0 (w_fld_u_0_datain_0),
			.dataout_0 (w_fld_u_0_dataout_0),
			.r_w_0 (w_fld_u_0_r_w_0),
			.ce_1 (w_fld_u_0_ce_1),
			.addr_1 (r_fld_u_0_addr_1),
			.datain_1 (r_fld_u_0_datain_1),
			.dataout_1 (w_fld_u_0_dataout_1),
			.r_w_1 (r_fld_u_0_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(9), .WORDS(484) )
		dpram_uu_1(
			.clk (clock),
			.ce_0 (w_fld_uu_1_ce_0),
			.addr_0 (w_fld_uu_1_addr_0),
			.datain_0 (w_fld_uu_1_datain_0),
			.dataout_0 (w_fld_uu_1_dataout_0),
			.r_w_0 (w_fld_uu_1_r_w_0),
			.ce_1 (w_fld_uu_1_ce_1),
			.addr_1 (r_fld_uu_1_addr_1),
			.datain_1 (r_fld_uu_1_datain_1),
			.dataout_1 (w_fld_uu_1_dataout_1),
			.r_w_1 (r_fld_uu_1_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(9), .WORDS(484) )
		dpram_q_2(
			.clk (clock),
			.ce_0 (w_fld_q_2_ce_0),
			.addr_0 (w_fld_q_2_addr_0),
			.datain_0 (w_fld_q_2_datain_0),
			.dataout_0 (w_fld_q_2_dataout_0),
			.r_w_0 (w_fld_q_2_r_w_0),
			.ce_1 (w_fld_q_2_ce_1),
			.addr_1 (r_fld_q_2_addr_1),
			.datain_1 (r_fld_q_2_datain_1),
			.dataout_1 (w_fld_q_2_dataout_1),
			.r_w_1 (r_fld_q_2_r_w_1)
		);

	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h36: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 6'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_phase <= 6'h2;
						end

						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h4;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6) ? 6'h9 : 6'hf);

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'ha;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp9) ? 6'hd : 6'h6);

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h13)) begin
										r_sys_run_phase <= 6'ha;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h10;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp252) ? 6'h14 : 6'h36);

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h10;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h15;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp255) ? 6'h18 : 6'h1a);

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h4f)) begin
										r_sys_run_phase <= 6'h15;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h1b;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp718) ? 6'h1e : 6'h1f);

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h16)) begin
										r_sys_run_phase <= 6'h1b;

									end
								end

							endcase
						end

						6'h1f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_phase <= 6'h21;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h22;

									end
								end

							endcase
						end

						6'h22: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp850) ? 6'h25 : 6'h26);

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h16)) begin
										r_sys_run_phase <= 6'h22;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_phase <= 6'h28;

									end
								end

							endcase
						end

						6'h28: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_phase <= 6'h2a;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h2b;

									end
								end

							endcase
						end

						6'h2b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp981) ? 6'h2e : 6'h30);

									end
								end

							endcase
						end

						6'h2e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h14)) begin
										r_sys_run_phase <= 6'h2b;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h31;

									end
								end

							endcase
						end

						6'h31: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1101) ? 6'h34 : 6'h11);

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h14)) begin
										r_sys_run_phase <= 6'h31;

									end
								end

							endcase
						end

						6'h36: begin
							r_sys_run_phase <= 6'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h13)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h4f)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h16)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h1f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h22: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h16)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h28: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h2b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h2e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h14)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h31: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h14)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 7'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h12)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h4e)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h4f)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h15)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h1f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h22: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h16)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h15)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h28: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub00_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub01_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h2b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h2e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h31: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h14)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						6'h36: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_addr_1 <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp13[8:0] );

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1) || (r_sys_run_step==7'h5) || (r_sys_run_step==7'h9) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h45) || (r_sys_run_step==7'h49) || (r_sys_run_step==7'h4d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp263[8:0] );

									end
									else
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h3e) || (r_sys_run_step==7'h42) || (r_sys_run_step==7'h46) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h4e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp268[8:0] );

									end
									else
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h2b) || (r_sys_run_step==7'h2f) || (r_sys_run_step==7'h33) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h3b) || (r_sys_run_step==7'h3f) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h47) || (r_sys_run_step==7'h4b) || (r_sys_run_step==7'h4f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp273[8:0] );

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h4) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h38) || (r_sys_run_step==7'h3c) || (r_sys_run_step==7'h40) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h48) || (r_sys_run_step==7'h4c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp259[8:0] );

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp837[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp723[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp765[8:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp789[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp807[8:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp783[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp747[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp753[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp831[8:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp795[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp759[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp813[8:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp801[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp777[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp735[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp729[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp819[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp843[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp741[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp825[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp771[8:0] );

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp920[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp938[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp854[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp860[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp950[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp968[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp956[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp902[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp878[8:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp932[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp890[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp908[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp962[8:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp914[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp884[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp866[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp944[8:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp926[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp974[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp872[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp896[8:0] );

									end
								end

							endcase
						end

						6'h2e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp986[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1088[8:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1040[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1010[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1016[8:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1052[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1094[8:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1034[8:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1046[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1070[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1058[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1082[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1022[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp998[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1004[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1028[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1064[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1076[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp992[8:0] );

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1178[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1184[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1124[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1202[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1148[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1112[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1130[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1196[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1142[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1106[8:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1166[8:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1154[8:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1160[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1214[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1136[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1118[8:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1172[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1208[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1190[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp16;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1) || (r_sys_run_step==7'h3) || (r_sys_run_step==7'h5) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'h9) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h2b) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h2f) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h33) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h3b) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h3f) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h45) || (r_sys_run_step==7'h47) || (r_sys_run_step==7'h49) || (r_sys_run_step==7'h4b) || (r_sys_run_step==7'h4d) || (r_sys_run_step==7'h4f)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp266;

									end
									else
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h3e) || (r_sys_run_step==7'h42) || (r_sys_run_step==7'h46) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h4e)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp271;

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h4) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h38) || (r_sys_run_step==7'h3c) || (r_sys_run_step==7'h40) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h48) || (r_sys_run_step==7'h4c)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp261;

									end
								end

							endcase
						end

						6'h2e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h14)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp988;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h14)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp1108;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h4f)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h14)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h14)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h14)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h14)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h36: begin
							r_fld_u_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_uu_1_addr_1 <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_fld_uu_1_addr_1 <= $signed( w_sys_tmp18[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_fld_uu_1_datain_1 <= w_sys_tmp16;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_uu_1_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_fld_uu_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h36: begin
							r_fld_uu_1_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_q_2_addr_1 <= 9'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_q_2_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h36: begin
							r_fld_q_2_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_5 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_5 <= w_sys_tmp8;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_5 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h16)) begin
										r_run_k_5 <= w_sys_tmp848;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_5 <= w_sys_tmp849;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h16)) begin
										r_run_k_5 <= w_sys_tmp979;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_5 <= w_sys_tmp980;

									end
								end

							endcase
						end

						6'h2e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h14)) begin
										r_run_k_5 <= w_sys_tmp1099;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_5 <= w_sys_tmp1100;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h14)) begin
										r_run_k_5 <= w_sys_tmp1219;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_6 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_run_j_6 <= w_sys_tmp23;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_6 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h4) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h38) || (r_sys_run_step==7'h3c) || (r_sys_run_step==7'h40) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h48) || (r_sys_run_step==7'h4c)) begin
										r_run_j_6 <= w_sys_tmp280;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_n_7 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_n_7 <= w_sys_tmp254;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_mx_8 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_my_9 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_nlast_10 <= w_sys_tmp5;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_dx_11 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_dy_12 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_13 <= r_run_j_6;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_run_copy0_j_13 <= w_sys_tmp22;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_14 <= r_run_j_6;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h2b) || (r_sys_run_step==7'h2f) || (r_sys_run_step==7'h33) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h3b) || (r_sys_run_step==7'h3f) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h47) || (r_sys_run_step==7'h4b) || (r_sys_run_step==7'h4f)) begin
										r_run_copy0_j_14 <= w_sys_tmp277;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_15 <= r_run_j_6;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h3e) || (r_sys_run_step==7'h42) || (r_sys_run_step==7'h46) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h4e)) begin
										r_run_copy1_j_15 <= w_sys_tmp278;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy2_j_16 <= r_run_j_6;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1) || (r_sys_run_step==7'h5) || (r_sys_run_step==7'h9) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h45) || (r_sys_run_step==7'h49) || (r_sys_run_step==7'h4d)) begin
										r_run_copy2_j_16 <= w_sys_tmp279;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h26: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp920[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp938[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp854[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp860[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp950[8:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp968[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp956[8:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp902[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp878[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp932[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp890[8:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp908[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp962[8:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp914[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp884[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp866[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp944[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp926[8:0] );

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp974[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp872[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp896[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h16)) begin
										r_sub01_u_datain <= w_sys_tmp856;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h16)) begin
										r_sub01_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h36: begin
							r_sub01_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_q_addr <= 9'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_q_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_q_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_q_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h36: begin
							r_sub01_q_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'hc)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1178[8:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1184[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1124[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1202[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1148[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1112[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1130[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1196[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1142[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1106[8:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1166[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1154[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1160[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1214[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1136[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1118[8:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1172[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1208[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1190[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h12)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h36: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h15)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp837[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp723[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp765[8:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp789[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp807[8:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp783[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp747[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp753[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp831[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp795[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp759[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp813[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp801[8:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp777[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp735[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp729[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp819[8:0] );

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp843[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp741[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp825[8:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp771[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h16)) begin
										r_sub00_u_datain <= w_sys_tmp725;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h16)) begin
										r_sub00_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h1f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h36: begin
							r_sub00_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_q_addr <= 9'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_q_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_q_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_q_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h36: begin
							r_sub00_q_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp986[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1088[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1040[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1010[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1016[8:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1052[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1094[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1034[8:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1046[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1070[8:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1058[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1082[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1022[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp998[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1004[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1028[8:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1064[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1076[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp992[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h12)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h36: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


endmodule
