/*
TimeStamp:	2016/9/9		16:20
*/


module c1(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy,	
	output signed  [31:0] o_run_return	
);

	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [31:0] r_sys_run_return;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 6:0] r_sys_run_phase;
	reg         [ 2:0] r_sys_run_stage;
	reg         [ 4:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 2:0] w_sys_run_stage_p1;
	wire        [ 4:0] w_sys_run_step_p1;
	wire signed [14:0] w_fld_u_0_addr_0;
	wire        [31:0] w_fld_u_0_datain_0;
	wire        [31:0] w_fld_u_0_dataout_0;
	wire               w_fld_u_0_r_w_0;
	wire               w_fld_u_0_ce_0;
	reg  signed [14:0] r_fld_u_0_addr_1;
	reg         [31:0] r_fld_u_0_datain_1;
	wire        [31:0] w_fld_u_0_dataout_1;
	reg                r_fld_u_0_r_w_1;
	wire               w_fld_u_0_ce_1;
	reg  signed [31:0] r_run_k_5;
	reg  signed [31:0] r_run_j_6;
	reg  signed [31:0] r_run_n_7;
	reg  signed [31:0] r_run_mx_8;
	reg  signed [31:0] r_run_my_9;
	reg  signed [31:0] r_run_nlast_10;
	reg         [31:0] r_run_dx_11;
	reg         [31:0] r_run_dy_12;
	reg         [31:0] r_run_r1_13;
	reg         [31:0] r_run_r2_14;
	reg         [31:0] r_run_dt_15;
	reg  signed [31:0] r_run_copy0_j_16;
	reg  signed [31:0] r_run_copy1_j_17;
	reg  signed [31:0] r_run_copy2_j_18;
	reg  signed [31:0] r_run_copy0_j_19;
	reg  signed [31:0] r_run_copy0_j_20;
	reg  signed [31:0] r_run_copy0_j_21;
	reg  signed [31:0] r_run_copy0_j_22;
	reg  signed [31:0] r_run_copy0_j_23;
	reg  signed [31:0] r_run_copy0_j_24;
	reg  signed [31:0] r_run_copy0_j_25;
	reg  signed [31:0] r_run_copy0_j_26;
	reg                r_sub03_run_req;
	wire               w_sub03_run_busy;
	wire signed [14:0] w_sub03_u_addr;
	reg  signed [14:0] r_sub03_u_addr;
	wire        [31:0] w_sub03_u_datain;
	reg         [31:0] r_sub03_u_datain;
	wire        [31:0] w_sub03_u_dataout;
	wire               w_sub03_u_r_w;
	reg                r_sub03_u_r_w;
	wire signed [14:0] w_sub03_result_addr;
	reg  signed [14:0] r_sub03_result_addr;
	wire        [31:0] w_sub03_result_datain;
	reg         [31:0] r_sub03_result_datain;
	wire        [31:0] w_sub03_result_dataout;
	wire               w_sub03_result_r_w;
	reg                r_sub03_result_r_w;
	reg                r_sub02_run_req;
	wire               w_sub02_run_busy;
	wire signed [14:0] w_sub02_u_addr;
	reg  signed [14:0] r_sub02_u_addr;
	wire        [31:0] w_sub02_u_datain;
	reg         [31:0] r_sub02_u_datain;
	wire        [31:0] w_sub02_u_dataout;
	wire               w_sub02_u_r_w;
	reg                r_sub02_u_r_w;
	wire signed [14:0] w_sub02_result_addr;
	reg  signed [14:0] r_sub02_result_addr;
	wire        [31:0] w_sub02_result_datain;
	reg         [31:0] r_sub02_result_datain;
	wire        [31:0] w_sub02_result_dataout;
	wire               w_sub02_result_r_w;
	reg                r_sub02_result_r_w;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [14:0] w_sub01_u_addr;
	reg  signed [14:0] r_sub01_u_addr;
	wire        [31:0] w_sub01_u_datain;
	reg         [31:0] r_sub01_u_datain;
	wire        [31:0] w_sub01_u_dataout;
	wire               w_sub01_u_r_w;
	reg                r_sub01_u_r_w;
	wire signed [14:0] w_sub01_result_addr;
	reg  signed [14:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [14:0] w_sub00_u_addr;
	reg  signed [14:0] r_sub00_u_addr;
	wire        [31:0] w_sub00_u_datain;
	reg         [31:0] r_sub00_u_datain;
	wire        [31:0] w_sub00_u_dataout;
	wire               w_sub00_u_r_w;
	reg                r_sub00_u_r_w;
	wire signed [14:0] w_sub00_result_addr;
	reg  signed [14:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	reg         [31:0] r_sys_tmp0_float;
	wire signed [31:0] w_sys_tmp1;
	wire        [31:0] w_sys_tmp3;
	wire        [31:0] w_sys_tmp4;
	wire        [31:0] w_sys_tmp6;
	wire               w_sys_tmp8;
	wire               w_sys_tmp9;
	wire signed [31:0] w_sys_tmp10;
	wire               w_sys_tmp11;
	wire               w_sys_tmp12;
	wire signed [31:0] w_sys_tmp15;
	wire signed [31:0] w_sys_tmp16;
	wire signed [31:0] w_sys_tmp17;
	wire        [31:0] w_sys_tmp18;
	wire signed [31:0] w_sys_tmp19;
	wire               w_sys_tmp56;
	wire               w_sys_tmp57;
	wire signed [31:0] w_sys_tmp58;
	wire               w_sys_tmp59;
	wire               w_sys_tmp60;
	wire signed [31:0] w_sys_tmp63;
	wire signed [31:0] w_sys_tmp64;
	wire        [31:0] w_sys_tmp65;
	wire signed [31:0] w_sys_tmp67;
	wire signed [31:0] w_sys_tmp68;
	wire        [31:0] w_sys_tmp70;
	wire signed [31:0] w_sys_tmp72;
	wire signed [31:0] w_sys_tmp73;
	wire        [31:0] w_sys_tmp75;
	wire signed [31:0] w_sys_tmp77;
	wire signed [31:0] w_sys_tmp78;
	wire signed [31:0] w_sys_tmp81;
	wire signed [31:0] w_sys_tmp82;
	wire signed [31:0] w_sys_tmp83;
	wire signed [31:0] w_sys_tmp84;
	wire               w_sys_tmp223;
	wire               w_sys_tmp224;
	wire signed [31:0] w_sys_tmp225;
	wire signed [31:0] w_sys_tmp226;
	wire               w_sys_tmp227;
	wire               w_sys_tmp228;
	wire signed [31:0] w_sys_tmp229;
	wire signed [31:0] w_sys_tmp232;
	wire signed [31:0] w_sys_tmp233;
	wire signed [31:0] w_sys_tmp234;
	wire        [31:0] w_sys_tmp235;
	wire signed [31:0] w_sys_tmp236;
	wire signed [31:0] w_sys_tmp237;
	wire signed [31:0] w_sys_tmp239;
	wire signed [31:0] w_sys_tmp240;
	wire signed [31:0] w_sys_tmp301;
	wire               w_sys_tmp302;
	wire               w_sys_tmp303;
	wire signed [31:0] w_sys_tmp304;
	wire signed [31:0] w_sys_tmp307;
	wire signed [31:0] w_sys_tmp308;
	wire signed [31:0] w_sys_tmp309;
	wire        [31:0] w_sys_tmp310;
	wire signed [31:0] w_sys_tmp311;
	wire signed [31:0] w_sys_tmp312;
	wire signed [31:0] w_sys_tmp314;
	wire signed [31:0] w_sys_tmp315;
	wire signed [31:0] w_sys_tmp376;
	wire               w_sys_tmp377;
	wire               w_sys_tmp378;
	wire signed [31:0] w_sys_tmp379;
	wire signed [31:0] w_sys_tmp380;
	wire               w_sys_tmp381;
	wire               w_sys_tmp382;
	wire signed [31:0] w_sys_tmp383;
	wire signed [31:0] w_sys_tmp386;
	wire signed [31:0] w_sys_tmp387;
	wire signed [31:0] w_sys_tmp388;
	wire        [31:0] w_sys_tmp389;
	wire signed [31:0] w_sys_tmp390;
	wire signed [31:0] w_sys_tmp391;
	wire signed [31:0] w_sys_tmp393;
	wire signed [31:0] w_sys_tmp394;
	wire signed [31:0] w_sys_tmp455;
	wire               w_sys_tmp456;
	wire               w_sys_tmp457;
	wire signed [31:0] w_sys_tmp458;
	wire signed [31:0] w_sys_tmp461;
	wire signed [31:0] w_sys_tmp462;
	wire signed [31:0] w_sys_tmp463;
	wire        [31:0] w_sys_tmp464;
	wire signed [31:0] w_sys_tmp465;
	wire signed [31:0] w_sys_tmp466;
	wire signed [31:0] w_sys_tmp468;
	wire signed [31:0] w_sys_tmp469;
	wire signed [31:0] w_sys_tmp530;
	wire               w_sys_tmp531;
	wire               w_sys_tmp532;
	wire signed [31:0] w_sys_tmp533;
	wire signed [31:0] w_sys_tmp534;
	wire signed [31:0] w_sys_tmp535;
	wire               w_sys_tmp536;
	wire               w_sys_tmp537;
	wire signed [31:0] w_sys_tmp538;
	wire signed [31:0] w_sys_tmp541;
	wire signed [31:0] w_sys_tmp542;
	wire signed [31:0] w_sys_tmp543;
	wire        [31:0] w_sys_tmp544;
	wire signed [31:0] w_sys_tmp545;
	wire signed [31:0] w_sys_tmp546;
	wire signed [31:0] w_sys_tmp548;
	wire signed [31:0] w_sys_tmp549;
	wire signed [31:0] w_sys_tmp610;
	wire               w_sys_tmp611;
	wire               w_sys_tmp612;
	wire signed [31:0] w_sys_tmp613;
	wire signed [31:0] w_sys_tmp616;
	wire signed [31:0] w_sys_tmp617;
	wire signed [31:0] w_sys_tmp618;
	wire        [31:0] w_sys_tmp619;
	wire signed [31:0] w_sys_tmp620;
	wire signed [31:0] w_sys_tmp621;
	wire signed [31:0] w_sys_tmp623;
	wire signed [31:0] w_sys_tmp624;
	wire signed [31:0] w_sys_tmp685;
	wire               w_sys_tmp686;
	wire               w_sys_tmp687;
	wire signed [31:0] w_sys_tmp688;
	wire signed [31:0] w_sys_tmp689;
	wire signed [31:0] w_sys_tmp690;
	wire               w_sys_tmp691;
	wire               w_sys_tmp692;
	wire signed [31:0] w_sys_tmp693;
	wire signed [31:0] w_sys_tmp696;
	wire signed [31:0] w_sys_tmp697;
	wire signed [31:0] w_sys_tmp698;
	wire        [31:0] w_sys_tmp699;
	wire signed [31:0] w_sys_tmp700;
	wire signed [31:0] w_sys_tmp701;
	wire signed [31:0] w_sys_tmp703;
	wire signed [31:0] w_sys_tmp704;
	wire signed [31:0] w_sys_tmp765;
	wire               w_sys_tmp766;
	wire               w_sys_tmp767;
	wire signed [31:0] w_sys_tmp768;
	wire signed [31:0] w_sys_tmp771;
	wire signed [31:0] w_sys_tmp772;
	wire signed [31:0] w_sys_tmp773;
	wire        [31:0] w_sys_tmp774;
	wire signed [31:0] w_sys_tmp775;
	wire signed [31:0] w_sys_tmp776;
	wire signed [31:0] w_sys_tmp778;
	wire signed [31:0] w_sys_tmp779;
	wire        [31:0] w_sys_tmp840;
	wire signed [31:0] w_sys_tmp841;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign o_run_return = r_sys_run_return;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 3'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 5'h1);
	assign w_fld_u_0_addr_0 = 15'sh0;
	assign w_fld_u_0_datain_0 = 32'h0;
	assign w_fld_u_0_r_w_0 = 1'h0;
	assign w_fld_u_0_ce_0 = w_sys_ce;
	assign w_fld_u_0_ce_1 = w_sys_ce;
	assign w_sub03_u_addr = ( (|r_sys_processing_methodID) ? r_sub03_u_addr : 15'sh0 ) ;
	assign w_sub03_u_datain = ( (|r_sys_processing_methodID) ? r_sub03_u_datain : 32'h0 ) ;
	assign w_sub03_u_r_w = ( (|r_sys_processing_methodID) ? r_sub03_u_r_w : 1'h0 ) ;
	assign w_sub03_result_addr = ( (|r_sys_processing_methodID) ? r_sub03_result_addr : 15'sh0 ) ;
	assign w_sub03_result_datain = ( (|r_sys_processing_methodID) ? r_sub03_result_datain : 32'h0 ) ;
	assign w_sub03_result_r_w = ( (|r_sys_processing_methodID) ? r_sub03_result_r_w : 1'h0 ) ;
	assign w_sub02_u_addr = ( (|r_sys_processing_methodID) ? r_sub02_u_addr : 15'sh0 ) ;
	assign w_sub02_u_datain = ( (|r_sys_processing_methodID) ? r_sub02_u_datain : 32'h0 ) ;
	assign w_sub02_u_r_w = ( (|r_sys_processing_methodID) ? r_sub02_u_r_w : 1'h0 ) ;
	assign w_sub02_result_addr = ( (|r_sys_processing_methodID) ? r_sub02_result_addr : 15'sh0 ) ;
	assign w_sub02_result_datain = ( (|r_sys_processing_methodID) ? r_sub02_result_datain : 32'h0 ) ;
	assign w_sub02_result_r_w = ( (|r_sys_processing_methodID) ? r_sub02_result_r_w : 1'h0 ) ;
	assign w_sub01_u_addr = ( (|r_sys_processing_methodID) ? r_sub01_u_addr : 15'sh0 ) ;
	assign w_sub01_u_datain = ( (|r_sys_processing_methodID) ? r_sub01_u_datain : 32'h0 ) ;
	assign w_sub01_u_r_w = ( (|r_sys_processing_methodID) ? r_sub01_u_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 15'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub00_u_addr = ( (|r_sys_processing_methodID) ? r_sub00_u_addr : 15'sh0 ) ;
	assign w_sub00_u_datain = ( (|r_sys_processing_methodID) ? r_sub00_u_datain : 32'h0 ) ;
	assign w_sub00_u_r_w = ( (|r_sys_processing_methodID) ? r_sub00_u_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 15'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh00000081;
	assign w_sys_tmp3 = 32'h3a03126f;
	assign w_sys_tmp4 = 32'h3c000000;
	assign w_sys_tmp6 = 32'h4103126f;
	assign w_sys_tmp8 = ( !w_sys_tmp9 );
	assign w_sys_tmp9 = (r_run_my_9 < r_run_k_5);
	assign w_sys_tmp10 = (r_run_k_5 + w_sys_intOne);
	assign w_sys_tmp11 = ( !w_sys_tmp12 );
	assign w_sys_tmp12 = (r_run_mx_8 < r_run_j_6);
	assign w_sys_tmp15 = (w_sys_tmp16 + r_run_k_5);
	assign w_sys_tmp16 = (r_run_j_6 * w_sys_tmp17);
	assign w_sys_tmp17 = 32'sh00000081;
	assign w_sys_tmp18 = 32'h0;
	assign w_sys_tmp19 = (r_run_j_6 + w_sys_intOne);
	assign w_sys_tmp56 = ( !w_sys_tmp57 );
	assign w_sys_tmp57 = (r_run_nlast_10 < r_run_n_7);
	assign w_sys_tmp58 = (r_run_n_7 + w_sys_intOne);
	assign w_sys_tmp59 = ( !w_sys_tmp60 );
	assign w_sys_tmp60 = (r_run_my_9 < r_run_j_6);
	assign w_sys_tmp63 = (w_sys_tmp64 + r_run_j_6);
	assign w_sys_tmp64 = 32'sh00000081;
	assign w_sys_tmp65 = 32'h3f000000;
	assign w_sys_tmp67 = (w_sys_tmp68 + r_run_copy2_j_18);
	assign w_sys_tmp68 = (r_run_mx_8 * w_sys_tmp64);
	assign w_sys_tmp70 = 32'h0;
	assign w_sys_tmp72 = (w_sys_tmp73 + w_sys_intOne);
	assign w_sys_tmp73 = (r_run_copy1_j_17 * w_sys_tmp64);
	assign w_sys_tmp75 = 32'h3f800000;
	assign w_sys_tmp77 = (w_sys_tmp78 + r_run_my_9);
	assign w_sys_tmp78 = (r_run_copy0_j_16 * w_sys_tmp64);
	assign w_sys_tmp81 = (r_run_copy0_j_16 + w_sys_intOne);
	assign w_sys_tmp82 = (r_run_copy1_j_17 + w_sys_intOne);
	assign w_sys_tmp83 = (r_run_copy2_j_18 + w_sys_intOne);
	assign w_sys_tmp84 = (r_run_j_6 + w_sys_intOne);
	assign w_sys_tmp223 = ( !w_sys_tmp224 );
	assign w_sys_tmp224 = (w_sys_tmp225 < r_run_k_5);
	assign w_sys_tmp225 = 32'sh00000041;
	assign w_sys_tmp226 = (r_run_k_5 + w_sys_intOne);
	assign w_sys_tmp227 = ( !w_sys_tmp228 );
	assign w_sys_tmp228 = (w_sys_tmp229 < r_run_j_6);
	assign w_sys_tmp229 = 32'sh00000041;
	assign w_sys_tmp232 = (w_sys_tmp233 + r_run_k_5);
	assign w_sys_tmp233 = (r_run_j_6 * w_sys_tmp234);
	assign w_sys_tmp234 = 32'sh00000081;
	assign w_sys_tmp235 = w_fld_u_0_dataout_1;
	assign w_sys_tmp236 = (w_sys_tmp237 + r_run_k_5);
	assign w_sys_tmp237 = (r_run_copy0_j_19 * w_sys_tmp234);
	assign w_sys_tmp239 = (r_run_copy0_j_19 + w_sys_intOne);
	assign w_sys_tmp240 = (r_run_j_6 + w_sys_intOne);
	assign w_sys_tmp301 = 32'sh00000041;
	assign w_sys_tmp302 = ( !w_sys_tmp303 );
	assign w_sys_tmp303 = (w_sys_tmp304 < r_run_j_6);
	assign w_sys_tmp304 = 32'sh00000081;
	assign w_sys_tmp307 = (w_sys_tmp308 + r_run_k_5);
	assign w_sys_tmp308 = (r_run_j_6 * w_sys_tmp309);
	assign w_sys_tmp309 = 32'sh00000081;
	assign w_sys_tmp310 = w_fld_u_0_dataout_1;
	assign w_sys_tmp311 = (w_sys_tmp312 + r_run_k_5);
	assign w_sys_tmp312 = (r_run_copy0_j_20 * w_sys_tmp309);
	assign w_sys_tmp314 = (r_run_copy0_j_20 + w_sys_intOne);
	assign w_sys_tmp315 = (r_run_j_6 + w_sys_intOne);
	assign w_sys_tmp376 = 32'sh00000040;
	assign w_sys_tmp377 = ( !w_sys_tmp378 );
	assign w_sys_tmp378 = (w_sys_tmp379 < r_run_k_5);
	assign w_sys_tmp379 = 32'sh00000081;
	assign w_sys_tmp380 = (r_run_k_5 + w_sys_intOne);
	assign w_sys_tmp381 = ( !w_sys_tmp382 );
	assign w_sys_tmp382 = (w_sys_tmp383 < r_run_j_6);
	assign w_sys_tmp383 = 32'sh00000041;
	assign w_sys_tmp386 = (w_sys_tmp387 + r_run_k_5);
	assign w_sys_tmp387 = (r_run_j_6 * w_sys_tmp388);
	assign w_sys_tmp388 = 32'sh00000081;
	assign w_sys_tmp389 = w_fld_u_0_dataout_1;
	assign w_sys_tmp390 = (w_sys_tmp391 + r_run_k_5);
	assign w_sys_tmp391 = (r_run_copy0_j_21 * w_sys_tmp388);
	assign w_sys_tmp393 = (r_run_copy0_j_21 + w_sys_intOne);
	assign w_sys_tmp394 = (r_run_j_6 + w_sys_intOne);
	assign w_sys_tmp455 = 32'sh00000041;
	assign w_sys_tmp456 = ( !w_sys_tmp457 );
	assign w_sys_tmp457 = (w_sys_tmp458 < r_run_j_6);
	assign w_sys_tmp458 = 32'sh00000081;
	assign w_sys_tmp461 = (w_sys_tmp462 + r_run_k_5);
	assign w_sys_tmp462 = (r_run_j_6 * w_sys_tmp463);
	assign w_sys_tmp463 = 32'sh00000081;
	assign w_sys_tmp464 = w_fld_u_0_dataout_1;
	assign w_sys_tmp465 = (w_sys_tmp466 + r_run_k_5);
	assign w_sys_tmp466 = (r_run_copy0_j_22 * w_sys_tmp463);
	assign w_sys_tmp468 = (r_run_copy0_j_22 + w_sys_intOne);
	assign w_sys_tmp469 = (r_run_j_6 + w_sys_intOne);
	assign w_sys_tmp530 = 32'sh00000002;
	assign w_sys_tmp531 = ( !w_sys_tmp532 );
	assign w_sys_tmp532 = (w_sys_tmp533 < r_run_k_5);
	assign w_sys_tmp533 = 32'sh00000040;
	assign w_sys_tmp534 = (r_run_k_5 + w_sys_intOne);
	assign w_sys_tmp535 = 32'sh00000002;
	assign w_sys_tmp536 = ( !w_sys_tmp537 );
	assign w_sys_tmp537 = (w_sys_tmp538 < r_run_j_6);
	assign w_sys_tmp538 = 32'sh00000040;
	assign w_sys_tmp541 = (w_sys_tmp542 + r_run_k_5);
	assign w_sys_tmp542 = (r_run_j_6 * w_sys_tmp543);
	assign w_sys_tmp543 = 32'sh00000081;
	assign w_sys_tmp544 = w_sub00_result_dataout;
	assign w_sys_tmp545 = (w_sys_tmp546 + r_run_k_5);
	assign w_sys_tmp546 = (r_run_copy0_j_23 * w_sys_tmp543);
	assign w_sys_tmp548 = (r_run_copy0_j_23 + w_sys_intOne);
	assign w_sys_tmp549 = (r_run_j_6 + w_sys_intOne);
	assign w_sys_tmp610 = 32'sh00000041;
	assign w_sys_tmp611 = ( !w_sys_tmp612 );
	assign w_sys_tmp612 = (w_sys_tmp613 < r_run_j_6);
	assign w_sys_tmp613 = 32'sh00000080;
	assign w_sys_tmp616 = (w_sys_tmp617 + r_run_k_5);
	assign w_sys_tmp617 = (r_run_j_6 * w_sys_tmp618);
	assign w_sys_tmp618 = 32'sh00000081;
	assign w_sys_tmp619 = w_sub01_result_dataout;
	assign w_sys_tmp620 = (w_sys_tmp621 + r_run_k_5);
	assign w_sys_tmp621 = (r_run_copy0_j_24 * w_sys_tmp618);
	assign w_sys_tmp623 = (r_run_copy0_j_24 + w_sys_intOne);
	assign w_sys_tmp624 = (r_run_j_6 + w_sys_intOne);
	assign w_sys_tmp685 = 32'sh00000041;
	assign w_sys_tmp686 = ( !w_sys_tmp687 );
	assign w_sys_tmp687 = (w_sys_tmp688 < r_run_k_5);
	assign w_sys_tmp688 = 32'sh00000080;
	assign w_sys_tmp689 = (r_run_k_5 + w_sys_intOne);
	assign w_sys_tmp690 = 32'sh00000002;
	assign w_sys_tmp691 = ( !w_sys_tmp692 );
	assign w_sys_tmp692 = (w_sys_tmp693 < r_run_j_6);
	assign w_sys_tmp693 = 32'sh00000040;
	assign w_sys_tmp696 = (w_sys_tmp697 + r_run_k_5);
	assign w_sys_tmp697 = (r_run_j_6 * w_sys_tmp698);
	assign w_sys_tmp698 = 32'sh00000081;
	assign w_sys_tmp699 = w_sub02_result_dataout;
	assign w_sys_tmp700 = (w_sys_tmp701 + r_run_k_5);
	assign w_sys_tmp701 = (r_run_copy0_j_25 * w_sys_tmp698);
	assign w_sys_tmp703 = (r_run_copy0_j_25 + w_sys_intOne);
	assign w_sys_tmp704 = (r_run_j_6 + w_sys_intOne);
	assign w_sys_tmp765 = 32'sh00000041;
	assign w_sys_tmp766 = ( !w_sys_tmp767 );
	assign w_sys_tmp767 = (w_sys_tmp768 < r_run_j_6);
	assign w_sys_tmp768 = 32'sh00000080;
	assign w_sys_tmp771 = (w_sys_tmp772 + r_run_k_5);
	assign w_sys_tmp772 = (r_run_j_6 * w_sys_tmp773);
	assign w_sys_tmp773 = 32'sh00000081;
	assign w_sys_tmp774 = w_sub03_result_dataout;
	assign w_sys_tmp775 = (w_sys_tmp776 + r_run_k_5);
	assign w_sys_tmp776 = (r_run_copy0_j_26 * w_sys_tmp773);
	assign w_sys_tmp778 = (r_run_copy0_j_26 + w_sys_intOne);
	assign w_sys_tmp779 = (r_run_j_6 + w_sys_intOne);
	assign w_sys_tmp840 = w_fld_u_0_dataout_1;
	assign w_sys_tmp841 = 32'sh000000dc;


	sub03
		sub03_inst(
			.i_fld_result_1_addr_0 (w_sub03_result_addr),
			.i_fld_result_1_datain_0 (w_sub03_result_datain),
			.o_fld_result_1_dataout_0 (w_sub03_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub03_result_r_w),
			.i_fld_u_0_addr_0 (w_sub03_u_addr),
			.i_fld_u_0_datain_0 (w_sub03_u_datain),
			.o_fld_u_0_dataout_0 (w_sub03_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub03_u_r_w),
			.o_run_busy (w_sub03_run_busy),
			.i_run_req (r_sub03_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub02
		sub02_inst(
			.i_fld_result_1_addr_0 (w_sub02_result_addr),
			.i_fld_result_1_datain_0 (w_sub02_result_datain),
			.o_fld_result_1_dataout_0 (w_sub02_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub02_result_r_w),
			.i_fld_u_0_addr_0 (w_sub02_u_addr),
			.i_fld_u_0_datain_0 (w_sub02_u_datain),
			.o_fld_u_0_dataout_0 (w_sub02_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub02_u_r_w),
			.o_run_busy (w_sub02_run_busy),
			.i_run_req (r_sub02_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub01
		sub01_inst(
			.i_fld_result_1_addr_0 (w_sub01_result_addr),
			.i_fld_result_1_datain_0 (w_sub01_result_datain),
			.o_fld_result_1_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub01_result_r_w),
			.i_fld_u_0_addr_0 (w_sub01_u_addr),
			.i_fld_u_0_datain_0 (w_sub01_u_datain),
			.o_fld_u_0_dataout_0 (w_sub01_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub01_u_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub00
		sub00_inst(
			.i_fld_result_1_addr_0 (w_sub00_result_addr),
			.i_fld_result_1_datain_0 (w_sub00_result_datain),
			.o_fld_result_1_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub00_result_r_w),
			.i_fld_u_0_addr_0 (w_sub00_u_addr),
			.i_fld_u_0_datain_0 (w_sub00_u_datain),
			.o_fld_u_0_dataout_0 (w_sub00_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub00_u_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_u_0(
			.clk (clock),
			.ce_0 (w_fld_u_0_ce_0),
			.addr_0 (w_fld_u_0_addr_0),
			.datain_0 (w_fld_u_0_datain_0),
			.dataout_0 (w_fld_u_0_dataout_0),
			.r_w_0 (w_fld_u_0_r_w_0),
			.ce_1 (w_fld_u_0_ce_1),
			.addr_1 (r_fld_u_0_addr_1),
			.datain_1 (r_fld_u_0_datain_1),
			.dataout_1 (w_fld_u_0_dataout_1),
			.r_w_1 (r_fld_u_0_r_w_1)
		);

	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						7'h63: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_return <= 32'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h60: begin
							r_sys_run_return <= r_sys_tmp0_float;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 7'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h0: begin
							r_sys_run_phase <= 7'h2;
						end

						7'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h4;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h5;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp8) ? 7'h9 : 7'hf);

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h5;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'ha;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp11) ? 7'hd : 7'h6);

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h6)) begin
										r_sys_run_phase <= 7'ha;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h10;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp56) ? 7'h14 : 7'h61);

									end
								end

							endcase
						end

						7'h11: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h10;

									end
								end

							endcase
						end

						7'h14: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h15;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp59) ? 7'h18 : 7'h1a);

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1b)) begin
										r_sys_run_phase <= 7'h15;

									end
								end

							endcase
						end

						7'h1a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h1b;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp223) ? 7'h1f : 7'h2b);

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h1b;

									end
								end

							endcase
						end

						7'h1f: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h20;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp227) ? 7'h23 : 7'h25);

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 7'h20;

									end
								end

							endcase
						end

						7'h25: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h26;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp302) ? 7'h29 : 7'h1c);

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 7'h26;

									end
								end

							endcase
						end

						7'h2b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h2c;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp377) ? 7'h30 : 7'h3b);

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h2c;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h31;

									end
								end

							endcase
						end

						7'h31: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp381) ? 7'h34 : 7'h36);

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 7'h31;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h37;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp456) ? 7'h3a : 7'h2d);

									end
								end

							endcase
						end

						7'h3a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 7'h37;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								3'h3: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_phase <= 7'h3d;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								3'h3: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_phase <= 7'h3f;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h40;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp531) ? 7'h44 : 7'h50);

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h40;

									end
								end

							endcase
						end

						7'h44: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h45;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp536) ? 7'h48 : 7'h4a);

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 7'h45;

									end
								end

							endcase
						end

						7'h4a: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h4b;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp611) ? 7'h4e : 7'h41);

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 7'h4b;

									end
								end

							endcase
						end

						7'h50: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h51;

									end
								end

							endcase
						end

						7'h51: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp686) ? 7'h55 : 7'h11);

									end
								end

							endcase
						end

						7'h52: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h51;

									end
								end

							endcase
						end

						7'h55: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h56;

									end
								end

							endcase
						end

						7'h56: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp691) ? 7'h59 : 7'h5b);

									end
								end

							endcase
						end

						7'h59: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 7'h56;

									end
								end

							endcase
						end

						7'h5b: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h5c;

									end
								end

							endcase
						end

						7'h5c: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp766) ? 7'h5f : 7'h52);

									end
								end

							endcase
						end

						7'h5f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 7'h5c;

									end
								end

							endcase
						end

						7'h60: begin
							r_sys_run_phase <= 7'h63;
						end

						7'h61: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h2)) begin
										r_sys_run_phase <= 7'h60;

									end
								end

							endcase
						end

						7'h63: begin
							r_sys_run_phase <= 7'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 3'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h6)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h11: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h14: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1b)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h1a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h2b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h31: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h3a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h44: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h4a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h50: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h51: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h52: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h55: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h56: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h59: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h5b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h5c: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h5f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h61: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h2)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 5'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h5)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h6)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h11: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h14: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h1a)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h1b)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h1a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h2b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h31: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h3a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub00_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub01_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub02_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub03_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h44: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h4a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h50: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h51: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h52: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h55: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h56: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h59: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h5b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h5c: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h5f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h61: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0) || (r_sys_run_step==5'h1)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h2)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						7'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						7'h63: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp15[14:0] );

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h2) || (r_sys_run_step==5'h6) || (r_sys_run_step==5'ha) || (r_sys_run_step==5'he) || (r_sys_run_step==5'h12) || (r_sys_run_step==5'h16) || (r_sys_run_step==5'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp72[14:0] );

									end
									else
									if((r_sys_run_step==5'h1) || (r_sys_run_step==5'h5) || (r_sys_run_step==5'h9) || (r_sys_run_step==5'hd) || (r_sys_run_step==5'h11) || (r_sys_run_step==5'h15) || (r_sys_run_step==5'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp67[14:0] );

									end
									else
									if((r_sys_run_step==5'h0) || (r_sys_run_step==5'h4) || (r_sys_run_step==5'h8) || (r_sys_run_step==5'hc) || (r_sys_run_step==5'h10) || (r_sys_run_step==5'h14) || (r_sys_run_step==5'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp63[14:0] );

									end
									else
									if((r_sys_run_step==5'h3) || (r_sys_run_step==5'h7) || (r_sys_run_step==5'hb) || (r_sys_run_step==5'hf) || (r_sys_run_step==5'h13) || (r_sys_run_step==5'h17) || (r_sys_run_step==5'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp77[14:0] );

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp236[14:0] );

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp311[14:0] );

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp390[14:0] );

									end
								end

							endcase
						end

						7'h3a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp465[14:0] );

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp541[14:0] );

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp616[14:0] );

									end
								end

							endcase
						end

						7'h59: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp696[14:0] );

									end
								end

							endcase
						end

						7'h5f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp771[14:0] );

									end
								end

							endcase
						end

						7'h61: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp841[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp18;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h2) || (r_sys_run_step==5'h6) || (r_sys_run_step==5'ha) || (r_sys_run_step==5'he) || (r_sys_run_step==5'h12) || (r_sys_run_step==5'h16) || (r_sys_run_step==5'h1a)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp75;

									end
									else
									if((r_sys_run_step==5'h0) || (r_sys_run_step==5'h4) || (r_sys_run_step==5'h8) || (r_sys_run_step==5'hc) || (r_sys_run_step==5'h10) || (r_sys_run_step==5'h14) || (r_sys_run_step==5'h18)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp65;

									end
									else
									if((r_sys_run_step==5'h1) || (r_sys_run_step==5'h3) || (r_sys_run_step==5'h5) || (r_sys_run_step==5'h7) || (r_sys_run_step==5'h9) || (r_sys_run_step==5'hb) || (r_sys_run_step==5'hd) || (r_sys_run_step==5'hf) || (r_sys_run_step==5'h11) || (r_sys_run_step==5'h13) || (r_sys_run_step==5'h15) || (r_sys_run_step==5'h17) || (r_sys_run_step==5'h19) || (r_sys_run_step==5'h1b)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp70;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp544;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp619;

									end
								end

							endcase
						end

						7'h59: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp699;

									end
								end

							endcase
						end

						7'h5f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp774;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h1b)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h59: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h5f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h61: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h63: begin
							r_fld_u_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_5 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_5 <= w_sys_tmp10;

									end
								end

							endcase
						end

						7'h1a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_5 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_5 <= w_sys_tmp226;

									end
								end

							endcase
						end

						7'h2b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_5 <= w_sys_tmp376;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_5 <= w_sys_tmp380;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_5 <= w_sys_tmp530;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_5 <= w_sys_tmp534;

									end
								end

							endcase
						end

						7'h50: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_5 <= w_sys_tmp685;

									end
								end

							endcase
						end

						7'h52: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_5 <= w_sys_tmp689;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_6 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_j_6 <= w_sys_tmp19;

									end
								end

							endcase
						end

						7'h14: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_6 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0) || (r_sys_run_step==5'h4) || (r_sys_run_step==5'h8) || (r_sys_run_step==5'hc) || (r_sys_run_step==5'h10) || (r_sys_run_step==5'h14) || (r_sys_run_step==5'h18)) begin
										r_run_j_6 <= w_sys_tmp84;

									end
								end

							endcase
						end

						7'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_6 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_6 <= w_sys_tmp240;

									end
								end

							endcase
						end

						7'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_6 <= w_sys_tmp301;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_6 <= w_sys_tmp315;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_6 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_6 <= w_sys_tmp394;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_6 <= w_sys_tmp455;

									end
								end

							endcase
						end

						7'h3a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_6 <= w_sys_tmp469;

									end
								end

							endcase
						end

						7'h44: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_6 <= w_sys_tmp535;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_6 <= w_sys_tmp549;

									end
								end

							endcase
						end

						7'h4a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_6 <= w_sys_tmp610;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_6 <= w_sys_tmp624;

									end
								end

							endcase
						end

						7'h55: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_6 <= w_sys_tmp690;

									end
								end

							endcase
						end

						7'h59: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_6 <= w_sys_tmp704;

									end
								end

							endcase
						end

						7'h5b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_6 <= w_sys_tmp765;

									end
								end

							endcase
						end

						7'h5f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_6 <= w_sys_tmp779;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hf: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_n_7 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h11: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_n_7 <= w_sys_tmp58;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_mx_8 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_my_9 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_nlast_10 <= w_sys_intOne;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_dx_11 <= w_sys_tmp4;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_dy_12 <= w_sys_tmp4;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_r1_13 <= w_sys_tmp6;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_r2_14 <= w_sys_tmp6;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_dt_15 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h14: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_16 <= r_run_j_6;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h3) || (r_sys_run_step==5'h7) || (r_sys_run_step==5'hb) || (r_sys_run_step==5'hf) || (r_sys_run_step==5'h13) || (r_sys_run_step==5'h17) || (r_sys_run_step==5'h1b)) begin
										r_run_copy0_j_16 <= w_sys_tmp81;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h14: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy1_j_17 <= r_run_j_6;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h2) || (r_sys_run_step==5'h6) || (r_sys_run_step==5'ha) || (r_sys_run_step==5'he) || (r_sys_run_step==5'h12) || (r_sys_run_step==5'h16) || (r_sys_run_step==5'h1a)) begin
										r_run_copy1_j_17 <= w_sys_tmp82;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h14: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy2_j_18 <= r_run_j_6;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1) || (r_sys_run_step==5'h5) || (r_sys_run_step==5'h9) || (r_sys_run_step==5'hd) || (r_sys_run_step==5'h11) || (r_sys_run_step==5'h15) || (r_sys_run_step==5'h19)) begin
										r_run_copy2_j_18 <= w_sys_tmp83;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h1f: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_19 <= r_run_j_6;

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_19 <= w_sys_tmp239;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h25: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_20 <= r_run_j_6;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_20 <= w_sys_tmp314;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h30: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_21 <= r_run_j_6;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_21 <= w_sys_tmp393;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_22 <= r_run_j_6;

									end
								end

							endcase
						end

						7'h3a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_22 <= w_sys_tmp468;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h44: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_23 <= r_run_j_6;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_23 <= w_sys_tmp548;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4a: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_24 <= r_run_j_6;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_24 <= w_sys_tmp623;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h55: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_25 <= r_run_j_6;

									end
								end

							endcase
						end

						7'h59: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_25 <= w_sys_tmp703;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h5b: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_26 <= r_run_j_6;

									end
								end

							endcase
						end

						7'h5f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_26 <= w_sys_tmp778;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp461[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub03_u_datain <= w_sys_tmp464;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub03_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h63: begin
							r_sub03_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h5f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp775[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h5f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h63: begin
							r_sub03_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp386[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub02_u_datain <= w_sys_tmp389;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub02_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h63: begin
							r_sub02_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h59: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp700[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h59: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h63: begin
							r_sub02_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								3'h2: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h29: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp307[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h29: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub01_u_datain <= w_sys_tmp310;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h29: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub01_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h63: begin
							r_sub01_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp620[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h63: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								3'h3: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h23: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp232[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h23: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub00_u_datain <= w_sys_tmp235;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h23: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub00_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h63: begin
							r_sub00_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h48: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp545[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h63: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h61: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h2)) begin
										r_sys_tmp0_float <= w_sys_tmp840;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
