/*
TimeStamp:	2016/4/8		13:1
*/


module Test(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy	
);

	reg  signed [31:0] r_ip_Multint_multiplicand_0;
	reg  signed [31:0] r_ip_Multint_multiplier_0;
	wire signed [63:0] w_ip_Multint_product_0;
	reg  signed [31:0] r_ip_FixedToFloat_fixed_0;
	wire        [31:0] w_ip_FixedToFloat_floating_0;
	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 5:0] r_sys_run_phase;
	reg         [ 4:0] r_sys_run_stage;
	reg         [ 5:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 4:0] w_sys_run_stage_p1;
	wire        [ 5:0] w_sys_run_step_p1;
	wire signed [ 6:0] w_fld_a_0_addr_0;
	wire        [31:0] w_fld_a_0_datain_0;
	wire        [31:0] w_fld_a_0_dataout_0;
	wire               w_fld_a_0_r_w_0;
	wire               w_fld_a_0_ce_0;
	reg  signed [ 6:0] r_fld_a_0_addr_1;
	reg         [31:0] r_fld_a_0_datain_1;
	wire        [31:0] w_fld_a_0_dataout_1;
	reg                r_fld_a_0_r_w_1;
	wire               w_fld_a_0_ce_1;
	wire signed [ 6:0] w_fld_x_1_addr_0;
	wire        [31:0] w_fld_x_1_datain_0;
	wire        [31:0] w_fld_x_1_dataout_0;
	wire               w_fld_x_1_r_w_0;
	wire               w_fld_x_1_ce_0;
	reg  signed [ 6:0] r_fld_x_1_addr_1;
	reg         [31:0] r_fld_x_1_datain_1;
	wire        [31:0] w_fld_x_1_dataout_1;
	reg                r_fld_x_1_r_w_1;
	wire               w_fld_x_1_ce_1;
	reg  signed [31:0] r_fld_N_2;
	reg  signed [31:0] r_fld_end_3;
	reg         [31:0] r_run_r_24;
	reg  signed [31:0] r_run_j_25;
	reg  signed [31:0] r_run_t_26;
	reg  signed [31:0] r_run_i_27;
	reg  signed [31:0] r_run_i_28;
	reg  signed [31:0] r_run_k_29;
	reg  signed [31:0] r_run_l_30;
	reg  signed [31:0] r_run_j_31;
	reg  signed [31:0] r_run_copy0_i_32;
	reg  signed [31:0] r_run_copy1_i_33;
	reg  signed [31:0] r_run_copy2_i_34;
	reg  signed [31:0] r_run_copy3_i_35;
	reg  signed [31:0] r_run_copy4_i_36;
	reg  signed [31:0] r_run_copy5_i_37;
	reg  signed [31:0] r_run_copy6_i_38;
	reg  signed [31:0] r_run_copy7_i_39;
	reg  signed [31:0] r_run_copy8_i_40;
	reg  signed [31:0] r_run_copy9_i_41;
	reg  signed [31:0] r_run_copy10_i_42;
	reg  signed [31:0] r_run_copy11_i_43;
	reg  signed [31:0] r_run_copy12_i_44;
	reg  signed [31:0] r_run_copy13_i_45;
	reg  signed [31:0] r_run_copy14_i_46;
	reg  signed [31:0] r_run_copy15_i_47;
	reg  signed [31:0] r_run_copy16_i_48;
	reg  signed [31:0] r_run_copy17_i_49;
	reg  signed [31:0] r_run_copy18_i_50;
	reg  signed [31:0] r_run_copy19_i_51;
	reg  signed [31:0] r_run_copy20_i_52;
	reg  signed [31:0] r_run_copy21_i_53;
	reg  signed [31:0] r_run_copy22_i_54;
	reg  signed [31:0] r_run_copy23_i_55;
	reg  signed [31:0] r_run_copy24_i_56;
	reg  signed [31:0] r_run_copy25_i_57;
	reg  signed [31:0] r_run_copy26_i_58;
	reg  signed [31:0] r_run_copy27_i_59;
	reg  signed [31:0] r_run_copy28_i_60;
	reg  signed [31:0] r_run_copy29_i_61;
	reg  signed [31:0] r_run_copy30_i_62;
	reg  signed [31:0] r_run_copy31_i_63;
	reg  signed [31:0] r_run_copy32_i_64;
	reg  signed [31:0] r_run_copy33_i_65;
	reg  signed [31:0] r_run_copy34_i_66;
	reg  signed [31:0] r_run_copy35_i_67;
	reg  signed [31:0] r_run_copy36_i_68;
	reg  signed [31:0] r_run_copy37_i_69;
	reg  signed [31:0] r_run_copy38_i_70;
	reg  signed [31:0] r_run_copy0_i_71;
	reg  signed [31:0] r_run_copy1_i_72;
	reg  signed [31:0] r_run_copy2_i_73;
	reg  signed [31:0] r_run_copy3_i_74;
	reg  signed [31:0] r_run_copy4_i_75;
	reg  signed [31:0] r_run_copy5_i_76;
	reg  signed [31:0] r_run_copy6_i_77;
	reg  signed [31:0] r_run_copy7_i_78;
	reg  signed [31:0] r_run_copy8_i_79;
	reg  signed [31:0] r_run_copy9_i_80;
	reg  signed [31:0] r_run_copy10_i_81;
	reg  signed [31:0] r_run_copy11_i_82;
	reg  signed [31:0] r_run_copy12_i_83;
	reg  signed [31:0] r_run_copy13_i_84;
	reg  signed [31:0] r_run_copy14_i_85;
	reg  signed [31:0] r_run_copy15_i_86;
	reg  signed [31:0] r_run_copy16_i_87;
	reg  signed [31:0] r_run_copy17_i_88;
	reg  signed [31:0] r_run_copy18_i_89;
	reg  signed [31:0] r_run_copy19_i_90;
	reg                r_sub19_run_req;
	wire               w_sub19_run_busy;
	wire signed [ 2:0] w_sub19_arrayA_addr;
	reg  signed [ 2:0] r_sub19_arrayA_addr;
	wire        [31:0] w_sub19_arrayA_datain;
	reg         [31:0] r_sub19_arrayA_datain;
	wire        [31:0] w_sub19_arrayA_dataout;
	wire               w_sub19_arrayA_r_w;
	reg                r_sub19_arrayA_r_w;
	wire signed [ 2:0] w_sub19_arrayX_addr;
	reg  signed [ 2:0] r_sub19_arrayX_addr;
	wire        [31:0] w_sub19_arrayX_datain;
	reg         [31:0] r_sub19_arrayX_datain;
	wire        [31:0] w_sub19_arrayX_dataout;
	wire               w_sub19_arrayX_r_w;
	reg                r_sub19_arrayX_r_w;
	reg                r_sub09_run_req;
	wire               w_sub09_run_busy;
	wire signed [ 2:0] w_sub09_arrayA_addr;
	reg  signed [ 2:0] r_sub09_arrayA_addr;
	wire        [31:0] w_sub09_arrayA_datain;
	reg         [31:0] r_sub09_arrayA_datain;
	wire        [31:0] w_sub09_arrayA_dataout;
	wire               w_sub09_arrayA_r_w;
	reg                r_sub09_arrayA_r_w;
	wire signed [ 2:0] w_sub09_arrayX_addr;
	reg  signed [ 2:0] r_sub09_arrayX_addr;
	wire        [31:0] w_sub09_arrayX_datain;
	reg         [31:0] r_sub09_arrayX_datain;
	wire        [31:0] w_sub09_arrayX_dataout;
	wire               w_sub09_arrayX_r_w;
	reg                r_sub09_arrayX_r_w;
	reg                r_sub08_run_req;
	wire               w_sub08_run_busy;
	wire signed [ 2:0] w_sub08_arrayA_addr;
	reg  signed [ 2:0] r_sub08_arrayA_addr;
	wire        [31:0] w_sub08_arrayA_datain;
	reg         [31:0] r_sub08_arrayA_datain;
	wire        [31:0] w_sub08_arrayA_dataout;
	wire               w_sub08_arrayA_r_w;
	reg                r_sub08_arrayA_r_w;
	wire signed [ 2:0] w_sub08_arrayX_addr;
	reg  signed [ 2:0] r_sub08_arrayX_addr;
	wire        [31:0] w_sub08_arrayX_datain;
	reg         [31:0] r_sub08_arrayX_datain;
	wire        [31:0] w_sub08_arrayX_dataout;
	wire               w_sub08_arrayX_r_w;
	reg                r_sub08_arrayX_r_w;
	reg                r_sub12_run_req;
	wire               w_sub12_run_busy;
	wire signed [ 2:0] w_sub12_arrayA_addr;
	reg  signed [ 2:0] r_sub12_arrayA_addr;
	wire        [31:0] w_sub12_arrayA_datain;
	reg         [31:0] r_sub12_arrayA_datain;
	wire        [31:0] w_sub12_arrayA_dataout;
	wire               w_sub12_arrayA_r_w;
	reg                r_sub12_arrayA_r_w;
	wire signed [ 2:0] w_sub12_arrayX_addr;
	reg  signed [ 2:0] r_sub12_arrayX_addr;
	wire        [31:0] w_sub12_arrayX_datain;
	reg         [31:0] r_sub12_arrayX_datain;
	wire        [31:0] w_sub12_arrayX_dataout;
	wire               w_sub12_arrayX_r_w;
	reg                r_sub12_arrayX_r_w;
	reg                r_sub03_run_req;
	wire               w_sub03_run_busy;
	wire signed [ 2:0] w_sub03_arrayA_addr;
	reg  signed [ 2:0] r_sub03_arrayA_addr;
	wire        [31:0] w_sub03_arrayA_datain;
	reg         [31:0] r_sub03_arrayA_datain;
	wire        [31:0] w_sub03_arrayA_dataout;
	wire               w_sub03_arrayA_r_w;
	reg                r_sub03_arrayA_r_w;
	wire signed [ 2:0] w_sub03_arrayX_addr;
	reg  signed [ 2:0] r_sub03_arrayX_addr;
	wire        [31:0] w_sub03_arrayX_datain;
	reg         [31:0] r_sub03_arrayX_datain;
	wire        [31:0] w_sub03_arrayX_dataout;
	wire               w_sub03_arrayX_r_w;
	reg                r_sub03_arrayX_r_w;
	reg                r_sub02_run_req;
	wire               w_sub02_run_busy;
	wire signed [ 2:0] w_sub02_arrayA_addr;
	reg  signed [ 2:0] r_sub02_arrayA_addr;
	wire        [31:0] w_sub02_arrayA_datain;
	reg         [31:0] r_sub02_arrayA_datain;
	wire        [31:0] w_sub02_arrayA_dataout;
	wire               w_sub02_arrayA_r_w;
	reg                r_sub02_arrayA_r_w;
	wire signed [ 2:0] w_sub02_arrayX_addr;
	reg  signed [ 2:0] r_sub02_arrayX_addr;
	wire        [31:0] w_sub02_arrayX_datain;
	reg         [31:0] r_sub02_arrayX_datain;
	wire        [31:0] w_sub02_arrayX_dataout;
	wire               w_sub02_arrayX_r_w;
	reg                r_sub02_arrayX_r_w;
	reg                r_sub11_run_req;
	wire               w_sub11_run_busy;
	wire signed [ 2:0] w_sub11_arrayA_addr;
	reg  signed [ 2:0] r_sub11_arrayA_addr;
	wire        [31:0] w_sub11_arrayA_datain;
	reg         [31:0] r_sub11_arrayA_datain;
	wire        [31:0] w_sub11_arrayA_dataout;
	wire               w_sub11_arrayA_r_w;
	reg                r_sub11_arrayA_r_w;
	wire signed [ 2:0] w_sub11_arrayX_addr;
	reg  signed [ 2:0] r_sub11_arrayX_addr;
	wire        [31:0] w_sub11_arrayX_datain;
	reg         [31:0] r_sub11_arrayX_datain;
	wire        [31:0] w_sub11_arrayX_dataout;
	wire               w_sub11_arrayX_r_w;
	reg                r_sub11_arrayX_r_w;
	reg                r_sub14_run_req;
	wire               w_sub14_run_busy;
	wire signed [ 2:0] w_sub14_arrayA_addr;
	reg  signed [ 2:0] r_sub14_arrayA_addr;
	wire        [31:0] w_sub14_arrayA_datain;
	reg         [31:0] r_sub14_arrayA_datain;
	wire        [31:0] w_sub14_arrayA_dataout;
	wire               w_sub14_arrayA_r_w;
	reg                r_sub14_arrayA_r_w;
	wire signed [ 2:0] w_sub14_arrayX_addr;
	reg  signed [ 2:0] r_sub14_arrayX_addr;
	wire        [31:0] w_sub14_arrayX_datain;
	reg         [31:0] r_sub14_arrayX_datain;
	wire        [31:0] w_sub14_arrayX_dataout;
	wire               w_sub14_arrayX_r_w;
	reg                r_sub14_arrayX_r_w;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [ 2:0] w_sub01_arrayA_addr;
	reg  signed [ 2:0] r_sub01_arrayA_addr;
	wire        [31:0] w_sub01_arrayA_datain;
	reg         [31:0] r_sub01_arrayA_datain;
	wire        [31:0] w_sub01_arrayA_dataout;
	wire               w_sub01_arrayA_r_w;
	reg                r_sub01_arrayA_r_w;
	wire signed [ 2:0] w_sub01_arrayX_addr;
	reg  signed [ 2:0] r_sub01_arrayX_addr;
	wire        [31:0] w_sub01_arrayX_datain;
	reg         [31:0] r_sub01_arrayX_datain;
	wire        [31:0] w_sub01_arrayX_dataout;
	wire               w_sub01_arrayX_r_w;
	reg                r_sub01_arrayX_r_w;
	reg                r_sub13_run_req;
	wire               w_sub13_run_busy;
	wire signed [ 2:0] w_sub13_arrayA_addr;
	reg  signed [ 2:0] r_sub13_arrayA_addr;
	wire        [31:0] w_sub13_arrayA_datain;
	reg         [31:0] r_sub13_arrayA_datain;
	wire        [31:0] w_sub13_arrayA_dataout;
	wire               w_sub13_arrayA_r_w;
	reg                r_sub13_arrayA_r_w;
	wire signed [ 2:0] w_sub13_arrayX_addr;
	reg  signed [ 2:0] r_sub13_arrayX_addr;
	wire        [31:0] w_sub13_arrayX_datain;
	reg         [31:0] r_sub13_arrayX_datain;
	wire        [31:0] w_sub13_arrayX_dataout;
	wire               w_sub13_arrayX_r_w;
	reg                r_sub13_arrayX_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [ 2:0] w_sub00_arrayA_addr;
	reg  signed [ 2:0] r_sub00_arrayA_addr;
	wire        [31:0] w_sub00_arrayA_datain;
	reg         [31:0] r_sub00_arrayA_datain;
	wire        [31:0] w_sub00_arrayA_dataout;
	wire               w_sub00_arrayA_r_w;
	reg                r_sub00_arrayA_r_w;
	wire signed [ 2:0] w_sub00_arrayX_addr;
	reg  signed [ 2:0] r_sub00_arrayX_addr;
	wire        [31:0] w_sub00_arrayX_datain;
	reg         [31:0] r_sub00_arrayX_datain;
	wire        [31:0] w_sub00_arrayX_dataout;
	wire               w_sub00_arrayX_r_w;
	reg                r_sub00_arrayX_r_w;
	reg                r_sub07_run_req;
	wire               w_sub07_run_busy;
	wire signed [ 2:0] w_sub07_arrayA_addr;
	reg  signed [ 2:0] r_sub07_arrayA_addr;
	wire        [31:0] w_sub07_arrayA_datain;
	reg         [31:0] r_sub07_arrayA_datain;
	wire        [31:0] w_sub07_arrayA_dataout;
	wire               w_sub07_arrayA_r_w;
	reg                r_sub07_arrayA_r_w;
	wire signed [ 2:0] w_sub07_arrayX_addr;
	reg  signed [ 2:0] r_sub07_arrayX_addr;
	wire        [31:0] w_sub07_arrayX_datain;
	reg         [31:0] r_sub07_arrayX_datain;
	wire        [31:0] w_sub07_arrayX_dataout;
	wire               w_sub07_arrayX_r_w;
	reg                r_sub07_arrayX_r_w;
	reg                r_sub16_run_req;
	wire               w_sub16_run_busy;
	wire signed [ 2:0] w_sub16_arrayA_addr;
	reg  signed [ 2:0] r_sub16_arrayA_addr;
	wire        [31:0] w_sub16_arrayA_datain;
	reg         [31:0] r_sub16_arrayA_datain;
	wire        [31:0] w_sub16_arrayA_dataout;
	wire               w_sub16_arrayA_r_w;
	reg                r_sub16_arrayA_r_w;
	wire signed [ 2:0] w_sub16_arrayX_addr;
	reg  signed [ 2:0] r_sub16_arrayX_addr;
	wire        [31:0] w_sub16_arrayX_datain;
	reg         [31:0] r_sub16_arrayX_datain;
	wire        [31:0] w_sub16_arrayX_dataout;
	wire               w_sub16_arrayX_r_w;
	reg                r_sub16_arrayX_r_w;
	reg                r_sub06_run_req;
	wire               w_sub06_run_busy;
	wire signed [ 2:0] w_sub06_arrayA_addr;
	reg  signed [ 2:0] r_sub06_arrayA_addr;
	wire        [31:0] w_sub06_arrayA_datain;
	reg         [31:0] r_sub06_arrayA_datain;
	wire        [31:0] w_sub06_arrayA_dataout;
	wire               w_sub06_arrayA_r_w;
	reg                r_sub06_arrayA_r_w;
	wire signed [ 2:0] w_sub06_arrayX_addr;
	reg  signed [ 2:0] r_sub06_arrayX_addr;
	wire        [31:0] w_sub06_arrayX_datain;
	reg         [31:0] r_sub06_arrayX_datain;
	wire        [31:0] w_sub06_arrayX_dataout;
	wire               w_sub06_arrayX_r_w;
	reg                r_sub06_arrayX_r_w;
	reg                r_sub15_run_req;
	wire               w_sub15_run_busy;
	wire signed [ 2:0] w_sub15_arrayA_addr;
	reg  signed [ 2:0] r_sub15_arrayA_addr;
	wire        [31:0] w_sub15_arrayA_datain;
	reg         [31:0] r_sub15_arrayA_datain;
	wire        [31:0] w_sub15_arrayA_dataout;
	wire               w_sub15_arrayA_r_w;
	reg                r_sub15_arrayA_r_w;
	wire signed [ 2:0] w_sub15_arrayX_addr;
	reg  signed [ 2:0] r_sub15_arrayX_addr;
	wire        [31:0] w_sub15_arrayX_datain;
	reg         [31:0] r_sub15_arrayX_datain;
	wire        [31:0] w_sub15_arrayX_dataout;
	wire               w_sub15_arrayX_r_w;
	reg                r_sub15_arrayX_r_w;
	reg                r_sub05_run_req;
	wire               w_sub05_run_busy;
	wire signed [ 2:0] w_sub05_arrayA_addr;
	reg  signed [ 2:0] r_sub05_arrayA_addr;
	wire        [31:0] w_sub05_arrayA_datain;
	reg         [31:0] r_sub05_arrayA_datain;
	wire        [31:0] w_sub05_arrayA_dataout;
	wire               w_sub05_arrayA_r_w;
	reg                r_sub05_arrayA_r_w;
	wire signed [ 2:0] w_sub05_arrayX_addr;
	reg  signed [ 2:0] r_sub05_arrayX_addr;
	wire        [31:0] w_sub05_arrayX_datain;
	reg         [31:0] r_sub05_arrayX_datain;
	wire        [31:0] w_sub05_arrayX_dataout;
	wire               w_sub05_arrayX_r_w;
	reg                r_sub05_arrayX_r_w;
	reg                r_sub18_run_req;
	wire               w_sub18_run_busy;
	wire signed [ 2:0] w_sub18_arrayA_addr;
	reg  signed [ 2:0] r_sub18_arrayA_addr;
	wire        [31:0] w_sub18_arrayA_datain;
	reg         [31:0] r_sub18_arrayA_datain;
	wire        [31:0] w_sub18_arrayA_dataout;
	wire               w_sub18_arrayA_r_w;
	reg                r_sub18_arrayA_r_w;
	wire signed [ 2:0] w_sub18_arrayX_addr;
	reg  signed [ 2:0] r_sub18_arrayX_addr;
	wire        [31:0] w_sub18_arrayX_datain;
	reg         [31:0] r_sub18_arrayX_datain;
	wire        [31:0] w_sub18_arrayX_dataout;
	wire               w_sub18_arrayX_r_w;
	reg                r_sub18_arrayX_r_w;
	reg                r_sub04_run_req;
	wire               w_sub04_run_busy;
	wire signed [ 2:0] w_sub04_arrayA_addr;
	reg  signed [ 2:0] r_sub04_arrayA_addr;
	wire        [31:0] w_sub04_arrayA_datain;
	reg         [31:0] r_sub04_arrayA_datain;
	wire        [31:0] w_sub04_arrayA_dataout;
	wire               w_sub04_arrayA_r_w;
	reg                r_sub04_arrayA_r_w;
	wire signed [ 2:0] w_sub04_arrayX_addr;
	reg  signed [ 2:0] r_sub04_arrayX_addr;
	wire        [31:0] w_sub04_arrayX_datain;
	reg         [31:0] r_sub04_arrayX_datain;
	wire        [31:0] w_sub04_arrayX_dataout;
	wire               w_sub04_arrayX_r_w;
	reg                r_sub04_arrayX_r_w;
	reg                r_sub17_run_req;
	wire               w_sub17_run_busy;
	wire signed [ 2:0] w_sub17_arrayA_addr;
	reg  signed [ 2:0] r_sub17_arrayA_addr;
	wire        [31:0] w_sub17_arrayA_datain;
	reg         [31:0] r_sub17_arrayA_datain;
	wire        [31:0] w_sub17_arrayA_dataout;
	wire               w_sub17_arrayA_r_w;
	reg                r_sub17_arrayA_r_w;
	wire signed [ 2:0] w_sub17_arrayX_addr;
	reg  signed [ 2:0] r_sub17_arrayX_addr;
	wire        [31:0] w_sub17_arrayX_datain;
	reg         [31:0] r_sub17_arrayX_datain;
	wire        [31:0] w_sub17_arrayX_dataout;
	wire               w_sub17_arrayX_r_w;
	reg                r_sub17_arrayX_r_w;
	reg                r_sub10_run_req;
	wire               w_sub10_run_busy;
	wire signed [ 2:0] w_sub10_arrayA_addr;
	reg  signed [ 2:0] r_sub10_arrayA_addr;
	wire        [31:0] w_sub10_arrayA_datain;
	reg         [31:0] r_sub10_arrayA_datain;
	wire        [31:0] w_sub10_arrayA_dataout;
	wire               w_sub10_arrayA_r_w;
	reg                r_sub10_arrayA_r_w;
	wire signed [ 2:0] w_sub10_arrayX_addr;
	reg  signed [ 2:0] r_sub10_arrayX_addr;
	wire        [31:0] w_sub10_arrayX_datain;
	reg         [31:0] r_sub10_arrayX_datain;
	wire        [31:0] w_sub10_arrayX_dataout;
	wire               w_sub10_arrayX_r_w;
	reg                r_sub10_arrayX_r_w;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg         [31:0] r_sys_tmp4_float;
	reg         [31:0] r_sys_tmp5_float;
	reg         [31:0] r_sys_tmp6_float;
	reg         [31:0] r_sys_tmp7_float;
	reg         [31:0] r_sys_tmp8_float;
	reg         [31:0] r_sys_tmp9_float;
	reg         [31:0] r_sys_tmp10_float;
	reg         [31:0] r_sys_tmp11_float;
	reg         [31:0] r_sys_tmp12_float;
	reg         [31:0] r_sys_tmp13_float;
	reg         [31:0] r_sys_tmp14_float;
	reg         [31:0] r_sys_tmp15_float;
	reg         [31:0] r_sys_tmp16_float;
	reg         [31:0] r_sys_tmp17_float;
	reg         [31:0] r_sys_tmp18_float;
	reg         [31:0] r_sys_tmp19_float;
	reg         [31:0] r_sys_tmp20_float;
	reg         [31:0] r_sys_tmp21_float;
	reg         [31:0] r_sys_tmp22_float;
	reg         [31:0] r_sys_tmp23_float;
	reg         [31:0] r_sys_tmp24_float;
	reg         [31:0] r_sys_tmp25_float;
	reg         [31:0] r_sys_tmp26_float;
	reg         [31:0] r_sys_tmp27_float;
	reg         [31:0] r_sys_tmp28_float;
	reg         [31:0] r_sys_tmp29_float;
	reg         [31:0] r_sys_tmp30_float;
	reg         [31:0] r_sys_tmp31_float;
	reg         [31:0] r_sys_tmp32_float;
	reg         [31:0] r_sys_tmp33_float;
	reg         [31:0] r_sys_tmp34_float;
	reg         [31:0] r_sys_tmp35_float;
	reg         [31:0] r_sys_tmp36_float;
	reg         [31:0] r_sys_tmp37_float;
	reg         [31:0] r_sys_tmp38_float;
	reg         [31:0] r_sys_tmp39_float;
	reg         [31:0] r_sys_tmp40_float;
	reg         [31:0] r_sys_tmp41_float;
	reg         [31:0] r_sys_tmp42_float;
	reg         [31:0] r_sys_tmp43_float;
	reg         [31:0] r_sys_tmp44_float;
	reg         [31:0] r_sys_tmp45_float;
	reg         [31:0] r_sys_tmp46_float;
	reg         [31:0] r_sys_tmp47_float;
	reg         [31:0] r_sys_tmp48_float;
	reg         [31:0] r_sys_tmp49_float;
	reg         [31:0] r_sys_tmp50_float;
	reg         [31:0] r_sys_tmp51_float;
	reg         [31:0] r_sys_tmp52_float;
	reg         [31:0] r_sys_tmp53_float;
	reg         [31:0] r_sys_tmp54_float;
	reg         [31:0] r_sys_tmp55_float;
	reg         [31:0] r_sys_tmp56_float;
	wire        [31:0] w_sys_tmp1;
	wire               w_sys_tmp2;
	wire        [31:0] w_sys_tmp5;
	wire signed [31:0] w_sys_tmp6;
	wire signed [31:0] w_sys_tmp7;
	wire               w_sys_tmp8;
	wire signed [31:0] w_sys_tmp9;
	wire               w_sys_tmp10;
	wire signed [31:0] w_sys_tmp11;
	wire        [31:0] w_sys_tmp14;
	wire signed [31:0] w_sys_tmp17;
	wire signed [31:0] w_sys_tmp18;
	wire signed [31:0] w_sys_tmp21;
	wire signed [31:0] w_sys_tmp22;
	wire signed [31:0] w_sys_tmp25;
	wire signed [31:0] w_sys_tmp26;
	wire signed [31:0] w_sys_tmp29;
	wire signed [31:0] w_sys_tmp30;
	wire signed [31:0] w_sys_tmp33;
	wire signed [31:0] w_sys_tmp34;
	wire signed [31:0] w_sys_tmp37;
	wire signed [31:0] w_sys_tmp38;
	wire signed [31:0] w_sys_tmp41;
	wire signed [31:0] w_sys_tmp42;
	wire signed [31:0] w_sys_tmp45;
	wire signed [31:0] w_sys_tmp46;
	wire signed [31:0] w_sys_tmp49;
	wire signed [31:0] w_sys_tmp50;
	wire signed [31:0] w_sys_tmp53;
	wire signed [31:0] w_sys_tmp54;
	wire signed [31:0] w_sys_tmp57;
	wire signed [31:0] w_sys_tmp58;
	wire signed [31:0] w_sys_tmp61;
	wire signed [31:0] w_sys_tmp62;
	wire signed [31:0] w_sys_tmp65;
	wire signed [31:0] w_sys_tmp66;
	wire signed [31:0] w_sys_tmp69;
	wire signed [31:0] w_sys_tmp70;
	wire signed [31:0] w_sys_tmp73;
	wire signed [31:0] w_sys_tmp74;
	wire signed [31:0] w_sys_tmp77;
	wire signed [31:0] w_sys_tmp78;
	wire signed [31:0] w_sys_tmp81;
	wire signed [31:0] w_sys_tmp82;
	wire signed [31:0] w_sys_tmp85;
	wire signed [31:0] w_sys_tmp86;
	wire signed [31:0] w_sys_tmp89;
	wire signed [31:0] w_sys_tmp90;
	wire signed [31:0] w_sys_tmp91;
	wire signed [31:0] w_sys_tmp92;
	wire signed [31:0] w_sys_tmp93;
	wire signed [31:0] w_sys_tmp94;
	wire signed [31:0] w_sys_tmp95;
	wire signed [31:0] w_sys_tmp96;
	wire signed [31:0] w_sys_tmp97;
	wire signed [31:0] w_sys_tmp98;
	wire signed [31:0] w_sys_tmp99;
	wire signed [31:0] w_sys_tmp100;
	wire signed [31:0] w_sys_tmp101;
	wire signed [31:0] w_sys_tmp102;
	wire signed [31:0] w_sys_tmp103;
	wire signed [31:0] w_sys_tmp104;
	wire signed [31:0] w_sys_tmp105;
	wire signed [31:0] w_sys_tmp106;
	wire signed [31:0] w_sys_tmp107;
	wire signed [31:0] w_sys_tmp108;
	wire signed [31:0] w_sys_tmp109;
	wire signed [31:0] w_sys_tmp110;
	wire signed [31:0] w_sys_tmp111;
	wire signed [31:0] w_sys_tmp112;
	wire signed [31:0] w_sys_tmp113;
	wire signed [31:0] w_sys_tmp114;
	wire signed [31:0] w_sys_tmp115;
	wire signed [31:0] w_sys_tmp116;
	wire signed [31:0] w_sys_tmp117;
	wire signed [31:0] w_sys_tmp118;
	wire signed [31:0] w_sys_tmp119;
	wire signed [31:0] w_sys_tmp120;
	wire signed [31:0] w_sys_tmp121;
	wire signed [31:0] w_sys_tmp122;
	wire signed [31:0] w_sys_tmp123;
	wire signed [31:0] w_sys_tmp124;
	wire signed [31:0] w_sys_tmp125;
	wire signed [31:0] w_sys_tmp126;
	wire signed [31:0] w_sys_tmp127;
	wire signed [31:0] w_sys_tmp128;
	wire signed [31:0] w_sys_tmp129;
	wire signed [31:0] w_sys_tmp130;
	wire signed [31:0] w_sys_tmp367;
	wire               w_sys_tmp368;
	wire signed [31:0] w_sys_tmp369;
	wire        [31:0] w_sys_tmp374;
	wire signed [31:0] w_sys_tmp376;
	wire signed [31:0] w_sys_tmp377;
	wire signed [31:0] w_sys_tmp379;
	wire signed [31:0] w_sys_tmp380;
	wire signed [31:0] w_sys_tmp382;
	wire signed [31:0] w_sys_tmp383;
	wire signed [31:0] w_sys_tmp385;
	wire signed [31:0] w_sys_tmp386;
	wire signed [31:0] w_sys_tmp388;
	wire signed [31:0] w_sys_tmp389;
	wire signed [31:0] w_sys_tmp391;
	wire signed [31:0] w_sys_tmp392;
	wire signed [31:0] w_sys_tmp394;
	wire signed [31:0] w_sys_tmp395;
	wire signed [31:0] w_sys_tmp397;
	wire signed [31:0] w_sys_tmp398;
	wire signed [31:0] w_sys_tmp400;
	wire signed [31:0] w_sys_tmp401;
	wire signed [31:0] w_sys_tmp403;
	wire signed [31:0] w_sys_tmp404;
	wire signed [31:0] w_sys_tmp406;
	wire signed [31:0] w_sys_tmp407;
	wire signed [31:0] w_sys_tmp409;
	wire signed [31:0] w_sys_tmp410;
	wire signed [31:0] w_sys_tmp412;
	wire signed [31:0] w_sys_tmp413;
	wire signed [31:0] w_sys_tmp415;
	wire signed [31:0] w_sys_tmp416;
	wire signed [31:0] w_sys_tmp418;
	wire signed [31:0] w_sys_tmp419;
	wire signed [31:0] w_sys_tmp421;
	wire signed [31:0] w_sys_tmp422;
	wire signed [31:0] w_sys_tmp424;
	wire signed [31:0] w_sys_tmp425;
	wire signed [31:0] w_sys_tmp427;
	wire signed [31:0] w_sys_tmp428;
	wire signed [31:0] w_sys_tmp430;
	wire signed [31:0] w_sys_tmp431;
	wire signed [31:0] w_sys_tmp432;
	wire signed [31:0] w_sys_tmp433;
	wire signed [31:0] w_sys_tmp434;
	wire signed [31:0] w_sys_tmp435;
	wire signed [31:0] w_sys_tmp436;
	wire signed [31:0] w_sys_tmp437;
	wire signed [31:0] w_sys_tmp438;
	wire signed [31:0] w_sys_tmp439;
	wire signed [31:0] w_sys_tmp440;
	wire signed [31:0] w_sys_tmp441;
	wire signed [31:0] w_sys_tmp442;
	wire signed [31:0] w_sys_tmp443;
	wire signed [31:0] w_sys_tmp444;
	wire signed [31:0] w_sys_tmp445;
	wire signed [31:0] w_sys_tmp446;
	wire signed [31:0] w_sys_tmp447;
	wire signed [31:0] w_sys_tmp448;
	wire signed [31:0] w_sys_tmp449;
	wire signed [31:0] w_sys_tmp450;
	wire signed [31:0] w_sys_tmp451;
	wire signed [31:0] w_sys_tmp452;
	wire signed [31:0] w_sys_tmp453;
	wire signed [31:0] w_sys_tmp454;
	wire               w_sys_tmp617;
	wire        [31:0] w_sys_tmp620;
	wire signed [31:0] w_sys_tmp621;
	wire signed [31:0] w_sys_tmp622;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 5'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 6'h1);
	assign w_fld_a_0_addr_0 = 7'sh0;
	assign w_fld_a_0_datain_0 = 32'h0;
	assign w_fld_a_0_r_w_0 = 1'h0;
	assign w_fld_a_0_ce_0 = w_sys_ce;
	assign w_fld_a_0_ce_1 = w_sys_ce;
	assign w_fld_x_1_addr_0 = 7'sh0;
	assign w_fld_x_1_datain_0 = 32'h0;
	assign w_fld_x_1_r_w_0 = 1'h0;
	assign w_fld_x_1_ce_0 = w_sys_ce;
	assign w_fld_x_1_ce_1 = w_sys_ce;
	assign w_sub19_arrayA_addr = ( (|r_sys_processing_methodID) ? r_sub19_arrayA_addr : 3'sh0 ) ;
	assign w_sub19_arrayA_datain = ( (|r_sys_processing_methodID) ? r_sub19_arrayA_datain : 32'h0 ) ;
	assign w_sub19_arrayA_r_w = ( (|r_sys_processing_methodID) ? r_sub19_arrayA_r_w : 1'h0 ) ;
	assign w_sub19_arrayX_addr = ( (|r_sys_processing_methodID) ? r_sub19_arrayX_addr : 3'sh0 ) ;
	assign w_sub19_arrayX_datain = ( (|r_sys_processing_methodID) ? r_sub19_arrayX_datain : 32'h0 ) ;
	assign w_sub19_arrayX_r_w = ( (|r_sys_processing_methodID) ? r_sub19_arrayX_r_w : 1'h0 ) ;
	assign w_sub09_arrayA_addr = ( (|r_sys_processing_methodID) ? r_sub09_arrayA_addr : 3'sh0 ) ;
	assign w_sub09_arrayA_datain = ( (|r_sys_processing_methodID) ? r_sub09_arrayA_datain : 32'h0 ) ;
	assign w_sub09_arrayA_r_w = ( (|r_sys_processing_methodID) ? r_sub09_arrayA_r_w : 1'h0 ) ;
	assign w_sub09_arrayX_addr = ( (|r_sys_processing_methodID) ? r_sub09_arrayX_addr : 3'sh0 ) ;
	assign w_sub09_arrayX_datain = ( (|r_sys_processing_methodID) ? r_sub09_arrayX_datain : 32'h0 ) ;
	assign w_sub09_arrayX_r_w = ( (|r_sys_processing_methodID) ? r_sub09_arrayX_r_w : 1'h0 ) ;
	assign w_sub08_arrayA_addr = ( (|r_sys_processing_methodID) ? r_sub08_arrayA_addr : 3'sh0 ) ;
	assign w_sub08_arrayA_datain = ( (|r_sys_processing_methodID) ? r_sub08_arrayA_datain : 32'h0 ) ;
	assign w_sub08_arrayA_r_w = ( (|r_sys_processing_methodID) ? r_sub08_arrayA_r_w : 1'h0 ) ;
	assign w_sub08_arrayX_addr = ( (|r_sys_processing_methodID) ? r_sub08_arrayX_addr : 3'sh0 ) ;
	assign w_sub08_arrayX_datain = ( (|r_sys_processing_methodID) ? r_sub08_arrayX_datain : 32'h0 ) ;
	assign w_sub08_arrayX_r_w = ( (|r_sys_processing_methodID) ? r_sub08_arrayX_r_w : 1'h0 ) ;
	assign w_sub12_arrayA_addr = ( (|r_sys_processing_methodID) ? r_sub12_arrayA_addr : 3'sh0 ) ;
	assign w_sub12_arrayA_datain = ( (|r_sys_processing_methodID) ? r_sub12_arrayA_datain : 32'h0 ) ;
	assign w_sub12_arrayA_r_w = ( (|r_sys_processing_methodID) ? r_sub12_arrayA_r_w : 1'h0 ) ;
	assign w_sub12_arrayX_addr = ( (|r_sys_processing_methodID) ? r_sub12_arrayX_addr : 3'sh0 ) ;
	assign w_sub12_arrayX_datain = ( (|r_sys_processing_methodID) ? r_sub12_arrayX_datain : 32'h0 ) ;
	assign w_sub12_arrayX_r_w = ( (|r_sys_processing_methodID) ? r_sub12_arrayX_r_w : 1'h0 ) ;
	assign w_sub03_arrayA_addr = ( (|r_sys_processing_methodID) ? r_sub03_arrayA_addr : 3'sh0 ) ;
	assign w_sub03_arrayA_datain = ( (|r_sys_processing_methodID) ? r_sub03_arrayA_datain : 32'h0 ) ;
	assign w_sub03_arrayA_r_w = ( (|r_sys_processing_methodID) ? r_sub03_arrayA_r_w : 1'h0 ) ;
	assign w_sub03_arrayX_addr = ( (|r_sys_processing_methodID) ? r_sub03_arrayX_addr : 3'sh0 ) ;
	assign w_sub03_arrayX_datain = ( (|r_sys_processing_methodID) ? r_sub03_arrayX_datain : 32'h0 ) ;
	assign w_sub03_arrayX_r_w = ( (|r_sys_processing_methodID) ? r_sub03_arrayX_r_w : 1'h0 ) ;
	assign w_sub02_arrayA_addr = ( (|r_sys_processing_methodID) ? r_sub02_arrayA_addr : 3'sh0 ) ;
	assign w_sub02_arrayA_datain = ( (|r_sys_processing_methodID) ? r_sub02_arrayA_datain : 32'h0 ) ;
	assign w_sub02_arrayA_r_w = ( (|r_sys_processing_methodID) ? r_sub02_arrayA_r_w : 1'h0 ) ;
	assign w_sub02_arrayX_addr = ( (|r_sys_processing_methodID) ? r_sub02_arrayX_addr : 3'sh0 ) ;
	assign w_sub02_arrayX_datain = ( (|r_sys_processing_methodID) ? r_sub02_arrayX_datain : 32'h0 ) ;
	assign w_sub02_arrayX_r_w = ( (|r_sys_processing_methodID) ? r_sub02_arrayX_r_w : 1'h0 ) ;
	assign w_sub11_arrayA_addr = ( (|r_sys_processing_methodID) ? r_sub11_arrayA_addr : 3'sh0 ) ;
	assign w_sub11_arrayA_datain = ( (|r_sys_processing_methodID) ? r_sub11_arrayA_datain : 32'h0 ) ;
	assign w_sub11_arrayA_r_w = ( (|r_sys_processing_methodID) ? r_sub11_arrayA_r_w : 1'h0 ) ;
	assign w_sub11_arrayX_addr = ( (|r_sys_processing_methodID) ? r_sub11_arrayX_addr : 3'sh0 ) ;
	assign w_sub11_arrayX_datain = ( (|r_sys_processing_methodID) ? r_sub11_arrayX_datain : 32'h0 ) ;
	assign w_sub11_arrayX_r_w = ( (|r_sys_processing_methodID) ? r_sub11_arrayX_r_w : 1'h0 ) ;
	assign w_sub14_arrayA_addr = ( (|r_sys_processing_methodID) ? r_sub14_arrayA_addr : 3'sh0 ) ;
	assign w_sub14_arrayA_datain = ( (|r_sys_processing_methodID) ? r_sub14_arrayA_datain : 32'h0 ) ;
	assign w_sub14_arrayA_r_w = ( (|r_sys_processing_methodID) ? r_sub14_arrayA_r_w : 1'h0 ) ;
	assign w_sub14_arrayX_addr = ( (|r_sys_processing_methodID) ? r_sub14_arrayX_addr : 3'sh0 ) ;
	assign w_sub14_arrayX_datain = ( (|r_sys_processing_methodID) ? r_sub14_arrayX_datain : 32'h0 ) ;
	assign w_sub14_arrayX_r_w = ( (|r_sys_processing_methodID) ? r_sub14_arrayX_r_w : 1'h0 ) ;
	assign w_sub01_arrayA_addr = ( (|r_sys_processing_methodID) ? r_sub01_arrayA_addr : 3'sh0 ) ;
	assign w_sub01_arrayA_datain = ( (|r_sys_processing_methodID) ? r_sub01_arrayA_datain : 32'h0 ) ;
	assign w_sub01_arrayA_r_w = ( (|r_sys_processing_methodID) ? r_sub01_arrayA_r_w : 1'h0 ) ;
	assign w_sub01_arrayX_addr = ( (|r_sys_processing_methodID) ? r_sub01_arrayX_addr : 3'sh0 ) ;
	assign w_sub01_arrayX_datain = ( (|r_sys_processing_methodID) ? r_sub01_arrayX_datain : 32'h0 ) ;
	assign w_sub01_arrayX_r_w = ( (|r_sys_processing_methodID) ? r_sub01_arrayX_r_w : 1'h0 ) ;
	assign w_sub13_arrayA_addr = ( (|r_sys_processing_methodID) ? r_sub13_arrayA_addr : 3'sh0 ) ;
	assign w_sub13_arrayA_datain = ( (|r_sys_processing_methodID) ? r_sub13_arrayA_datain : 32'h0 ) ;
	assign w_sub13_arrayA_r_w = ( (|r_sys_processing_methodID) ? r_sub13_arrayA_r_w : 1'h0 ) ;
	assign w_sub13_arrayX_addr = ( (|r_sys_processing_methodID) ? r_sub13_arrayX_addr : 3'sh0 ) ;
	assign w_sub13_arrayX_datain = ( (|r_sys_processing_methodID) ? r_sub13_arrayX_datain : 32'h0 ) ;
	assign w_sub13_arrayX_r_w = ( (|r_sys_processing_methodID) ? r_sub13_arrayX_r_w : 1'h0 ) ;
	assign w_sub00_arrayA_addr = ( (|r_sys_processing_methodID) ? r_sub00_arrayA_addr : 3'sh0 ) ;
	assign w_sub00_arrayA_datain = ( (|r_sys_processing_methodID) ? r_sub00_arrayA_datain : 32'h0 ) ;
	assign w_sub00_arrayA_r_w = ( (|r_sys_processing_methodID) ? r_sub00_arrayA_r_w : 1'h0 ) ;
	assign w_sub00_arrayX_addr = ( (|r_sys_processing_methodID) ? r_sub00_arrayX_addr : 3'sh0 ) ;
	assign w_sub00_arrayX_datain = ( (|r_sys_processing_methodID) ? r_sub00_arrayX_datain : 32'h0 ) ;
	assign w_sub00_arrayX_r_w = ( (|r_sys_processing_methodID) ? r_sub00_arrayX_r_w : 1'h0 ) ;
	assign w_sub07_arrayA_addr = ( (|r_sys_processing_methodID) ? r_sub07_arrayA_addr : 3'sh0 ) ;
	assign w_sub07_arrayA_datain = ( (|r_sys_processing_methodID) ? r_sub07_arrayA_datain : 32'h0 ) ;
	assign w_sub07_arrayA_r_w = ( (|r_sys_processing_methodID) ? r_sub07_arrayA_r_w : 1'h0 ) ;
	assign w_sub07_arrayX_addr = ( (|r_sys_processing_methodID) ? r_sub07_arrayX_addr : 3'sh0 ) ;
	assign w_sub07_arrayX_datain = ( (|r_sys_processing_methodID) ? r_sub07_arrayX_datain : 32'h0 ) ;
	assign w_sub07_arrayX_r_w = ( (|r_sys_processing_methodID) ? r_sub07_arrayX_r_w : 1'h0 ) ;
	assign w_sub16_arrayA_addr = ( (|r_sys_processing_methodID) ? r_sub16_arrayA_addr : 3'sh0 ) ;
	assign w_sub16_arrayA_datain = ( (|r_sys_processing_methodID) ? r_sub16_arrayA_datain : 32'h0 ) ;
	assign w_sub16_arrayA_r_w = ( (|r_sys_processing_methodID) ? r_sub16_arrayA_r_w : 1'h0 ) ;
	assign w_sub16_arrayX_addr = ( (|r_sys_processing_methodID) ? r_sub16_arrayX_addr : 3'sh0 ) ;
	assign w_sub16_arrayX_datain = ( (|r_sys_processing_methodID) ? r_sub16_arrayX_datain : 32'h0 ) ;
	assign w_sub16_arrayX_r_w = ( (|r_sys_processing_methodID) ? r_sub16_arrayX_r_w : 1'h0 ) ;
	assign w_sub06_arrayA_addr = ( (|r_sys_processing_methodID) ? r_sub06_arrayA_addr : 3'sh0 ) ;
	assign w_sub06_arrayA_datain = ( (|r_sys_processing_methodID) ? r_sub06_arrayA_datain : 32'h0 ) ;
	assign w_sub06_arrayA_r_w = ( (|r_sys_processing_methodID) ? r_sub06_arrayA_r_w : 1'h0 ) ;
	assign w_sub06_arrayX_addr = ( (|r_sys_processing_methodID) ? r_sub06_arrayX_addr : 3'sh0 ) ;
	assign w_sub06_arrayX_datain = ( (|r_sys_processing_methodID) ? r_sub06_arrayX_datain : 32'h0 ) ;
	assign w_sub06_arrayX_r_w = ( (|r_sys_processing_methodID) ? r_sub06_arrayX_r_w : 1'h0 ) ;
	assign w_sub15_arrayA_addr = ( (|r_sys_processing_methodID) ? r_sub15_arrayA_addr : 3'sh0 ) ;
	assign w_sub15_arrayA_datain = ( (|r_sys_processing_methodID) ? r_sub15_arrayA_datain : 32'h0 ) ;
	assign w_sub15_arrayA_r_w = ( (|r_sys_processing_methodID) ? r_sub15_arrayA_r_w : 1'h0 ) ;
	assign w_sub15_arrayX_addr = ( (|r_sys_processing_methodID) ? r_sub15_arrayX_addr : 3'sh0 ) ;
	assign w_sub15_arrayX_datain = ( (|r_sys_processing_methodID) ? r_sub15_arrayX_datain : 32'h0 ) ;
	assign w_sub15_arrayX_r_w = ( (|r_sys_processing_methodID) ? r_sub15_arrayX_r_w : 1'h0 ) ;
	assign w_sub05_arrayA_addr = ( (|r_sys_processing_methodID) ? r_sub05_arrayA_addr : 3'sh0 ) ;
	assign w_sub05_arrayA_datain = ( (|r_sys_processing_methodID) ? r_sub05_arrayA_datain : 32'h0 ) ;
	assign w_sub05_arrayA_r_w = ( (|r_sys_processing_methodID) ? r_sub05_arrayA_r_w : 1'h0 ) ;
	assign w_sub05_arrayX_addr = ( (|r_sys_processing_methodID) ? r_sub05_arrayX_addr : 3'sh0 ) ;
	assign w_sub05_arrayX_datain = ( (|r_sys_processing_methodID) ? r_sub05_arrayX_datain : 32'h0 ) ;
	assign w_sub05_arrayX_r_w = ( (|r_sys_processing_methodID) ? r_sub05_arrayX_r_w : 1'h0 ) ;
	assign w_sub18_arrayA_addr = ( (|r_sys_processing_methodID) ? r_sub18_arrayA_addr : 3'sh0 ) ;
	assign w_sub18_arrayA_datain = ( (|r_sys_processing_methodID) ? r_sub18_arrayA_datain : 32'h0 ) ;
	assign w_sub18_arrayA_r_w = ( (|r_sys_processing_methodID) ? r_sub18_arrayA_r_w : 1'h0 ) ;
	assign w_sub18_arrayX_addr = ( (|r_sys_processing_methodID) ? r_sub18_arrayX_addr : 3'sh0 ) ;
	assign w_sub18_arrayX_datain = ( (|r_sys_processing_methodID) ? r_sub18_arrayX_datain : 32'h0 ) ;
	assign w_sub18_arrayX_r_w = ( (|r_sys_processing_methodID) ? r_sub18_arrayX_r_w : 1'h0 ) ;
	assign w_sub04_arrayA_addr = ( (|r_sys_processing_methodID) ? r_sub04_arrayA_addr : 3'sh0 ) ;
	assign w_sub04_arrayA_datain = ( (|r_sys_processing_methodID) ? r_sub04_arrayA_datain : 32'h0 ) ;
	assign w_sub04_arrayA_r_w = ( (|r_sys_processing_methodID) ? r_sub04_arrayA_r_w : 1'h0 ) ;
	assign w_sub04_arrayX_addr = ( (|r_sys_processing_methodID) ? r_sub04_arrayX_addr : 3'sh0 ) ;
	assign w_sub04_arrayX_datain = ( (|r_sys_processing_methodID) ? r_sub04_arrayX_datain : 32'h0 ) ;
	assign w_sub04_arrayX_r_w = ( (|r_sys_processing_methodID) ? r_sub04_arrayX_r_w : 1'h0 ) ;
	assign w_sub17_arrayA_addr = ( (|r_sys_processing_methodID) ? r_sub17_arrayA_addr : 3'sh0 ) ;
	assign w_sub17_arrayA_datain = ( (|r_sys_processing_methodID) ? r_sub17_arrayA_datain : 32'h0 ) ;
	assign w_sub17_arrayA_r_w = ( (|r_sys_processing_methodID) ? r_sub17_arrayA_r_w : 1'h0 ) ;
	assign w_sub17_arrayX_addr = ( (|r_sys_processing_methodID) ? r_sub17_arrayX_addr : 3'sh0 ) ;
	assign w_sub17_arrayX_datain = ( (|r_sys_processing_methodID) ? r_sub17_arrayX_datain : 32'h0 ) ;
	assign w_sub17_arrayX_r_w = ( (|r_sys_processing_methodID) ? r_sub17_arrayX_r_w : 1'h0 ) ;
	assign w_sub10_arrayA_addr = ( (|r_sys_processing_methodID) ? r_sub10_arrayA_addr : 3'sh0 ) ;
	assign w_sub10_arrayA_datain = ( (|r_sys_processing_methodID) ? r_sub10_arrayA_datain : 32'h0 ) ;
	assign w_sub10_arrayA_r_w = ( (|r_sys_processing_methodID) ? r_sub10_arrayA_r_w : 1'h0 ) ;
	assign w_sub10_arrayX_addr = ( (|r_sys_processing_methodID) ? r_sub10_arrayX_addr : 3'sh0 ) ;
	assign w_sub10_arrayX_datain = ( (|r_sys_processing_methodID) ? r_sub10_arrayX_datain : 32'h0 ) ;
	assign w_sub10_arrayX_r_w = ( (|r_sys_processing_methodID) ? r_sub10_arrayX_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'h3a83126f;
	assign w_sys_tmp2 = (r_run_j_25 < r_fld_N_2);
	assign w_sys_tmp5 = w_ip_FixedToFloat_floating_0;
	assign w_sys_tmp6 = $signed( w_ip_Multint_product_0[31:0] );
	assign w_sys_tmp7 = (r_run_j_25 + w_sys_intOne);
	assign w_sys_tmp8 = (r_run_t_26 < r_fld_end_3);
	assign w_sys_tmp9 = (r_run_t_26 + w_sys_intOne);
	assign w_sys_tmp10 = (r_run_i_27 < w_sys_tmp11);
	assign w_sys_tmp11 = 32'sh00000007;
	assign w_sys_tmp14 = w_fld_a_0_dataout_1;
	assign w_sys_tmp17 = (r_run_copy36_i_68 + w_sys_tmp18);
	assign w_sys_tmp18 = 32'sh00000004;
	assign w_sys_tmp21 = (r_run_copy34_i_66 + w_sys_tmp22);
	assign w_sys_tmp22 = 32'sh00000009;
	assign w_sys_tmp25 = (r_run_copy32_i_64 + w_sys_tmp26);
	assign w_sys_tmp26 = 32'sh0000000e;
	assign w_sys_tmp29 = (r_run_copy30_i_62 + w_sys_tmp30);
	assign w_sys_tmp30 = 32'sh00000013;
	assign w_sys_tmp33 = (r_run_copy28_i_60 + w_sys_tmp34);
	assign w_sys_tmp34 = 32'sh00000018;
	assign w_sys_tmp37 = (r_run_copy26_i_58 + w_sys_tmp38);
	assign w_sys_tmp38 = 32'sh0000001d;
	assign w_sys_tmp41 = (r_run_copy24_i_56 + w_sys_tmp42);
	assign w_sys_tmp42 = 32'sh00000022;
	assign w_sys_tmp45 = (r_run_copy22_i_54 + w_sys_tmp46);
	assign w_sys_tmp46 = 32'sh00000027;
	assign w_sys_tmp49 = (r_run_copy20_i_52 + w_sys_tmp50);
	assign w_sys_tmp50 = 32'sh0000002c;
	assign w_sys_tmp53 = (r_run_copy18_i_50 + w_sys_tmp54);
	assign w_sys_tmp54 = 32'sh00000031;
	assign w_sys_tmp57 = (r_run_copy16_i_48 + w_sys_tmp58);
	assign w_sys_tmp58 = 32'sh00000036;
	assign w_sys_tmp61 = (r_run_copy14_i_46 + w_sys_tmp62);
	assign w_sys_tmp62 = 32'sh0000003b;
	assign w_sys_tmp65 = (r_run_copy12_i_44 + w_sys_tmp66);
	assign w_sys_tmp66 = 32'sh00000040;
	assign w_sys_tmp69 = (r_run_copy10_i_42 + w_sys_tmp70);
	assign w_sys_tmp70 = 32'sh00000045;
	assign w_sys_tmp73 = (r_run_copy8_i_40 + w_sys_tmp74);
	assign w_sys_tmp74 = 32'sh0000004a;
	assign w_sys_tmp77 = (r_run_copy6_i_38 + w_sys_tmp78);
	assign w_sys_tmp78 = 32'sh0000004f;
	assign w_sys_tmp81 = (r_run_copy4_i_36 + w_sys_tmp82);
	assign w_sys_tmp82 = 32'sh00000054;
	assign w_sys_tmp85 = (r_run_copy2_i_34 + w_sys_tmp86);
	assign w_sys_tmp86 = 32'sh00000059;
	assign w_sys_tmp89 = (r_run_copy0_i_32 + w_sys_tmp90);
	assign w_sys_tmp90 = 32'sh0000005d;
	assign w_sys_tmp91 = (r_run_copy0_i_32 + w_sys_intOne);
	assign w_sys_tmp92 = (r_run_copy1_i_33 + w_sys_intOne);
	assign w_sys_tmp93 = (r_run_copy2_i_34 + w_sys_intOne);
	assign w_sys_tmp94 = (r_run_copy3_i_35 + w_sys_intOne);
	assign w_sys_tmp95 = (r_run_copy4_i_36 + w_sys_intOne);
	assign w_sys_tmp96 = (r_run_copy5_i_37 + w_sys_intOne);
	assign w_sys_tmp97 = (r_run_copy6_i_38 + w_sys_intOne);
	assign w_sys_tmp98 = (r_run_copy7_i_39 + w_sys_intOne);
	assign w_sys_tmp99 = (r_run_copy8_i_40 + w_sys_intOne);
	assign w_sys_tmp100 = (r_run_copy9_i_41 + w_sys_intOne);
	assign w_sys_tmp101 = (r_run_copy10_i_42 + w_sys_intOne);
	assign w_sys_tmp102 = (r_run_copy11_i_43 + w_sys_intOne);
	assign w_sys_tmp103 = (r_run_copy12_i_44 + w_sys_intOne);
	assign w_sys_tmp104 = (r_run_copy13_i_45 + w_sys_intOne);
	assign w_sys_tmp105 = (r_run_copy14_i_46 + w_sys_intOne);
	assign w_sys_tmp106 = (r_run_copy15_i_47 + w_sys_intOne);
	assign w_sys_tmp107 = (r_run_copy16_i_48 + w_sys_intOne);
	assign w_sys_tmp108 = (r_run_copy17_i_49 + w_sys_intOne);
	assign w_sys_tmp109 = (r_run_copy18_i_50 + w_sys_intOne);
	assign w_sys_tmp110 = (r_run_copy19_i_51 + w_sys_intOne);
	assign w_sys_tmp111 = (r_run_copy20_i_52 + w_sys_intOne);
	assign w_sys_tmp112 = (r_run_copy21_i_53 + w_sys_intOne);
	assign w_sys_tmp113 = (r_run_copy22_i_54 + w_sys_intOne);
	assign w_sys_tmp114 = (r_run_copy23_i_55 + w_sys_intOne);
	assign w_sys_tmp115 = (r_run_copy24_i_56 + w_sys_intOne);
	assign w_sys_tmp116 = (r_run_copy25_i_57 + w_sys_intOne);
	assign w_sys_tmp117 = (r_run_copy26_i_58 + w_sys_intOne);
	assign w_sys_tmp118 = (r_run_copy27_i_59 + w_sys_intOne);
	assign w_sys_tmp119 = (r_run_copy28_i_60 + w_sys_intOne);
	assign w_sys_tmp120 = (r_run_copy29_i_61 + w_sys_intOne);
	assign w_sys_tmp121 = (r_run_copy30_i_62 + w_sys_intOne);
	assign w_sys_tmp122 = (r_run_copy31_i_63 + w_sys_intOne);
	assign w_sys_tmp123 = (r_run_copy32_i_64 + w_sys_intOne);
	assign w_sys_tmp124 = (r_run_copy33_i_65 + w_sys_intOne);
	assign w_sys_tmp125 = (r_run_copy34_i_66 + w_sys_intOne);
	assign w_sys_tmp126 = (r_run_copy35_i_67 + w_sys_intOne);
	assign w_sys_tmp127 = (r_run_copy36_i_68 + w_sys_intOne);
	assign w_sys_tmp128 = (r_run_copy37_i_69 + w_sys_intOne);
	assign w_sys_tmp129 = (r_run_copy38_i_70 + w_sys_intOne);
	assign w_sys_tmp130 = (r_run_i_27 + w_sys_intOne);
	assign w_sys_tmp367 = 32'sh00000002;
	assign w_sys_tmp368 = (r_run_i_28 < w_sys_tmp369);
	assign w_sys_tmp369 = 32'sh00000005;
	assign w_sys_tmp374 = w_sub00_arrayX_dataout;
	assign w_sys_tmp376 = (r_run_copy18_i_89 + w_sys_tmp377);
	assign w_sys_tmp377 = 32'sh00000005;
	assign w_sys_tmp379 = (r_run_copy17_i_88 + w_sys_tmp380);
	assign w_sys_tmp380 = 32'sh0000000a;
	assign w_sys_tmp382 = (r_run_copy16_i_87 + w_sys_tmp383);
	assign w_sys_tmp383 = 32'sh0000000f;
	assign w_sys_tmp385 = (r_run_copy15_i_86 + w_sys_tmp386);
	assign w_sys_tmp386 = 32'sh00000014;
	assign w_sys_tmp388 = (r_run_copy14_i_85 + w_sys_tmp389);
	assign w_sys_tmp389 = 32'sh00000019;
	assign w_sys_tmp391 = (r_run_copy13_i_84 + w_sys_tmp392);
	assign w_sys_tmp392 = 32'sh0000001e;
	assign w_sys_tmp394 = (r_run_copy12_i_83 + w_sys_tmp395);
	assign w_sys_tmp395 = 32'sh00000023;
	assign w_sys_tmp397 = (r_run_copy11_i_82 + w_sys_tmp398);
	assign w_sys_tmp398 = 32'sh00000028;
	assign w_sys_tmp400 = (r_run_copy10_i_81 + w_sys_tmp401);
	assign w_sys_tmp401 = 32'sh0000002d;
	assign w_sys_tmp403 = (r_run_copy9_i_80 + w_sys_tmp404);
	assign w_sys_tmp404 = 32'sh00000032;
	assign w_sys_tmp406 = (r_run_copy8_i_79 + w_sys_tmp407);
	assign w_sys_tmp407 = 32'sh00000037;
	assign w_sys_tmp409 = (r_run_copy7_i_78 + w_sys_tmp410);
	assign w_sys_tmp410 = 32'sh0000003c;
	assign w_sys_tmp412 = (r_run_copy6_i_77 + w_sys_tmp413);
	assign w_sys_tmp413 = 32'sh00000041;
	assign w_sys_tmp415 = (r_run_copy5_i_76 + w_sys_tmp416);
	assign w_sys_tmp416 = 32'sh00000046;
	assign w_sys_tmp418 = (r_run_copy4_i_75 + w_sys_tmp419);
	assign w_sys_tmp419 = 32'sh0000004b;
	assign w_sys_tmp421 = (r_run_copy3_i_74 + w_sys_tmp422);
	assign w_sys_tmp422 = 32'sh00000050;
	assign w_sys_tmp424 = (r_run_copy2_i_73 + w_sys_tmp425);
	assign w_sys_tmp425 = 32'sh00000055;
	assign w_sys_tmp427 = (r_run_copy1_i_72 + w_sys_tmp428);
	assign w_sys_tmp428 = 32'sh0000005a;
	assign w_sys_tmp430 = (r_run_copy0_i_71 + w_sys_tmp431);
	assign w_sys_tmp431 = 32'sh0000005f;
	assign w_sys_tmp432 = (r_run_copy0_i_71 + w_sys_intOne);
	assign w_sys_tmp433 = (r_run_copy1_i_72 + w_sys_intOne);
	assign w_sys_tmp434 = (r_run_copy2_i_73 + w_sys_intOne);
	assign w_sys_tmp435 = (r_run_copy3_i_74 + w_sys_intOne);
	assign w_sys_tmp436 = (r_run_copy4_i_75 + w_sys_intOne);
	assign w_sys_tmp437 = (r_run_copy5_i_76 + w_sys_intOne);
	assign w_sys_tmp438 = (r_run_copy6_i_77 + w_sys_intOne);
	assign w_sys_tmp439 = (r_run_copy7_i_78 + w_sys_intOne);
	assign w_sys_tmp440 = (r_run_copy8_i_79 + w_sys_intOne);
	assign w_sys_tmp441 = (r_run_copy9_i_80 + w_sys_intOne);
	assign w_sys_tmp442 = (r_run_copy10_i_81 + w_sys_intOne);
	assign w_sys_tmp443 = (r_run_copy11_i_82 + w_sys_intOne);
	assign w_sys_tmp444 = (r_run_copy12_i_83 + w_sys_intOne);
	assign w_sys_tmp445 = (r_run_copy13_i_84 + w_sys_intOne);
	assign w_sys_tmp446 = (r_run_copy14_i_85 + w_sys_intOne);
	assign w_sys_tmp447 = (r_run_copy15_i_86 + w_sys_intOne);
	assign w_sys_tmp448 = (r_run_copy16_i_87 + w_sys_intOne);
	assign w_sys_tmp449 = (r_run_copy17_i_88 + w_sys_intOne);
	assign w_sys_tmp450 = (r_run_copy18_i_89 + w_sys_intOne);
	assign w_sys_tmp451 = (r_run_copy19_i_90 + w_sys_intOne);
	assign w_sys_tmp452 = (r_run_i_28 + w_sys_intOne);
	assign w_sys_tmp453 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp454 = (r_run_l_30 + w_sys_intOne);
	assign w_sys_tmp617 = (r_run_j_31 < r_fld_N_2);
	assign w_sys_tmp620 = w_fld_x_1_dataout_1;
	assign w_sys_tmp621 = (r_run_j_31 + w_sys_intOne);
	assign w_sys_tmp622 = 32'sh00000064;


	SubUnder
		sub19_inst(
			.i_fld_arrayA_0_addr_0 (w_sub19_arrayA_addr),
			.i_fld_arrayA_0_datain_0 (w_sub19_arrayA_datain),
			.o_fld_arrayA_0_dataout_0 (w_sub19_arrayA_dataout),
			.i_fld_arrayA_0_r_w_0 (w_sub19_arrayA_r_w),
			.i_fld_arrayX_1_addr_0 (w_sub19_arrayX_addr),
			.i_fld_arrayX_1_datain_0 (w_sub19_arrayX_datain),
			.o_fld_arrayX_1_dataout_0 (w_sub19_arrayX_dataout),
			.i_fld_arrayX_1_r_w_0 (w_sub19_arrayX_r_w),
			.o_run_busy (w_sub19_run_busy),
			.i_run_req (r_sub19_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	Sub
		sub09_inst(
			.i_fld_arrayA_0_addr_0 (w_sub09_arrayA_addr),
			.i_fld_arrayA_0_datain_0 (w_sub09_arrayA_datain),
			.o_fld_arrayA_0_dataout_0 (w_sub09_arrayA_dataout),
			.i_fld_arrayA_0_r_w_0 (w_sub09_arrayA_r_w),
			.i_fld_arrayX_1_addr_0 (w_sub09_arrayX_addr),
			.i_fld_arrayX_1_datain_0 (w_sub09_arrayX_datain),
			.o_fld_arrayX_1_dataout_0 (w_sub09_arrayX_dataout),
			.i_fld_arrayX_1_r_w_0 (w_sub09_arrayX_r_w),
			.o_run_busy (w_sub09_run_busy),
			.i_run_req (r_sub09_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	Sub
		sub08_inst(
			.i_fld_arrayA_0_addr_0 (w_sub08_arrayA_addr),
			.i_fld_arrayA_0_datain_0 (w_sub08_arrayA_datain),
			.o_fld_arrayA_0_dataout_0 (w_sub08_arrayA_dataout),
			.i_fld_arrayA_0_r_w_0 (w_sub08_arrayA_r_w),
			.i_fld_arrayX_1_addr_0 (w_sub08_arrayX_addr),
			.i_fld_arrayX_1_datain_0 (w_sub08_arrayX_datain),
			.o_fld_arrayX_1_dataout_0 (w_sub08_arrayX_dataout),
			.i_fld_arrayX_1_r_w_0 (w_sub08_arrayX_r_w),
			.o_run_busy (w_sub08_run_busy),
			.i_run_req (r_sub08_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	Sub
		sub12_inst(
			.i_fld_arrayA_0_addr_0 (w_sub12_arrayA_addr),
			.i_fld_arrayA_0_datain_0 (w_sub12_arrayA_datain),
			.o_fld_arrayA_0_dataout_0 (w_sub12_arrayA_dataout),
			.i_fld_arrayA_0_r_w_0 (w_sub12_arrayA_r_w),
			.i_fld_arrayX_1_addr_0 (w_sub12_arrayX_addr),
			.i_fld_arrayX_1_datain_0 (w_sub12_arrayX_datain),
			.o_fld_arrayX_1_dataout_0 (w_sub12_arrayX_dataout),
			.i_fld_arrayX_1_r_w_0 (w_sub12_arrayX_r_w),
			.o_run_busy (w_sub12_run_busy),
			.i_run_req (r_sub12_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	Sub
		sub03_inst(
			.i_fld_arrayA_0_addr_0 (w_sub03_arrayA_addr),
			.i_fld_arrayA_0_datain_0 (w_sub03_arrayA_datain),
			.o_fld_arrayA_0_dataout_0 (w_sub03_arrayA_dataout),
			.i_fld_arrayA_0_r_w_0 (w_sub03_arrayA_r_w),
			.i_fld_arrayX_1_addr_0 (w_sub03_arrayX_addr),
			.i_fld_arrayX_1_datain_0 (w_sub03_arrayX_datain),
			.o_fld_arrayX_1_dataout_0 (w_sub03_arrayX_dataout),
			.i_fld_arrayX_1_r_w_0 (w_sub03_arrayX_r_w),
			.o_run_busy (w_sub03_run_busy),
			.i_run_req (r_sub03_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	Sub
		sub02_inst(
			.i_fld_arrayA_0_addr_0 (w_sub02_arrayA_addr),
			.i_fld_arrayA_0_datain_0 (w_sub02_arrayA_datain),
			.o_fld_arrayA_0_dataout_0 (w_sub02_arrayA_dataout),
			.i_fld_arrayA_0_r_w_0 (w_sub02_arrayA_r_w),
			.i_fld_arrayX_1_addr_0 (w_sub02_arrayX_addr),
			.i_fld_arrayX_1_datain_0 (w_sub02_arrayX_datain),
			.o_fld_arrayX_1_dataout_0 (w_sub02_arrayX_dataout),
			.i_fld_arrayX_1_r_w_0 (w_sub02_arrayX_r_w),
			.o_run_busy (w_sub02_run_busy),
			.i_run_req (r_sub02_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	Sub
		sub11_inst(
			.i_fld_arrayA_0_addr_0 (w_sub11_arrayA_addr),
			.i_fld_arrayA_0_datain_0 (w_sub11_arrayA_datain),
			.o_fld_arrayA_0_dataout_0 (w_sub11_arrayA_dataout),
			.i_fld_arrayA_0_r_w_0 (w_sub11_arrayA_r_w),
			.i_fld_arrayX_1_addr_0 (w_sub11_arrayX_addr),
			.i_fld_arrayX_1_datain_0 (w_sub11_arrayX_datain),
			.o_fld_arrayX_1_dataout_0 (w_sub11_arrayX_dataout),
			.i_fld_arrayX_1_r_w_0 (w_sub11_arrayX_r_w),
			.o_run_busy (w_sub11_run_busy),
			.i_run_req (r_sub11_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	Sub
		sub14_inst(
			.i_fld_arrayA_0_addr_0 (w_sub14_arrayA_addr),
			.i_fld_arrayA_0_datain_0 (w_sub14_arrayA_datain),
			.o_fld_arrayA_0_dataout_0 (w_sub14_arrayA_dataout),
			.i_fld_arrayA_0_r_w_0 (w_sub14_arrayA_r_w),
			.i_fld_arrayX_1_addr_0 (w_sub14_arrayX_addr),
			.i_fld_arrayX_1_datain_0 (w_sub14_arrayX_datain),
			.o_fld_arrayX_1_dataout_0 (w_sub14_arrayX_dataout),
			.i_fld_arrayX_1_r_w_0 (w_sub14_arrayX_r_w),
			.o_run_busy (w_sub14_run_busy),
			.i_run_req (r_sub14_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	Sub
		sub01_inst(
			.i_fld_arrayA_0_addr_0 (w_sub01_arrayA_addr),
			.i_fld_arrayA_0_datain_0 (w_sub01_arrayA_datain),
			.o_fld_arrayA_0_dataout_0 (w_sub01_arrayA_dataout),
			.i_fld_arrayA_0_r_w_0 (w_sub01_arrayA_r_w),
			.i_fld_arrayX_1_addr_0 (w_sub01_arrayX_addr),
			.i_fld_arrayX_1_datain_0 (w_sub01_arrayX_datain),
			.o_fld_arrayX_1_dataout_0 (w_sub01_arrayX_dataout),
			.i_fld_arrayX_1_r_w_0 (w_sub01_arrayX_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	Sub
		sub13_inst(
			.i_fld_arrayA_0_addr_0 (w_sub13_arrayA_addr),
			.i_fld_arrayA_0_datain_0 (w_sub13_arrayA_datain),
			.o_fld_arrayA_0_dataout_0 (w_sub13_arrayA_dataout),
			.i_fld_arrayA_0_r_w_0 (w_sub13_arrayA_r_w),
			.i_fld_arrayX_1_addr_0 (w_sub13_arrayX_addr),
			.i_fld_arrayX_1_datain_0 (w_sub13_arrayX_datain),
			.o_fld_arrayX_1_dataout_0 (w_sub13_arrayX_dataout),
			.i_fld_arrayX_1_r_w_0 (w_sub13_arrayX_r_w),
			.o_run_busy (w_sub13_run_busy),
			.i_run_req (r_sub13_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	SubUp
		sub00_inst(
			.i_fld_arrayA_0_addr_0 (w_sub00_arrayA_addr),
			.i_fld_arrayA_0_datain_0 (w_sub00_arrayA_datain),
			.o_fld_arrayA_0_dataout_0 (w_sub00_arrayA_dataout),
			.i_fld_arrayA_0_r_w_0 (w_sub00_arrayA_r_w),
			.i_fld_arrayX_1_addr_0 (w_sub00_arrayX_addr),
			.i_fld_arrayX_1_datain_0 (w_sub00_arrayX_datain),
			.o_fld_arrayX_1_dataout_0 (w_sub00_arrayX_dataout),
			.i_fld_arrayX_1_r_w_0 (w_sub00_arrayX_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	Sub
		sub07_inst(
			.i_fld_arrayA_0_addr_0 (w_sub07_arrayA_addr),
			.i_fld_arrayA_0_datain_0 (w_sub07_arrayA_datain),
			.o_fld_arrayA_0_dataout_0 (w_sub07_arrayA_dataout),
			.i_fld_arrayA_0_r_w_0 (w_sub07_arrayA_r_w),
			.i_fld_arrayX_1_addr_0 (w_sub07_arrayX_addr),
			.i_fld_arrayX_1_datain_0 (w_sub07_arrayX_datain),
			.o_fld_arrayX_1_dataout_0 (w_sub07_arrayX_dataout),
			.i_fld_arrayX_1_r_w_0 (w_sub07_arrayX_r_w),
			.o_run_busy (w_sub07_run_busy),
			.i_run_req (r_sub07_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	Sub
		sub16_inst(
			.i_fld_arrayA_0_addr_0 (w_sub16_arrayA_addr),
			.i_fld_arrayA_0_datain_0 (w_sub16_arrayA_datain),
			.o_fld_arrayA_0_dataout_0 (w_sub16_arrayA_dataout),
			.i_fld_arrayA_0_r_w_0 (w_sub16_arrayA_r_w),
			.i_fld_arrayX_1_addr_0 (w_sub16_arrayX_addr),
			.i_fld_arrayX_1_datain_0 (w_sub16_arrayX_datain),
			.o_fld_arrayX_1_dataout_0 (w_sub16_arrayX_dataout),
			.i_fld_arrayX_1_r_w_0 (w_sub16_arrayX_r_w),
			.o_run_busy (w_sub16_run_busy),
			.i_run_req (r_sub16_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	Sub
		sub06_inst(
			.i_fld_arrayA_0_addr_0 (w_sub06_arrayA_addr),
			.i_fld_arrayA_0_datain_0 (w_sub06_arrayA_datain),
			.o_fld_arrayA_0_dataout_0 (w_sub06_arrayA_dataout),
			.i_fld_arrayA_0_r_w_0 (w_sub06_arrayA_r_w),
			.i_fld_arrayX_1_addr_0 (w_sub06_arrayX_addr),
			.i_fld_arrayX_1_datain_0 (w_sub06_arrayX_datain),
			.o_fld_arrayX_1_dataout_0 (w_sub06_arrayX_dataout),
			.i_fld_arrayX_1_r_w_0 (w_sub06_arrayX_r_w),
			.o_run_busy (w_sub06_run_busy),
			.i_run_req (r_sub06_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	Sub
		sub15_inst(
			.i_fld_arrayA_0_addr_0 (w_sub15_arrayA_addr),
			.i_fld_arrayA_0_datain_0 (w_sub15_arrayA_datain),
			.o_fld_arrayA_0_dataout_0 (w_sub15_arrayA_dataout),
			.i_fld_arrayA_0_r_w_0 (w_sub15_arrayA_r_w),
			.i_fld_arrayX_1_addr_0 (w_sub15_arrayX_addr),
			.i_fld_arrayX_1_datain_0 (w_sub15_arrayX_datain),
			.o_fld_arrayX_1_dataout_0 (w_sub15_arrayX_dataout),
			.i_fld_arrayX_1_r_w_0 (w_sub15_arrayX_r_w),
			.o_run_busy (w_sub15_run_busy),
			.i_run_req (r_sub15_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	Sub
		sub05_inst(
			.i_fld_arrayA_0_addr_0 (w_sub05_arrayA_addr),
			.i_fld_arrayA_0_datain_0 (w_sub05_arrayA_datain),
			.o_fld_arrayA_0_dataout_0 (w_sub05_arrayA_dataout),
			.i_fld_arrayA_0_r_w_0 (w_sub05_arrayA_r_w),
			.i_fld_arrayX_1_addr_0 (w_sub05_arrayX_addr),
			.i_fld_arrayX_1_datain_0 (w_sub05_arrayX_datain),
			.o_fld_arrayX_1_dataout_0 (w_sub05_arrayX_dataout),
			.i_fld_arrayX_1_r_w_0 (w_sub05_arrayX_r_w),
			.o_run_busy (w_sub05_run_busy),
			.i_run_req (r_sub05_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	Sub
		sub18_inst(
			.i_fld_arrayA_0_addr_0 (w_sub18_arrayA_addr),
			.i_fld_arrayA_0_datain_0 (w_sub18_arrayA_datain),
			.o_fld_arrayA_0_dataout_0 (w_sub18_arrayA_dataout),
			.i_fld_arrayA_0_r_w_0 (w_sub18_arrayA_r_w),
			.i_fld_arrayX_1_addr_0 (w_sub18_arrayX_addr),
			.i_fld_arrayX_1_datain_0 (w_sub18_arrayX_datain),
			.o_fld_arrayX_1_dataout_0 (w_sub18_arrayX_dataout),
			.i_fld_arrayX_1_r_w_0 (w_sub18_arrayX_r_w),
			.o_run_busy (w_sub18_run_busy),
			.i_run_req (r_sub18_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	Sub
		sub04_inst(
			.i_fld_arrayA_0_addr_0 (w_sub04_arrayA_addr),
			.i_fld_arrayA_0_datain_0 (w_sub04_arrayA_datain),
			.o_fld_arrayA_0_dataout_0 (w_sub04_arrayA_dataout),
			.i_fld_arrayA_0_r_w_0 (w_sub04_arrayA_r_w),
			.i_fld_arrayX_1_addr_0 (w_sub04_arrayX_addr),
			.i_fld_arrayX_1_datain_0 (w_sub04_arrayX_datain),
			.o_fld_arrayX_1_dataout_0 (w_sub04_arrayX_dataout),
			.i_fld_arrayX_1_r_w_0 (w_sub04_arrayX_r_w),
			.o_run_busy (w_sub04_run_busy),
			.i_run_req (r_sub04_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	Sub
		sub17_inst(
			.i_fld_arrayA_0_addr_0 (w_sub17_arrayA_addr),
			.i_fld_arrayA_0_datain_0 (w_sub17_arrayA_datain),
			.o_fld_arrayA_0_dataout_0 (w_sub17_arrayA_dataout),
			.i_fld_arrayA_0_r_w_0 (w_sub17_arrayA_r_w),
			.i_fld_arrayX_1_addr_0 (w_sub17_arrayX_addr),
			.i_fld_arrayX_1_datain_0 (w_sub17_arrayX_datain),
			.o_fld_arrayX_1_dataout_0 (w_sub17_arrayX_dataout),
			.i_fld_arrayX_1_r_w_0 (w_sub17_arrayX_r_w),
			.o_run_busy (w_sub17_run_busy),
			.i_run_req (r_sub17_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	Sub
		sub10_inst(
			.i_fld_arrayA_0_addr_0 (w_sub10_arrayA_addr),
			.i_fld_arrayA_0_datain_0 (w_sub10_arrayA_datain),
			.o_fld_arrayA_0_dataout_0 (w_sub10_arrayA_dataout),
			.i_fld_arrayA_0_r_w_0 (w_sub10_arrayA_r_w),
			.i_fld_arrayX_1_addr_0 (w_sub10_arrayX_addr),
			.i_fld_arrayX_1_datain_0 (w_sub10_arrayX_datain),
			.o_fld_arrayX_1_dataout_0 (w_sub10_arrayX_dataout),
			.i_fld_arrayX_1_r_w_0 (w_sub10_arrayX_r_w),
			.o_run_busy (w_sub10_run_busy),
			.i_run_req (r_sub10_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(7), .WORDS(100) )
		dpram_a_0(
			.clk (clock),
			.ce_0 (w_fld_a_0_ce_0),
			.addr_0 (w_fld_a_0_addr_0),
			.datain_0 (w_fld_a_0_datain_0),
			.dataout_0 (w_fld_a_0_dataout_0),
			.r_w_0 (w_fld_a_0_r_w_0),
			.ce_1 (w_fld_a_0_ce_1),
			.addr_1 (r_fld_a_0_addr_1),
			.datain_1 (r_fld_a_0_datain_1),
			.dataout_1 (w_fld_a_0_dataout_1),
			.r_w_1 (r_fld_a_0_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(7), .WORDS(100) )
		dpram_x_1(
			.clk (clock),
			.ce_0 (w_fld_x_1_ce_0),
			.addr_0 (w_fld_x_1_addr_0),
			.datain_0 (w_fld_x_1_datain_0),
			.dataout_0 (w_fld_x_1_dataout_0),
			.r_w_0 (w_fld_x_1_r_w_0),
			.ce_1 (w_fld_x_1_ce_1),
			.addr_1 (r_fld_x_1_addr_1),
			.datain_1 (r_fld_x_1_datain_1),
			.dataout_1 (w_fld_x_1_dataout_1),
			.r_w_1 (r_fld_x_1_r_w_1)
		);

	Multint
		Multint_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_Multint_multiplicand_0),
			.b (r_ip_Multint_multiplier_0),
			.p (w_ip_Multint_product_0)
		);

	FixedToFloat
		FixedToFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_FixedToFloat_fixed_0),
			.result (w_ip_FixedToFloat_floating_0)
		);

	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_ip_Multint_multiplicand_0 <= r_run_j_25;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_ip_Multint_multiplier_0 <= r_run_j_25;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5)) begin
										r_ip_FixedToFloat_fixed_0 <= w_sys_tmp6;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 6'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_phase <= 6'h2;
						end

						6'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 6'h4;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2) ? 6'h8 : 6'ha);

									end
								end

							endcase
						end

						6'h8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hc)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 6'hb;

									end
								end

							endcase
						end

						6'hb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp8) ? 6'hf : 6'h24);

									end
								end

							endcase
						end

						6'hc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 6'hb;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 6'h10;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp10) ? 6'h13 : 6'h14);

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 6'h10;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h13: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_phase <= 6'h16;

									end
								end

							endcase
						end

						6'h16: begin

							case(r_sys_run_stage) 
								5'h13: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_phase <= 6'h18;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 6'h19;

									end
								end

							endcase
						end

						6'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp368) ? 6'h1c : 6'h1e);

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 6'h19;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 6'h1f;

									end
								end

							endcase
						end

						6'h1f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp617) ? 6'h22 : 6'hc);

									end
								end

							endcase
						end

						6'h22: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_run_phase <= 6'h1f;

									end
								end

							endcase
						end

						6'h24: begin
							r_sys_run_phase <= 6'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 5'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hc)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'hb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'hc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h16: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h1f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h22: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 6'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hc)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'hb)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'hb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'hc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h16: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub00_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub01_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub02_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub03_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub04_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub05_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub06_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub07_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub08_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub09_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub10_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub11_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub12_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub13_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub14_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub15_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub16_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub17_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub18_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub19_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h1f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h22: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						6'h24: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_a_0_addr_1 <= 7'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hc)) begin
										r_fld_a_0_addr_1 <= $signed( r_run_j_25[6:0] );

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h30)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp45[6:0] );

									end
									else
									if((r_sys_run_step==6'h10) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h38)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp77[6:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h2a)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp21[6:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h2e)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp37[6:0] );

									end
									else
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h2f)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp41[6:0] );

									end
									else
									if((r_sys_run_step==6'hf) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h37)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp73[6:0] );

									end
									else
									if((r_sys_run_step==6'hc) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h34)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp61[6:0] );

									end
									else
									if((r_sys_run_step==6'h4) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h2c)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp29[6:0] );

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h32)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp53[6:0] );

									end
									else
									if((r_sys_run_step==6'h11) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h39)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp81[6:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h31)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp49[6:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h28)) begin
										r_fld_a_0_addr_1 <= $signed( r_run_copy38_i_70[6:0] );

									end
									else
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h33)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp57[6:0] );

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h35)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp65[6:0] );

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h2b)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp25[6:0] );

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h2d)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp33[6:0] );

									end
									else
									if((r_sys_run_step==6'h13) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h3b)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp89[6:0] );

									end
									else
									if((r_sys_run_step==6'h1) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h29)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp17[6:0] );

									end
									else
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h36)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp69[6:0] );

									end
									else
									if((r_sys_run_step==6'h12) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h3a)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp85[6:0] );

									end
								end

							endcase
						end

						6'h22: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_fld_a_0_addr_1 <= $signed( r_run_j_31[6:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hc)) begin
										r_fld_a_0_datain_1 <= w_sys_tmp5;

									end
								end

							endcase
						end

						6'h22: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_fld_a_0_datain_1 <= w_sys_tmp620;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_a_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hc)) begin
										r_fld_a_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3b)) begin
										r_fld_a_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h22: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_fld_a_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h24: begin
							r_fld_a_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_x_1_addr_1 <= 7'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hc) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h34)) begin
										r_fld_x_1_addr_1 <= $signed( w_sys_tmp403[6:0] );

									end
									else
									if((r_sys_run_step==6'h10) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h38)) begin
										r_fld_x_1_addr_1 <= $signed( w_sys_tmp415[6:0] );

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h32)) begin
										r_fld_x_1_addr_1 <= $signed( w_sys_tmp397[6:0] );

									end
									else
									if((r_sys_run_step==6'h4) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h2c)) begin
										r_fld_x_1_addr_1 <= $signed( w_sys_tmp379[6:0] );

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h2d)) begin
										r_fld_x_1_addr_1 <= $signed( w_sys_tmp382[6:0] );

									end
									else
									if((r_sys_run_step==6'h15) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h3d)) begin
										r_fld_x_1_addr_1 <= $signed( w_sys_tmp430[6:0] );

									end
									else
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h36)) begin
										r_fld_x_1_addr_1 <= $signed( w_sys_tmp409[6:0] );

									end
									else
									if((r_sys_run_step==6'h8) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h30)) begin
										r_fld_x_1_addr_1 <= $signed( w_sys_tmp391[6:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h2a)) begin
										r_fld_x_1_addr_1 <= $signed( r_run_i_28[6:0] );

									end
									else
									if((r_sys_run_step==6'hf) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h37)) begin
										r_fld_x_1_addr_1 <= $signed( w_sys_tmp412[6:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h2e)) begin
										r_fld_x_1_addr_1 <= $signed( w_sys_tmp385[6:0] );

									end
									else
									if((r_sys_run_step==6'h11) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h39)) begin
										r_fld_x_1_addr_1 <= $signed( w_sys_tmp418[6:0] );

									end
									else
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h33)) begin
										r_fld_x_1_addr_1 <= $signed( w_sys_tmp400[6:0] );

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h2b)) begin
										r_fld_x_1_addr_1 <= $signed( w_sys_tmp376[6:0] );

									end
									else
									if((r_sys_run_step==6'h14) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h3c)) begin
										r_fld_x_1_addr_1 <= $signed( w_sys_tmp427[6:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h31)) begin
										r_fld_x_1_addr_1 <= $signed( w_sys_tmp394[6:0] );

									end
									else
									if((r_sys_run_step==6'h13) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h3b)) begin
										r_fld_x_1_addr_1 <= $signed( w_sys_tmp424[6:0] );

									end
									else
									if((r_sys_run_step==6'h12) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h3a)) begin
										r_fld_x_1_addr_1 <= $signed( w_sys_tmp421[6:0] );

									end
									else
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h2f)) begin
										r_fld_x_1_addr_1 <= $signed( w_sys_tmp388[6:0] );

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h35)) begin
										r_fld_x_1_addr_1 <= $signed( w_sys_tmp406[6:0] );

									end
								end

							endcase
						end

						6'h22: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_fld_x_1_addr_1 <= $signed( r_run_j_31[6:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp53_float;

									end
									else
									if((r_sys_run_step==6'h1c)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp22_float;

									end
									else
									if((r_sys_run_step==6'he)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp42_float;

									end
									else
									if((r_sys_run_step==6'h32)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==6'h2d)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp52_float;

									end
									else
									if((r_sys_run_step==6'h1f)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp36_float;

									end
									else
									if((r_sys_run_step==6'h25)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp31_float;

									end
									else
									if((r_sys_run_step==6'h3b)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==6'h12)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp44_float;

									end
									else
									if((r_sys_run_step==6'h19)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp24_float;

									end
									else
									if((r_sys_run_step==6'h31)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==6'h21)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp34_float;

									end
									else
									if((r_sys_run_step==6'h3d)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp14_float;

									end
									else
									if((r_sys_run_step==6'h38)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp18_float;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp38_float;

									end
									else
									if((r_sys_run_step==6'h2b)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_fld_x_1_datain_1 <= w_sys_tmp374;

									end
									else
									if((r_sys_run_step==6'h13)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp47_float;

									end
									else
									if((r_sys_run_step==6'h36)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==6'h18)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp20_float;

									end
									else
									if((r_sys_run_step==6'h16)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp19_float;

									end
									else
									if((r_sys_run_step==6'h14)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp45_float;

									end
									else
									if((r_sys_run_step==6'h37)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==6'h2a)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h3c)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==6'hf)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp49_float;

									end
									else
									if((r_sys_run_step==6'h23)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp33_float;

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp40_float;

									end
									else
									if((r_sys_run_step==6'h26)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp27_float;

									end
									else
									if((r_sys_run_step==6'h39)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==6'h1e)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp25_float;

									end
									else
									if((r_sys_run_step==6'h11)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp48_float;

									end
									else
									if((r_sys_run_step==6'h1b)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp23_float;

									end
									else
									if((r_sys_run_step==6'h24)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp32_float;

									end
									else
									if((r_sys_run_step==6'h20)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp35_float;

									end
									else
									if((r_sys_run_step==6'h22)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp26_float;

									end
									else
									if((r_sys_run_step==6'hc)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp41_float;

									end
									else
									if((r_sys_run_step==6'h1d)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp37_float;

									end
									else
									if((r_sys_run_step==6'h10)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp43_float;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp39_float;

									end
									else
									if((r_sys_run_step==6'h29)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp28_float;

									end
									else
									if((r_sys_run_step==6'hb)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp51_float;

									end
									else
									if((r_sys_run_step==6'h28)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp29_float;

									end
									else
									if((r_sys_run_step==6'h2f)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h17)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp55_float;

									end
									else
									if((r_sys_run_step==6'h4) || (r_sys_run_step==6'h2c)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp56_float;

									end
									else
									if((r_sys_run_step==6'h3a)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==6'h15)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp46_float;

									end
									else
									if((r_sys_run_step==6'h1a)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp21_float;

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp54_float;

									end
									else
									if((r_sys_run_step==6'h35)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==6'h33)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==6'h30)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==6'h34)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp50_float;

									end
									else
									if((r_sys_run_step==6'h27)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp30_float;

									end
									else
									if((r_sys_run_step==6'h2e)) begin
										r_fld_x_1_datain_1 <= r_sys_tmp3_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_x_1_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h3d)) begin
										r_fld_x_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h22: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_fld_x_1_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_fld_x_1_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_N_2 <= w_sys_tmp622;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_end_3 <= w_sys_intOne;

		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_r_24 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_25 <= w_sys_intZero;

									end
								end

							endcase
						end

						6'h8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hc)) begin
										r_run_j_25 <= w_sys_tmp7;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_t_26 <= w_sys_intZero;

									end
								end

							endcase
						end

						6'hc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_t_26 <= w_sys_tmp9;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_i_27 <= w_sys_intZero;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h2a)) begin
										r_run_i_27 <= w_sys_tmp130;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_i_28 <= w_sys_intZero;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h2a)) begin
										r_run_i_28 <= w_sys_tmp452;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_29 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_run_k_29 <= w_sys_tmp453;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_l_30 <= w_sys_tmp367;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_run_l_30 <= w_sys_tmp454;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_31 <= w_sys_intZero;

									end
								end

							endcase
						end

						6'h22: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_run_j_31 <= w_sys_tmp621;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_i_32 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h13) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_i_32 <= w_sys_tmp91;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_i_33 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h15) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_i_33 <= w_sys_tmp92;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_i_34 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h12) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h3a)) begin
										r_run_copy2_i_34 <= w_sys_tmp93;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_i_35 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h14) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h3c)) begin
										r_run_copy3_i_35 <= w_sys_tmp94;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_i_36 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h11) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h39)) begin
										r_run_copy4_i_36 <= w_sys_tmp95;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_i_37 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h13) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h3b)) begin
										r_run_copy5_i_37 <= w_sys_tmp96;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_i_38 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h10) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h38)) begin
										r_run_copy6_i_38 <= w_sys_tmp97;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_i_39 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h12) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h3a)) begin
										r_run_copy7_i_39 <= w_sys_tmp98;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_i_40 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hf) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h37)) begin
										r_run_copy8_i_40 <= w_sys_tmp99;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_i_41 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h11) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h39)) begin
										r_run_copy9_i_41 <= w_sys_tmp100;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_i_42 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h36)) begin
										r_run_copy10_i_42 <= w_sys_tmp101;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy11_i_43 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h10) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h38)) begin
										r_run_copy11_i_43 <= w_sys_tmp102;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy12_i_44 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h35)) begin
										r_run_copy12_i_44 <= w_sys_tmp103;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy13_i_45 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hf) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h37)) begin
										r_run_copy13_i_45 <= w_sys_tmp104;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy14_i_46 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hc) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h34)) begin
										r_run_copy14_i_46 <= w_sys_tmp105;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy15_i_47 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h36)) begin
										r_run_copy15_i_47 <= w_sys_tmp106;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy16_i_48 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h33)) begin
										r_run_copy16_i_48 <= w_sys_tmp107;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy17_i_49 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h35)) begin
										r_run_copy17_i_49 <= w_sys_tmp108;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy18_i_50 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h32)) begin
										r_run_copy18_i_50 <= w_sys_tmp109;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy19_i_51 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hc) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h34)) begin
										r_run_copy19_i_51 <= w_sys_tmp110;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy20_i_52 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h31)) begin
										r_run_copy20_i_52 <= w_sys_tmp111;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy21_i_53 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h33)) begin
										r_run_copy21_i_53 <= w_sys_tmp112;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy22_i_54 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h30)) begin
										r_run_copy22_i_54 <= w_sys_tmp113;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy23_i_55 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h32)) begin
										r_run_copy23_i_55 <= w_sys_tmp114;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy24_i_56 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h2f)) begin
										r_run_copy24_i_56 <= w_sys_tmp115;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy25_i_57 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h31)) begin
										r_run_copy25_i_57 <= w_sys_tmp116;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy26_i_58 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h2e)) begin
										r_run_copy26_i_58 <= w_sys_tmp117;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy27_i_59 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h30)) begin
										r_run_copy27_i_59 <= w_sys_tmp118;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy28_i_60 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h2d)) begin
										r_run_copy28_i_60 <= w_sys_tmp119;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy29_i_61 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h2f)) begin
										r_run_copy29_i_61 <= w_sys_tmp120;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy30_i_62 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h2c)) begin
										r_run_copy30_i_62 <= w_sys_tmp121;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy31_i_63 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h2e)) begin
										r_run_copy31_i_63 <= w_sys_tmp122;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy32_i_64 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h2b)) begin
										r_run_copy32_i_64 <= w_sys_tmp123;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy33_i_65 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h2d)) begin
										r_run_copy33_i_65 <= w_sys_tmp124;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy34_i_66 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h2a)) begin
										r_run_copy34_i_66 <= w_sys_tmp125;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy35_i_67 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h2c)) begin
										r_run_copy35_i_67 <= w_sys_tmp126;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy36_i_68 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h29)) begin
										r_run_copy36_i_68 <= w_sys_tmp127;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy37_i_69 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h2b)) begin
										r_run_copy37_i_69 <= w_sys_tmp128;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy38_i_70 <= r_run_i_27;

									end
								end

							endcase
						end

						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h28)) begin
										r_run_copy38_i_70 <= w_sys_tmp129;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h18: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_i_71 <= r_run_i_28;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h15) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h3d)) begin
										r_run_copy0_i_71 <= w_sys_tmp432;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h18: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_i_72 <= r_run_i_28;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h14) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h3c)) begin
										r_run_copy1_i_72 <= w_sys_tmp433;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h18: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_i_73 <= r_run_i_28;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h13) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h3b)) begin
										r_run_copy2_i_73 <= w_sys_tmp434;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h18: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_i_74 <= r_run_i_28;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h12) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_i_74 <= w_sys_tmp435;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h18: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_i_75 <= r_run_i_28;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h11) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h39)) begin
										r_run_copy4_i_75 <= w_sys_tmp436;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h18: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_i_76 <= r_run_i_28;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h10) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h38)) begin
										r_run_copy5_i_76 <= w_sys_tmp437;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h18: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_i_77 <= r_run_i_28;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hf) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h37)) begin
										r_run_copy6_i_77 <= w_sys_tmp438;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h18: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_i_78 <= r_run_i_28;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_i_78 <= w_sys_tmp439;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h18: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_i_79 <= r_run_i_28;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h35)) begin
										r_run_copy8_i_79 <= w_sys_tmp440;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h18: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_i_80 <= r_run_i_28;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hc) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h34)) begin
										r_run_copy9_i_80 <= w_sys_tmp441;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h18: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_i_81 <= r_run_i_28;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h33)) begin
										r_run_copy10_i_81 <= w_sys_tmp442;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h18: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy11_i_82 <= r_run_i_28;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h32)) begin
										r_run_copy11_i_82 <= w_sys_tmp443;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h18: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy12_i_83 <= r_run_i_28;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h31)) begin
										r_run_copy12_i_83 <= w_sys_tmp444;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h18: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy13_i_84 <= r_run_i_28;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h30)) begin
										r_run_copy13_i_84 <= w_sys_tmp445;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h18: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy14_i_85 <= r_run_i_28;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h2f)) begin
										r_run_copy14_i_85 <= w_sys_tmp446;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h18: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy15_i_86 <= r_run_i_28;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h2e)) begin
										r_run_copy15_i_86 <= w_sys_tmp447;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h18: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy16_i_87 <= r_run_i_28;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h2d)) begin
										r_run_copy16_i_87 <= w_sys_tmp448;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h18: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy17_i_88 <= r_run_i_28;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h2c)) begin
										r_run_copy17_i_88 <= w_sys_tmp449;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h18: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy18_i_89 <= r_run_i_28;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h2b)) begin
										r_run_copy18_i_89 <= w_sys_tmp450;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h18: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy19_i_90 <= r_run_i_28;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_run_copy19_i_90 <= w_sys_tmp451;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h13: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub19_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub19_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_arrayA_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h15) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h3d)) begin
										r_sub19_arrayA_addr <= $signed( r_run_copy1_i_33[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h15) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h3d)) begin
										r_sub19_arrayA_datain <= w_sys_tmp14;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_arrayA_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h15) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h3d)) begin
										r_sub19_arrayA_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayA_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub19_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_arrayX_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub19_arrayX_addr <= $signed( r_run_l_30[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_arrayX_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub19_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub19_arrayX_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h9: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub09_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub09_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_arrayA_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h33)) begin
										r_sub09_arrayA_addr <= $signed( r_run_copy21_i_53[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h33)) begin
										r_sub09_arrayA_datain <= w_sys_tmp14;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_arrayA_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h33)) begin
										r_sub09_arrayA_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayA_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub09_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_arrayX_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub09_arrayX_addr <= $signed( r_run_k_29[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_arrayX_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub09_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub09_arrayX_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub08_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub08_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_arrayA_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h32)) begin
										r_sub08_arrayA_addr <= $signed( r_run_copy23_i_55[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h32)) begin
										r_sub08_arrayA_datain <= w_sys_tmp14;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_arrayA_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h32)) begin
										r_sub08_arrayA_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayA_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub08_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_arrayX_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub08_arrayX_addr <= $signed( r_run_k_29[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_arrayX_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub08_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub08_arrayX_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub12_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub12_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_arrayA_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h36)) begin
										r_sub12_arrayA_addr <= $signed( r_run_copy15_i_47[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h36)) begin
										r_sub12_arrayA_datain <= w_sys_tmp14;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_arrayA_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h36)) begin
										r_sub12_arrayA_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayA_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub12_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_arrayX_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub12_arrayX_addr <= $signed( r_run_k_29[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_arrayX_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub12_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub12_arrayX_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_arrayA_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h2d)) begin
										r_sub03_arrayA_addr <= $signed( r_run_copy33_i_65[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h2d)) begin
										r_sub03_arrayA_datain <= w_sys_tmp14;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_arrayA_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h2d)) begin
										r_sub03_arrayA_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayA_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub03_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_arrayX_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub03_arrayX_addr <= $signed( r_run_k_29[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_arrayX_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub03_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub03_arrayX_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h2: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_arrayA_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h2c)) begin
										r_sub02_arrayA_addr <= $signed( r_run_copy35_i_67[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h2c)) begin
										r_sub02_arrayA_datain <= w_sys_tmp14;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_arrayA_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h2c)) begin
										r_sub02_arrayA_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayA_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub02_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_arrayX_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub02_arrayX_addr <= $signed( r_run_k_29[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_arrayX_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub02_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub02_arrayX_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'hb: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub11_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub11_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_arrayA_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h35)) begin
										r_sub11_arrayA_addr <= $signed( r_run_copy17_i_49[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h35)) begin
										r_sub11_arrayA_datain <= w_sys_tmp14;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_arrayA_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h35)) begin
										r_sub11_arrayA_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayA_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub11_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_arrayX_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub11_arrayX_addr <= $signed( r_run_k_29[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_arrayX_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub11_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub11_arrayX_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'he: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub14_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub14_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_arrayA_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h10) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h38)) begin
										r_sub14_arrayA_addr <= $signed( r_run_copy11_i_43[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h10) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h38)) begin
										r_sub14_arrayA_datain <= w_sys_tmp14;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_arrayA_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h10) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h38)) begin
										r_sub14_arrayA_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayA_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub14_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_arrayX_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub14_arrayX_addr <= $signed( r_run_k_29[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_arrayX_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub14_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub14_arrayX_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_arrayA_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h2b)) begin
										r_sub01_arrayA_addr <= $signed( r_run_copy37_i_69[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h2b)) begin
										r_sub01_arrayA_datain <= w_sys_tmp14;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_arrayA_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h2b)) begin
										r_sub01_arrayA_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayA_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub01_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_arrayX_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub01_arrayX_addr <= $signed( r_run_k_29[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_arrayX_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub01_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub01_arrayX_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'hd: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub13_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub13_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_arrayA_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hf) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h37)) begin
										r_sub13_arrayA_addr <= $signed( r_run_copy13_i_45[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hf) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h37)) begin
										r_sub13_arrayA_datain <= w_sys_tmp14;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_arrayA_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hf) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h37)) begin
										r_sub13_arrayA_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayA_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub13_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_arrayX_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub13_arrayX_addr <= $signed( r_run_k_29[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_arrayX_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub13_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub13_arrayX_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_arrayA_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h2a)) begin
										r_sub00_arrayA_addr <= $signed( r_run_i_27[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h2a)) begin
										r_sub00_arrayA_datain <= w_sys_tmp14;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_arrayA_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h2a)) begin
										r_sub00_arrayA_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayA_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub00_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_arrayX_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub00_arrayX_addr <= $signed( r_run_copy19_i_90[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_arrayX_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub00_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub00_arrayX_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub07_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub07_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_arrayA_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h31)) begin
										r_sub07_arrayA_addr <= $signed( r_run_copy25_i_57[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h31)) begin
										r_sub07_arrayA_datain <= w_sys_tmp14;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_arrayA_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h31)) begin
										r_sub07_arrayA_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayA_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub07_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_arrayX_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub07_arrayX_addr <= $signed( r_run_k_29[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_arrayX_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub07_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub07_arrayX_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h10: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub16_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub16_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_arrayA_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h12) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h3a)) begin
										r_sub16_arrayA_addr <= $signed( r_run_copy7_i_39[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h12) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h3a)) begin
										r_sub16_arrayA_datain <= w_sys_tmp14;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_arrayA_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h12) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h3a)) begin
										r_sub16_arrayA_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayA_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub16_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_arrayX_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub16_arrayX_addr <= $signed( r_run_k_29[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_arrayX_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub16_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub16_arrayX_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub06_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub06_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_arrayA_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h30)) begin
										r_sub06_arrayA_addr <= $signed( r_run_copy27_i_59[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h30)) begin
										r_sub06_arrayA_datain <= w_sys_tmp14;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_arrayA_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h30)) begin
										r_sub06_arrayA_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayA_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub06_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_arrayX_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub06_arrayX_addr <= $signed( r_run_k_29[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_arrayX_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub06_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub06_arrayX_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub15_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub15_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_arrayA_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h11) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h39)) begin
										r_sub15_arrayA_addr <= $signed( r_run_copy9_i_41[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h11) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h39)) begin
										r_sub15_arrayA_datain <= w_sys_tmp14;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_arrayA_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h11) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h39)) begin
										r_sub15_arrayA_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayA_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub15_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_arrayX_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub15_arrayX_addr <= $signed( r_run_k_29[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_arrayX_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub15_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub15_arrayX_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub05_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub05_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_arrayA_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h2f)) begin
										r_sub05_arrayA_addr <= $signed( r_run_copy29_i_61[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h2f)) begin
										r_sub05_arrayA_datain <= w_sys_tmp14;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_arrayA_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h2f)) begin
										r_sub05_arrayA_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayA_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub05_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_arrayX_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub05_arrayX_addr <= $signed( r_run_k_29[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_arrayX_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub05_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub05_arrayX_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h12: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub18_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub18_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_arrayA_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h14) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h3c)) begin
										r_sub18_arrayA_addr <= $signed( r_run_copy3_i_35[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h14) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h3c)) begin
										r_sub18_arrayA_datain <= w_sys_tmp14;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_arrayA_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h14) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h3c)) begin
										r_sub18_arrayA_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayA_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub18_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_arrayX_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub18_arrayX_addr <= $signed( r_run_k_29[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_arrayX_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub18_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub18_arrayX_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub04_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub04_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_arrayA_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h2e)) begin
										r_sub04_arrayA_addr <= $signed( r_run_copy31_i_63[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h2e)) begin
										r_sub04_arrayA_datain <= w_sys_tmp14;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_arrayA_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h2e)) begin
										r_sub04_arrayA_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayA_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub04_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_arrayX_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub04_arrayX_addr <= $signed( r_run_k_29[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_arrayX_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub04_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub04_arrayX_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h11: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub17_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub17_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_arrayA_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h13) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h3b)) begin
										r_sub17_arrayA_addr <= $signed( r_run_copy5_i_37[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h13) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h3b)) begin
										r_sub17_arrayA_datain <= w_sys_tmp14;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_arrayA_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h13) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h3b)) begin
										r_sub17_arrayA_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayA_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub17_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_arrayX_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub17_arrayX_addr <= $signed( r_run_k_29[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_arrayX_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub17_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub17_arrayX_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'ha: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub10_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub10_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_arrayA_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hc) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h34)) begin
										r_sub10_arrayA_addr <= $signed( r_run_copy19_i_51[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hc) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h34)) begin
										r_sub10_arrayA_datain <= w_sys_tmp14;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_arrayA_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hc) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h34)) begin
										r_sub10_arrayA_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayA_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub10_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_arrayX_addr <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub10_arrayX_addr <= $signed( r_run_k_29[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_arrayX_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayX_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub10_arrayX_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin
							r_sub10_arrayX_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4)) begin
										r_sys_tmp0_float <= w_sub00_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4)) begin
										r_sys_tmp1_float <= w_sub01_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4)) begin
										r_sys_tmp2_float <= w_sub05_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4)) begin
										r_sys_tmp3_float <= w_sub04_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4)) begin
										r_sys_tmp4_float <= w_sub03_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4)) begin
										r_sys_tmp5_float <= w_sub08_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4)) begin
										r_sys_tmp6_float <= w_sub13_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4)) begin
										r_sys_tmp7_float <= w_sub12_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4)) begin
										r_sys_tmp8_float <= w_sub11_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4)) begin
										r_sys_tmp9_float <= w_sub10_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4)) begin
										r_sys_tmp10_float <= w_sub09_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4)) begin
										r_sys_tmp11_float <= w_sub07_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4)) begin
										r_sys_tmp12_float <= w_sub06_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4)) begin
										r_sys_tmp13_float <= w_sub16_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4)) begin
										r_sys_tmp14_float <= w_sub19_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4)) begin
										r_sys_tmp15_float <= w_sub18_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4)) begin
										r_sys_tmp16_float <= w_sub17_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4)) begin
										r_sys_tmp17_float <= w_sub15_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4)) begin
										r_sys_tmp18_float <= w_sub14_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp19_float <= w_sub00_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp20_float <= w_sub02_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp21_float <= w_sub04_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp22_float <= w_sub06_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp23_float <= w_sub05_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp24_float <= w_sub03_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp25_float <= w_sub08_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp26_float <= w_sub12_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp27_float <= w_sub16_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp28_float <= w_sub19_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp29_float <= w_sub18_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp30_float <= w_sub17_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp31_float <= w_sub15_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp32_float <= w_sub14_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp33_float <= w_sub13_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp34_float <= w_sub11_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp35_float <= w_sub10_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp36_float <= w_sub09_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp37_float <= w_sub07_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp38_float <= w_sub04_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp39_float <= w_sub06_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp40_float <= w_sub08_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp41_float <= w_sub10_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp42_float <= w_sub12_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp43_float <= w_sub14_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp44_float <= w_sub16_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp45_float <= w_sub18_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp46_float <= w_sub19_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp47_float <= w_sub17_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp48_float <= w_sub15_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp49_float <= w_sub13_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp50_float <= w_sub11_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp51_float <= w_sub09_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp52_float <= w_sub07_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp53_float <= w_sub05_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp54_float <= w_sub03_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h3)) begin
										r_sys_tmp55_float <= w_sub01_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h4)) begin
										r_sys_tmp56_float <= w_sub02_arrayX_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
