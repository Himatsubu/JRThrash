/*
TimeStamp:	2016/5/25		7:17
*/


module P3_2dim(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy	
);

	reg  signed [31:0] r_ip_DivInt_dividend_0;
	reg  signed [31:0] r_ip_DivInt_divisor_0;
	wire signed [31:0] w_ip_DivInt_quotient_0;
	wire signed [31:0] w_ip_DivInt_fractional_0;
	reg  signed [31:0] r_ip_DivInt_dividend_1;
	reg  signed [31:0] r_ip_DivInt_divisor_1;
	wire signed [31:0] w_ip_DivInt_quotient_1;
	wire signed [31:0] w_ip_DivInt_fractional_1;
	reg         [31:0] r_ip_AddFloat_portA_0;
	reg         [31:0] r_ip_AddFloat_portB_0;
	wire        [31:0] w_ip_AddFloat_result_0;
	reg         [31:0] r_ip_MultFloat_multiplicand_0;
	reg         [31:0] r_ip_MultFloat_multiplier_0;
	wire        [31:0] w_ip_MultFloat_product_0;
	reg  signed [31:0] r_ip_FixedToFloat_fixed_0;
	wire        [31:0] w_ip_FixedToFloat_floating_0;
	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 6:0] r_sys_run_phase;
	reg         [ 4:0] r_sys_run_stage;
	reg         [ 7:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 4:0] w_sys_run_stage_p1;
	wire        [ 7:0] w_sys_run_step_p1;
	wire signed [ 9:0] w_fld_T_0_addr_0;
	wire        [31:0] w_fld_T_0_datain_0;
	wire        [31:0] w_fld_T_0_dataout_0;
	wire               w_fld_T_0_r_w_0;
	wire               w_fld_T_0_ce_0;
	reg  signed [ 9:0] r_fld_T_0_addr_1;
	reg         [31:0] r_fld_T_0_datain_1;
	wire        [31:0] w_fld_T_0_dataout_1;
	reg                r_fld_T_0_r_w_1;
	wire               w_fld_T_0_ce_1;
	wire signed [ 9:0] w_fld_TT_1_addr_0;
	wire        [31:0] w_fld_TT_1_datain_0;
	wire        [31:0] w_fld_TT_1_dataout_0;
	wire               w_fld_TT_1_r_w_0;
	wire               w_fld_TT_1_ce_0;
	reg  signed [ 9:0] r_fld_TT_1_addr_1;
	reg         [31:0] r_fld_TT_1_datain_1;
	wire        [31:0] w_fld_TT_1_dataout_1;
	reg                r_fld_TT_1_r_w_1;
	wire               w_fld_TT_1_ce_1;
	wire signed [ 9:0] w_fld_U_2_addr_0;
	wire        [31:0] w_fld_U_2_datain_0;
	wire        [31:0] w_fld_U_2_dataout_0;
	wire               w_fld_U_2_r_w_0;
	wire               w_fld_U_2_ce_0;
	reg  signed [ 9:0] r_fld_U_2_addr_1;
	reg         [31:0] r_fld_U_2_datain_1;
	wire        [31:0] w_fld_U_2_dataout_1;
	reg                r_fld_U_2_r_w_1;
	wire               w_fld_U_2_ce_1;
	wire signed [ 9:0] w_fld_V_3_addr_0;
	wire        [31:0] w_fld_V_3_datain_0;
	wire        [31:0] w_fld_V_3_dataout_0;
	wire               w_fld_V_3_r_w_0;
	wire               w_fld_V_3_ce_0;
	reg  signed [ 9:0] r_fld_V_3_addr_1;
	reg         [31:0] r_fld_V_3_datain_1;
	wire        [31:0] w_fld_V_3_dataout_1;
	reg                r_fld_V_3_r_w_1;
	wire               w_fld_V_3_ce_1;
	reg  signed [31:0] r_run_k_29;
	reg  signed [31:0] r_run_j_30;
	reg  signed [31:0] r_run_n_31;
	reg  signed [31:0] r_run_mx_32;
	reg  signed [31:0] r_run_my_33;
	reg         [31:0] r_run_dt_34;
	reg         [31:0] r_run_dx_35;
	reg         [31:0] r_run_dy_36;
	reg         [31:0] r_run_r1_37;
	reg         [31:0] r_run_r2_38;
	reg         [31:0] r_run_r3_39;
	reg         [31:0] r_run_r4_40;
	reg         [31:0] r_run_YY_41;
	reg  signed [31:0] r_run_kx_42;
	reg  signed [31:0] r_run_ky_43;
	reg  signed [31:0] r_run_nlast_44;
	reg  signed [31:0] r_run_copy0_j_45;
	reg  signed [31:0] r_run_copy1_j_46;
	reg  signed [31:0] r_run_copy2_j_47;
	reg  signed [31:0] r_run_copy0_j_48;
	reg                r_sub19_run_req;
	wire               w_sub19_run_busy;
	wire signed [ 9:0] w_sub19_T_addr;
	reg  signed [ 9:0] r_sub19_T_addr;
	wire        [31:0] w_sub19_T_datain;
	reg         [31:0] r_sub19_T_datain;
	wire        [31:0] w_sub19_T_dataout;
	wire               w_sub19_T_r_w;
	reg                r_sub19_T_r_w;
	wire signed [ 9:0] w_sub19_V_addr;
	reg  signed [ 9:0] r_sub19_V_addr;
	wire        [31:0] w_sub19_V_datain;
	reg         [31:0] r_sub19_V_datain;
	wire        [31:0] w_sub19_V_dataout;
	wire               w_sub19_V_r_w;
	reg                r_sub19_V_r_w;
	wire signed [ 9:0] w_sub19_U_addr;
	reg  signed [ 9:0] r_sub19_U_addr;
	wire        [31:0] w_sub19_U_datain;
	reg         [31:0] r_sub19_U_datain;
	wire        [31:0] w_sub19_U_dataout;
	wire               w_sub19_U_r_w;
	reg                r_sub19_U_r_w;
	wire signed [ 9:0] w_sub19_result_addr;
	reg  signed [ 9:0] r_sub19_result_addr;
	wire        [31:0] w_sub19_result_datain;
	reg         [31:0] r_sub19_result_datain;
	wire        [31:0] w_sub19_result_dataout;
	wire               w_sub19_result_r_w;
	reg                r_sub19_result_r_w;
	reg                r_sub09_run_req;
	wire               w_sub09_run_busy;
	wire signed [ 9:0] w_sub09_T_addr;
	reg  signed [ 9:0] r_sub09_T_addr;
	wire        [31:0] w_sub09_T_datain;
	reg         [31:0] r_sub09_T_datain;
	wire        [31:0] w_sub09_T_dataout;
	wire               w_sub09_T_r_w;
	reg                r_sub09_T_r_w;
	wire signed [ 9:0] w_sub09_V_addr;
	reg  signed [ 9:0] r_sub09_V_addr;
	wire        [31:0] w_sub09_V_datain;
	reg         [31:0] r_sub09_V_datain;
	wire        [31:0] w_sub09_V_dataout;
	wire               w_sub09_V_r_w;
	reg                r_sub09_V_r_w;
	wire signed [ 9:0] w_sub09_U_addr;
	reg  signed [ 9:0] r_sub09_U_addr;
	wire        [31:0] w_sub09_U_datain;
	reg         [31:0] r_sub09_U_datain;
	wire        [31:0] w_sub09_U_dataout;
	wire               w_sub09_U_r_w;
	reg                r_sub09_U_r_w;
	wire signed [ 9:0] w_sub09_result_addr;
	reg  signed [ 9:0] r_sub09_result_addr;
	wire        [31:0] w_sub09_result_datain;
	reg         [31:0] r_sub09_result_datain;
	wire        [31:0] w_sub09_result_dataout;
	wire               w_sub09_result_r_w;
	reg                r_sub09_result_r_w;
	reg                r_sub08_run_req;
	wire               w_sub08_run_busy;
	wire signed [ 9:0] w_sub08_T_addr;
	reg  signed [ 9:0] r_sub08_T_addr;
	wire        [31:0] w_sub08_T_datain;
	reg         [31:0] r_sub08_T_datain;
	wire        [31:0] w_sub08_T_dataout;
	wire               w_sub08_T_r_w;
	reg                r_sub08_T_r_w;
	wire signed [ 9:0] w_sub08_V_addr;
	reg  signed [ 9:0] r_sub08_V_addr;
	wire        [31:0] w_sub08_V_datain;
	reg         [31:0] r_sub08_V_datain;
	wire        [31:0] w_sub08_V_dataout;
	wire               w_sub08_V_r_w;
	reg                r_sub08_V_r_w;
	wire signed [ 9:0] w_sub08_U_addr;
	reg  signed [ 9:0] r_sub08_U_addr;
	wire        [31:0] w_sub08_U_datain;
	reg         [31:0] r_sub08_U_datain;
	wire        [31:0] w_sub08_U_dataout;
	wire               w_sub08_U_r_w;
	reg                r_sub08_U_r_w;
	wire signed [ 9:0] w_sub08_result_addr;
	reg  signed [ 9:0] r_sub08_result_addr;
	wire        [31:0] w_sub08_result_datain;
	reg         [31:0] r_sub08_result_datain;
	wire        [31:0] w_sub08_result_dataout;
	wire               w_sub08_result_r_w;
	reg                r_sub08_result_r_w;
	reg                r_sub24_run_req;
	wire               w_sub24_run_busy;
	wire signed [ 9:0] w_sub24_T_addr;
	reg  signed [ 9:0] r_sub24_T_addr;
	wire        [31:0] w_sub24_T_datain;
	reg         [31:0] r_sub24_T_datain;
	wire        [31:0] w_sub24_T_dataout;
	wire               w_sub24_T_r_w;
	reg                r_sub24_T_r_w;
	wire signed [ 9:0] w_sub24_V_addr;
	reg  signed [ 9:0] r_sub24_V_addr;
	wire        [31:0] w_sub24_V_datain;
	reg         [31:0] r_sub24_V_datain;
	wire        [31:0] w_sub24_V_dataout;
	wire               w_sub24_V_r_w;
	reg                r_sub24_V_r_w;
	wire signed [ 9:0] w_sub24_U_addr;
	reg  signed [ 9:0] r_sub24_U_addr;
	wire        [31:0] w_sub24_U_datain;
	reg         [31:0] r_sub24_U_datain;
	wire        [31:0] w_sub24_U_dataout;
	wire               w_sub24_U_r_w;
	reg                r_sub24_U_r_w;
	wire signed [ 9:0] w_sub24_result_addr;
	reg  signed [ 9:0] r_sub24_result_addr;
	wire        [31:0] w_sub24_result_datain;
	reg         [31:0] r_sub24_result_datain;
	wire        [31:0] w_sub24_result_dataout;
	wire               w_sub24_result_r_w;
	reg                r_sub24_result_r_w;
	reg                r_sub22_run_req;
	wire               w_sub22_run_busy;
	wire signed [ 9:0] w_sub22_T_addr;
	reg  signed [ 9:0] r_sub22_T_addr;
	wire        [31:0] w_sub22_T_datain;
	reg         [31:0] r_sub22_T_datain;
	wire        [31:0] w_sub22_T_dataout;
	wire               w_sub22_T_r_w;
	reg                r_sub22_T_r_w;
	wire signed [ 9:0] w_sub22_V_addr;
	reg  signed [ 9:0] r_sub22_V_addr;
	wire        [31:0] w_sub22_V_datain;
	reg         [31:0] r_sub22_V_datain;
	wire        [31:0] w_sub22_V_dataout;
	wire               w_sub22_V_r_w;
	reg                r_sub22_V_r_w;
	wire signed [ 9:0] w_sub22_U_addr;
	reg  signed [ 9:0] r_sub22_U_addr;
	wire        [31:0] w_sub22_U_datain;
	reg         [31:0] r_sub22_U_datain;
	wire        [31:0] w_sub22_U_dataout;
	wire               w_sub22_U_r_w;
	reg                r_sub22_U_r_w;
	wire signed [ 9:0] w_sub22_result_addr;
	reg  signed [ 9:0] r_sub22_result_addr;
	wire        [31:0] w_sub22_result_datain;
	reg         [31:0] r_sub22_result_datain;
	wire        [31:0] w_sub22_result_dataout;
	wire               w_sub22_result_r_w;
	reg                r_sub22_result_r_w;
	reg                r_sub23_run_req;
	wire               w_sub23_run_busy;
	wire signed [ 9:0] w_sub23_T_addr;
	reg  signed [ 9:0] r_sub23_T_addr;
	wire        [31:0] w_sub23_T_datain;
	reg         [31:0] r_sub23_T_datain;
	wire        [31:0] w_sub23_T_dataout;
	wire               w_sub23_T_r_w;
	reg                r_sub23_T_r_w;
	wire signed [ 9:0] w_sub23_V_addr;
	reg  signed [ 9:0] r_sub23_V_addr;
	wire        [31:0] w_sub23_V_datain;
	reg         [31:0] r_sub23_V_datain;
	wire        [31:0] w_sub23_V_dataout;
	wire               w_sub23_V_r_w;
	reg                r_sub23_V_r_w;
	wire signed [ 9:0] w_sub23_U_addr;
	reg  signed [ 9:0] r_sub23_U_addr;
	wire        [31:0] w_sub23_U_datain;
	reg         [31:0] r_sub23_U_datain;
	wire        [31:0] w_sub23_U_dataout;
	wire               w_sub23_U_r_w;
	reg                r_sub23_U_r_w;
	wire signed [ 9:0] w_sub23_result_addr;
	reg  signed [ 9:0] r_sub23_result_addr;
	wire        [31:0] w_sub23_result_datain;
	reg         [31:0] r_sub23_result_datain;
	wire        [31:0] w_sub23_result_dataout;
	wire               w_sub23_result_r_w;
	reg                r_sub23_result_r_w;
	reg                r_sub12_run_req;
	wire               w_sub12_run_busy;
	wire signed [ 9:0] w_sub12_T_addr;
	reg  signed [ 9:0] r_sub12_T_addr;
	wire        [31:0] w_sub12_T_datain;
	reg         [31:0] r_sub12_T_datain;
	wire        [31:0] w_sub12_T_dataout;
	wire               w_sub12_T_r_w;
	reg                r_sub12_T_r_w;
	wire signed [ 9:0] w_sub12_V_addr;
	reg  signed [ 9:0] r_sub12_V_addr;
	wire        [31:0] w_sub12_V_datain;
	reg         [31:0] r_sub12_V_datain;
	wire        [31:0] w_sub12_V_dataout;
	wire               w_sub12_V_r_w;
	reg                r_sub12_V_r_w;
	wire signed [ 9:0] w_sub12_U_addr;
	reg  signed [ 9:0] r_sub12_U_addr;
	wire        [31:0] w_sub12_U_datain;
	reg         [31:0] r_sub12_U_datain;
	wire        [31:0] w_sub12_U_dataout;
	wire               w_sub12_U_r_w;
	reg                r_sub12_U_r_w;
	wire signed [ 9:0] w_sub12_result_addr;
	reg  signed [ 9:0] r_sub12_result_addr;
	wire        [31:0] w_sub12_result_datain;
	reg         [31:0] r_sub12_result_datain;
	wire        [31:0] w_sub12_result_dataout;
	wire               w_sub12_result_r_w;
	reg                r_sub12_result_r_w;
	reg                r_sub03_run_req;
	wire               w_sub03_run_busy;
	wire signed [ 9:0] w_sub03_T_addr;
	reg  signed [ 9:0] r_sub03_T_addr;
	wire        [31:0] w_sub03_T_datain;
	reg         [31:0] r_sub03_T_datain;
	wire        [31:0] w_sub03_T_dataout;
	wire               w_sub03_T_r_w;
	reg                r_sub03_T_r_w;
	wire signed [ 9:0] w_sub03_V_addr;
	reg  signed [ 9:0] r_sub03_V_addr;
	wire        [31:0] w_sub03_V_datain;
	reg         [31:0] r_sub03_V_datain;
	wire        [31:0] w_sub03_V_dataout;
	wire               w_sub03_V_r_w;
	reg                r_sub03_V_r_w;
	wire signed [ 9:0] w_sub03_U_addr;
	reg  signed [ 9:0] r_sub03_U_addr;
	wire        [31:0] w_sub03_U_datain;
	reg         [31:0] r_sub03_U_datain;
	wire        [31:0] w_sub03_U_dataout;
	wire               w_sub03_U_r_w;
	reg                r_sub03_U_r_w;
	wire signed [ 9:0] w_sub03_result_addr;
	reg  signed [ 9:0] r_sub03_result_addr;
	wire        [31:0] w_sub03_result_datain;
	reg         [31:0] r_sub03_result_datain;
	wire        [31:0] w_sub03_result_dataout;
	wire               w_sub03_result_r_w;
	reg                r_sub03_result_r_w;
	reg                r_sub02_run_req;
	wire               w_sub02_run_busy;
	wire signed [ 9:0] w_sub02_T_addr;
	reg  signed [ 9:0] r_sub02_T_addr;
	wire        [31:0] w_sub02_T_datain;
	reg         [31:0] r_sub02_T_datain;
	wire        [31:0] w_sub02_T_dataout;
	wire               w_sub02_T_r_w;
	reg                r_sub02_T_r_w;
	wire signed [ 9:0] w_sub02_V_addr;
	reg  signed [ 9:0] r_sub02_V_addr;
	wire        [31:0] w_sub02_V_datain;
	reg         [31:0] r_sub02_V_datain;
	wire        [31:0] w_sub02_V_dataout;
	wire               w_sub02_V_r_w;
	reg                r_sub02_V_r_w;
	wire signed [ 9:0] w_sub02_U_addr;
	reg  signed [ 9:0] r_sub02_U_addr;
	wire        [31:0] w_sub02_U_datain;
	reg         [31:0] r_sub02_U_datain;
	wire        [31:0] w_sub02_U_dataout;
	wire               w_sub02_U_r_w;
	reg                r_sub02_U_r_w;
	wire signed [ 9:0] w_sub02_result_addr;
	reg  signed [ 9:0] r_sub02_result_addr;
	wire        [31:0] w_sub02_result_datain;
	reg         [31:0] r_sub02_result_datain;
	wire        [31:0] w_sub02_result_dataout;
	wire               w_sub02_result_r_w;
	reg                r_sub02_result_r_w;
	reg                r_sub11_run_req;
	wire               w_sub11_run_busy;
	wire signed [ 9:0] w_sub11_T_addr;
	reg  signed [ 9:0] r_sub11_T_addr;
	wire        [31:0] w_sub11_T_datain;
	reg         [31:0] r_sub11_T_datain;
	wire        [31:0] w_sub11_T_dataout;
	wire               w_sub11_T_r_w;
	reg                r_sub11_T_r_w;
	wire signed [ 9:0] w_sub11_V_addr;
	reg  signed [ 9:0] r_sub11_V_addr;
	wire        [31:0] w_sub11_V_datain;
	reg         [31:0] r_sub11_V_datain;
	wire        [31:0] w_sub11_V_dataout;
	wire               w_sub11_V_r_w;
	reg                r_sub11_V_r_w;
	wire signed [ 9:0] w_sub11_U_addr;
	reg  signed [ 9:0] r_sub11_U_addr;
	wire        [31:0] w_sub11_U_datain;
	reg         [31:0] r_sub11_U_datain;
	wire        [31:0] w_sub11_U_dataout;
	wire               w_sub11_U_r_w;
	reg                r_sub11_U_r_w;
	wire signed [ 9:0] w_sub11_result_addr;
	reg  signed [ 9:0] r_sub11_result_addr;
	wire        [31:0] w_sub11_result_datain;
	reg         [31:0] r_sub11_result_datain;
	wire        [31:0] w_sub11_result_dataout;
	wire               w_sub11_result_r_w;
	reg                r_sub11_result_r_w;
	reg                r_sub14_run_req;
	wire               w_sub14_run_busy;
	wire signed [ 9:0] w_sub14_T_addr;
	reg  signed [ 9:0] r_sub14_T_addr;
	wire        [31:0] w_sub14_T_datain;
	reg         [31:0] r_sub14_T_datain;
	wire        [31:0] w_sub14_T_dataout;
	wire               w_sub14_T_r_w;
	reg                r_sub14_T_r_w;
	wire signed [ 9:0] w_sub14_V_addr;
	reg  signed [ 9:0] r_sub14_V_addr;
	wire        [31:0] w_sub14_V_datain;
	reg         [31:0] r_sub14_V_datain;
	wire        [31:0] w_sub14_V_dataout;
	wire               w_sub14_V_r_w;
	reg                r_sub14_V_r_w;
	wire signed [ 9:0] w_sub14_U_addr;
	reg  signed [ 9:0] r_sub14_U_addr;
	wire        [31:0] w_sub14_U_datain;
	reg         [31:0] r_sub14_U_datain;
	wire        [31:0] w_sub14_U_dataout;
	wire               w_sub14_U_r_w;
	reg                r_sub14_U_r_w;
	wire signed [ 9:0] w_sub14_result_addr;
	reg  signed [ 9:0] r_sub14_result_addr;
	wire        [31:0] w_sub14_result_datain;
	reg         [31:0] r_sub14_result_datain;
	wire        [31:0] w_sub14_result_dataout;
	wire               w_sub14_result_r_w;
	reg                r_sub14_result_r_w;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [ 9:0] w_sub01_T_addr;
	reg  signed [ 9:0] r_sub01_T_addr;
	wire        [31:0] w_sub01_T_datain;
	reg         [31:0] r_sub01_T_datain;
	wire        [31:0] w_sub01_T_dataout;
	wire               w_sub01_T_r_w;
	reg                r_sub01_T_r_w;
	wire signed [ 9:0] w_sub01_V_addr;
	reg  signed [ 9:0] r_sub01_V_addr;
	wire        [31:0] w_sub01_V_datain;
	reg         [31:0] r_sub01_V_datain;
	wire        [31:0] w_sub01_V_dataout;
	wire               w_sub01_V_r_w;
	reg                r_sub01_V_r_w;
	wire signed [ 9:0] w_sub01_U_addr;
	reg  signed [ 9:0] r_sub01_U_addr;
	wire        [31:0] w_sub01_U_datain;
	reg         [31:0] r_sub01_U_datain;
	wire        [31:0] w_sub01_U_dataout;
	wire               w_sub01_U_r_w;
	reg                r_sub01_U_r_w;
	wire signed [ 9:0] w_sub01_result_addr;
	reg  signed [ 9:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [ 9:0] w_sub00_T_addr;
	reg  signed [ 9:0] r_sub00_T_addr;
	wire        [31:0] w_sub00_T_datain;
	reg         [31:0] r_sub00_T_datain;
	wire        [31:0] w_sub00_T_dataout;
	wire               w_sub00_T_r_w;
	reg                r_sub00_T_r_w;
	wire signed [ 9:0] w_sub00_V_addr;
	reg  signed [ 9:0] r_sub00_V_addr;
	wire        [31:0] w_sub00_V_datain;
	reg         [31:0] r_sub00_V_datain;
	wire        [31:0] w_sub00_V_dataout;
	wire               w_sub00_V_r_w;
	reg                r_sub00_V_r_w;
	wire signed [ 9:0] w_sub00_U_addr;
	reg  signed [ 9:0] r_sub00_U_addr;
	wire        [31:0] w_sub00_U_datain;
	reg         [31:0] r_sub00_U_datain;
	wire        [31:0] w_sub00_U_dataout;
	wire               w_sub00_U_r_w;
	reg                r_sub00_U_r_w;
	wire signed [ 9:0] w_sub00_result_addr;
	reg  signed [ 9:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	reg                r_sub13_run_req;
	wire               w_sub13_run_busy;
	wire signed [ 9:0] w_sub13_T_addr;
	reg  signed [ 9:0] r_sub13_T_addr;
	wire        [31:0] w_sub13_T_datain;
	reg         [31:0] r_sub13_T_datain;
	wire        [31:0] w_sub13_T_dataout;
	wire               w_sub13_T_r_w;
	reg                r_sub13_T_r_w;
	wire signed [ 9:0] w_sub13_V_addr;
	reg  signed [ 9:0] r_sub13_V_addr;
	wire        [31:0] w_sub13_V_datain;
	reg         [31:0] r_sub13_V_datain;
	wire        [31:0] w_sub13_V_dataout;
	wire               w_sub13_V_r_w;
	reg                r_sub13_V_r_w;
	wire signed [ 9:0] w_sub13_U_addr;
	reg  signed [ 9:0] r_sub13_U_addr;
	wire        [31:0] w_sub13_U_datain;
	reg         [31:0] r_sub13_U_datain;
	wire        [31:0] w_sub13_U_dataout;
	wire               w_sub13_U_r_w;
	reg                r_sub13_U_r_w;
	wire signed [ 9:0] w_sub13_result_addr;
	reg  signed [ 9:0] r_sub13_result_addr;
	wire        [31:0] w_sub13_result_datain;
	reg         [31:0] r_sub13_result_datain;
	wire        [31:0] w_sub13_result_dataout;
	wire               w_sub13_result_r_w;
	reg                r_sub13_result_r_w;
	reg                r_sub07_run_req;
	wire               w_sub07_run_busy;
	wire signed [ 9:0] w_sub07_T_addr;
	reg  signed [ 9:0] r_sub07_T_addr;
	wire        [31:0] w_sub07_T_datain;
	reg         [31:0] r_sub07_T_datain;
	wire        [31:0] w_sub07_T_dataout;
	wire               w_sub07_T_r_w;
	reg                r_sub07_T_r_w;
	wire signed [ 9:0] w_sub07_V_addr;
	reg  signed [ 9:0] r_sub07_V_addr;
	wire        [31:0] w_sub07_V_datain;
	reg         [31:0] r_sub07_V_datain;
	wire        [31:0] w_sub07_V_dataout;
	wire               w_sub07_V_r_w;
	reg                r_sub07_V_r_w;
	wire signed [ 9:0] w_sub07_U_addr;
	reg  signed [ 9:0] r_sub07_U_addr;
	wire        [31:0] w_sub07_U_datain;
	reg         [31:0] r_sub07_U_datain;
	wire        [31:0] w_sub07_U_dataout;
	wire               w_sub07_U_r_w;
	reg                r_sub07_U_r_w;
	wire signed [ 9:0] w_sub07_result_addr;
	reg  signed [ 9:0] r_sub07_result_addr;
	wire        [31:0] w_sub07_result_datain;
	reg         [31:0] r_sub07_result_datain;
	wire        [31:0] w_sub07_result_dataout;
	wire               w_sub07_result_r_w;
	reg                r_sub07_result_r_w;
	reg                r_sub16_run_req;
	wire               w_sub16_run_busy;
	wire signed [ 9:0] w_sub16_T_addr;
	reg  signed [ 9:0] r_sub16_T_addr;
	wire        [31:0] w_sub16_T_datain;
	reg         [31:0] r_sub16_T_datain;
	wire        [31:0] w_sub16_T_dataout;
	wire               w_sub16_T_r_w;
	reg                r_sub16_T_r_w;
	wire signed [ 9:0] w_sub16_V_addr;
	reg  signed [ 9:0] r_sub16_V_addr;
	wire        [31:0] w_sub16_V_datain;
	reg         [31:0] r_sub16_V_datain;
	wire        [31:0] w_sub16_V_dataout;
	wire               w_sub16_V_r_w;
	reg                r_sub16_V_r_w;
	wire signed [ 9:0] w_sub16_U_addr;
	reg  signed [ 9:0] r_sub16_U_addr;
	wire        [31:0] w_sub16_U_datain;
	reg         [31:0] r_sub16_U_datain;
	wire        [31:0] w_sub16_U_dataout;
	wire               w_sub16_U_r_w;
	reg                r_sub16_U_r_w;
	wire signed [ 9:0] w_sub16_result_addr;
	reg  signed [ 9:0] r_sub16_result_addr;
	wire        [31:0] w_sub16_result_datain;
	reg         [31:0] r_sub16_result_datain;
	wire        [31:0] w_sub16_result_dataout;
	wire               w_sub16_result_r_w;
	reg                r_sub16_result_r_w;
	reg                r_sub06_run_req;
	wire               w_sub06_run_busy;
	wire signed [ 9:0] w_sub06_T_addr;
	reg  signed [ 9:0] r_sub06_T_addr;
	wire        [31:0] w_sub06_T_datain;
	reg         [31:0] r_sub06_T_datain;
	wire        [31:0] w_sub06_T_dataout;
	wire               w_sub06_T_r_w;
	reg                r_sub06_T_r_w;
	wire signed [ 9:0] w_sub06_V_addr;
	reg  signed [ 9:0] r_sub06_V_addr;
	wire        [31:0] w_sub06_V_datain;
	reg         [31:0] r_sub06_V_datain;
	wire        [31:0] w_sub06_V_dataout;
	wire               w_sub06_V_r_w;
	reg                r_sub06_V_r_w;
	wire signed [ 9:0] w_sub06_U_addr;
	reg  signed [ 9:0] r_sub06_U_addr;
	wire        [31:0] w_sub06_U_datain;
	reg         [31:0] r_sub06_U_datain;
	wire        [31:0] w_sub06_U_dataout;
	wire               w_sub06_U_r_w;
	reg                r_sub06_U_r_w;
	wire signed [ 9:0] w_sub06_result_addr;
	reg  signed [ 9:0] r_sub06_result_addr;
	wire        [31:0] w_sub06_result_datain;
	reg         [31:0] r_sub06_result_datain;
	wire        [31:0] w_sub06_result_dataout;
	wire               w_sub06_result_r_w;
	reg                r_sub06_result_r_w;
	reg                r_sub15_run_req;
	wire               w_sub15_run_busy;
	wire signed [ 9:0] w_sub15_T_addr;
	reg  signed [ 9:0] r_sub15_T_addr;
	wire        [31:0] w_sub15_T_datain;
	reg         [31:0] r_sub15_T_datain;
	wire        [31:0] w_sub15_T_dataout;
	wire               w_sub15_T_r_w;
	reg                r_sub15_T_r_w;
	wire signed [ 9:0] w_sub15_V_addr;
	reg  signed [ 9:0] r_sub15_V_addr;
	wire        [31:0] w_sub15_V_datain;
	reg         [31:0] r_sub15_V_datain;
	wire        [31:0] w_sub15_V_dataout;
	wire               w_sub15_V_r_w;
	reg                r_sub15_V_r_w;
	wire signed [ 9:0] w_sub15_U_addr;
	reg  signed [ 9:0] r_sub15_U_addr;
	wire        [31:0] w_sub15_U_datain;
	reg         [31:0] r_sub15_U_datain;
	wire        [31:0] w_sub15_U_dataout;
	wire               w_sub15_U_r_w;
	reg                r_sub15_U_r_w;
	wire signed [ 9:0] w_sub15_result_addr;
	reg  signed [ 9:0] r_sub15_result_addr;
	wire        [31:0] w_sub15_result_datain;
	reg         [31:0] r_sub15_result_datain;
	wire        [31:0] w_sub15_result_dataout;
	wire               w_sub15_result_r_w;
	reg                r_sub15_result_r_w;
	reg                r_sub05_run_req;
	wire               w_sub05_run_busy;
	wire signed [ 9:0] w_sub05_T_addr;
	reg  signed [ 9:0] r_sub05_T_addr;
	wire        [31:0] w_sub05_T_datain;
	reg         [31:0] r_sub05_T_datain;
	wire        [31:0] w_sub05_T_dataout;
	wire               w_sub05_T_r_w;
	reg                r_sub05_T_r_w;
	wire signed [ 9:0] w_sub05_V_addr;
	reg  signed [ 9:0] r_sub05_V_addr;
	wire        [31:0] w_sub05_V_datain;
	reg         [31:0] r_sub05_V_datain;
	wire        [31:0] w_sub05_V_dataout;
	wire               w_sub05_V_r_w;
	reg                r_sub05_V_r_w;
	wire signed [ 9:0] w_sub05_U_addr;
	reg  signed [ 9:0] r_sub05_U_addr;
	wire        [31:0] w_sub05_U_datain;
	reg         [31:0] r_sub05_U_datain;
	wire        [31:0] w_sub05_U_dataout;
	wire               w_sub05_U_r_w;
	reg                r_sub05_U_r_w;
	wire signed [ 9:0] w_sub05_result_addr;
	reg  signed [ 9:0] r_sub05_result_addr;
	wire        [31:0] w_sub05_result_datain;
	reg         [31:0] r_sub05_result_datain;
	wire        [31:0] w_sub05_result_dataout;
	wire               w_sub05_result_r_w;
	reg                r_sub05_result_r_w;
	reg                r_sub18_run_req;
	wire               w_sub18_run_busy;
	wire signed [ 9:0] w_sub18_T_addr;
	reg  signed [ 9:0] r_sub18_T_addr;
	wire        [31:0] w_sub18_T_datain;
	reg         [31:0] r_sub18_T_datain;
	wire        [31:0] w_sub18_T_dataout;
	wire               w_sub18_T_r_w;
	reg                r_sub18_T_r_w;
	wire signed [ 9:0] w_sub18_V_addr;
	reg  signed [ 9:0] r_sub18_V_addr;
	wire        [31:0] w_sub18_V_datain;
	reg         [31:0] r_sub18_V_datain;
	wire        [31:0] w_sub18_V_dataout;
	wire               w_sub18_V_r_w;
	reg                r_sub18_V_r_w;
	wire signed [ 9:0] w_sub18_U_addr;
	reg  signed [ 9:0] r_sub18_U_addr;
	wire        [31:0] w_sub18_U_datain;
	reg         [31:0] r_sub18_U_datain;
	wire        [31:0] w_sub18_U_dataout;
	wire               w_sub18_U_r_w;
	reg                r_sub18_U_r_w;
	wire signed [ 9:0] w_sub18_result_addr;
	reg  signed [ 9:0] r_sub18_result_addr;
	wire        [31:0] w_sub18_result_datain;
	reg         [31:0] r_sub18_result_datain;
	wire        [31:0] w_sub18_result_dataout;
	wire               w_sub18_result_r_w;
	reg                r_sub18_result_r_w;
	reg                r_sub04_run_req;
	wire               w_sub04_run_busy;
	wire signed [ 9:0] w_sub04_T_addr;
	reg  signed [ 9:0] r_sub04_T_addr;
	wire        [31:0] w_sub04_T_datain;
	reg         [31:0] r_sub04_T_datain;
	wire        [31:0] w_sub04_T_dataout;
	wire               w_sub04_T_r_w;
	reg                r_sub04_T_r_w;
	wire signed [ 9:0] w_sub04_V_addr;
	reg  signed [ 9:0] r_sub04_V_addr;
	wire        [31:0] w_sub04_V_datain;
	reg         [31:0] r_sub04_V_datain;
	wire        [31:0] w_sub04_V_dataout;
	wire               w_sub04_V_r_w;
	reg                r_sub04_V_r_w;
	wire signed [ 9:0] w_sub04_U_addr;
	reg  signed [ 9:0] r_sub04_U_addr;
	wire        [31:0] w_sub04_U_datain;
	reg         [31:0] r_sub04_U_datain;
	wire        [31:0] w_sub04_U_dataout;
	wire               w_sub04_U_r_w;
	reg                r_sub04_U_r_w;
	wire signed [ 9:0] w_sub04_result_addr;
	reg  signed [ 9:0] r_sub04_result_addr;
	wire        [31:0] w_sub04_result_datain;
	reg         [31:0] r_sub04_result_datain;
	wire        [31:0] w_sub04_result_dataout;
	wire               w_sub04_result_r_w;
	reg                r_sub04_result_r_w;
	reg                r_sub17_run_req;
	wire               w_sub17_run_busy;
	wire signed [ 9:0] w_sub17_T_addr;
	reg  signed [ 9:0] r_sub17_T_addr;
	wire        [31:0] w_sub17_T_datain;
	reg         [31:0] r_sub17_T_datain;
	wire        [31:0] w_sub17_T_dataout;
	wire               w_sub17_T_r_w;
	reg                r_sub17_T_r_w;
	wire signed [ 9:0] w_sub17_V_addr;
	reg  signed [ 9:0] r_sub17_V_addr;
	wire        [31:0] w_sub17_V_datain;
	reg         [31:0] r_sub17_V_datain;
	wire        [31:0] w_sub17_V_dataout;
	wire               w_sub17_V_r_w;
	reg                r_sub17_V_r_w;
	wire signed [ 9:0] w_sub17_U_addr;
	reg  signed [ 9:0] r_sub17_U_addr;
	wire        [31:0] w_sub17_U_datain;
	reg         [31:0] r_sub17_U_datain;
	wire        [31:0] w_sub17_U_dataout;
	wire               w_sub17_U_r_w;
	reg                r_sub17_U_r_w;
	wire signed [ 9:0] w_sub17_result_addr;
	reg  signed [ 9:0] r_sub17_result_addr;
	wire        [31:0] w_sub17_result_datain;
	reg         [31:0] r_sub17_result_datain;
	wire        [31:0] w_sub17_result_dataout;
	wire               w_sub17_result_r_w;
	reg                r_sub17_result_r_w;
	reg                r_sub10_run_req;
	wire               w_sub10_run_busy;
	wire signed [ 9:0] w_sub10_T_addr;
	reg  signed [ 9:0] r_sub10_T_addr;
	wire        [31:0] w_sub10_T_datain;
	reg         [31:0] r_sub10_T_datain;
	wire        [31:0] w_sub10_T_dataout;
	wire               w_sub10_T_r_w;
	reg                r_sub10_T_r_w;
	wire signed [ 9:0] w_sub10_V_addr;
	reg  signed [ 9:0] r_sub10_V_addr;
	wire        [31:0] w_sub10_V_datain;
	reg         [31:0] r_sub10_V_datain;
	wire        [31:0] w_sub10_V_dataout;
	wire               w_sub10_V_r_w;
	reg                r_sub10_V_r_w;
	wire signed [ 9:0] w_sub10_U_addr;
	reg  signed [ 9:0] r_sub10_U_addr;
	wire        [31:0] w_sub10_U_datain;
	reg         [31:0] r_sub10_U_datain;
	wire        [31:0] w_sub10_U_dataout;
	wire               w_sub10_U_r_w;
	reg                r_sub10_U_r_w;
	wire signed [ 9:0] w_sub10_result_addr;
	reg  signed [ 9:0] r_sub10_result_addr;
	wire        [31:0] w_sub10_result_datain;
	reg         [31:0] r_sub10_result_datain;
	wire        [31:0] w_sub10_result_dataout;
	wire               w_sub10_result_r_w;
	reg                r_sub10_result_r_w;
	reg                r_sub20_run_req;
	wire               w_sub20_run_busy;
	wire signed [ 9:0] w_sub20_T_addr;
	reg  signed [ 9:0] r_sub20_T_addr;
	wire        [31:0] w_sub20_T_datain;
	reg         [31:0] r_sub20_T_datain;
	wire        [31:0] w_sub20_T_dataout;
	wire               w_sub20_T_r_w;
	reg                r_sub20_T_r_w;
	wire signed [ 9:0] w_sub20_V_addr;
	reg  signed [ 9:0] r_sub20_V_addr;
	wire        [31:0] w_sub20_V_datain;
	reg         [31:0] r_sub20_V_datain;
	wire        [31:0] w_sub20_V_dataout;
	wire               w_sub20_V_r_w;
	reg                r_sub20_V_r_w;
	wire signed [ 9:0] w_sub20_U_addr;
	reg  signed [ 9:0] r_sub20_U_addr;
	wire        [31:0] w_sub20_U_datain;
	reg         [31:0] r_sub20_U_datain;
	wire        [31:0] w_sub20_U_dataout;
	wire               w_sub20_U_r_w;
	reg                r_sub20_U_r_w;
	wire signed [ 9:0] w_sub20_result_addr;
	reg  signed [ 9:0] r_sub20_result_addr;
	wire        [31:0] w_sub20_result_datain;
	reg         [31:0] r_sub20_result_datain;
	wire        [31:0] w_sub20_result_dataout;
	wire               w_sub20_result_r_w;
	reg                r_sub20_result_r_w;
	reg                r_sub21_run_req;
	wire               w_sub21_run_busy;
	wire signed [ 9:0] w_sub21_T_addr;
	reg  signed [ 9:0] r_sub21_T_addr;
	wire        [31:0] w_sub21_T_datain;
	reg         [31:0] r_sub21_T_datain;
	wire        [31:0] w_sub21_T_dataout;
	wire               w_sub21_T_r_w;
	reg                r_sub21_T_r_w;
	wire signed [ 9:0] w_sub21_V_addr;
	reg  signed [ 9:0] r_sub21_V_addr;
	wire        [31:0] w_sub21_V_datain;
	reg         [31:0] r_sub21_V_datain;
	wire        [31:0] w_sub21_V_dataout;
	wire               w_sub21_V_r_w;
	reg                r_sub21_V_r_w;
	wire signed [ 9:0] w_sub21_U_addr;
	reg  signed [ 9:0] r_sub21_U_addr;
	wire        [31:0] w_sub21_U_datain;
	reg         [31:0] r_sub21_U_datain;
	wire        [31:0] w_sub21_U_dataout;
	wire               w_sub21_U_r_w;
	reg                r_sub21_U_r_w;
	wire signed [ 9:0] w_sub21_result_addr;
	reg  signed [ 9:0] r_sub21_result_addr;
	wire        [31:0] w_sub21_result_datain;
	reg         [31:0] r_sub21_result_datain;
	wire        [31:0] w_sub21_result_dataout;
	wire               w_sub21_result_r_w;
	reg                r_sub21_result_r_w;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg         [31:0] r_sys_tmp4_float;
	reg         [31:0] r_sys_tmp5_float;
	reg         [31:0] r_sys_tmp6_float;
	reg         [31:0] r_sys_tmp7_float;
	reg         [31:0] r_sys_tmp8_float;
	reg         [31:0] r_sys_tmp9_float;
	reg         [31:0] r_sys_tmp10_float;
	reg         [31:0] r_sys_tmp11_float;
	reg         [31:0] r_sys_tmp12_float;
	reg         [31:0] r_sys_tmp13_float;
	reg         [31:0] r_sys_tmp14_float;
	reg         [31:0] r_sys_tmp15_float;
	reg         [31:0] r_sys_tmp16_float;
	reg         [31:0] r_sys_tmp17_float;
	reg         [31:0] r_sys_tmp18_float;
	reg         [31:0] r_sys_tmp19_float;
	reg         [31:0] r_sys_tmp20_float;
	reg         [31:0] r_sys_tmp21_float;
	reg         [31:0] r_sys_tmp22_float;
	reg         [31:0] r_sys_tmp23_float;
	reg         [31:0] r_sys_tmp24_float;
	reg         [31:0] r_sys_tmp25_float;
	reg         [31:0] r_sys_tmp26_float;
	reg         [31:0] r_sys_tmp27_float;
	reg         [31:0] r_sys_tmp28_float;
	reg         [31:0] r_sys_tmp29_float;
	reg         [31:0] r_sys_tmp30_float;
	reg         [31:0] r_sys_tmp31_float;
	reg         [31:0] r_sys_tmp32_float;
	reg         [31:0] r_sys_tmp33_float;
	reg         [31:0] r_sys_tmp34_float;
	reg         [31:0] r_sys_tmp35_float;
	reg         [31:0] r_sys_tmp36_float;
	reg         [31:0] r_sys_tmp37_float;
	reg         [31:0] r_sys_tmp38_float;
	reg         [31:0] r_sys_tmp39_float;
	reg         [31:0] r_sys_tmp40_float;
	reg         [31:0] r_sys_tmp41_float;
	reg         [31:0] r_sys_tmp42_float;
	reg         [31:0] r_sys_tmp43_float;
	reg         [31:0] r_sys_tmp44_float;
	reg         [31:0] r_sys_tmp45_float;
	reg         [31:0] r_sys_tmp46_float;
	reg         [31:0] r_sys_tmp47_float;
	reg         [31:0] r_sys_tmp48_float;
	reg         [31:0] r_sys_tmp49_float;
	reg         [31:0] r_sys_tmp50_float;
	reg         [31:0] r_sys_tmp51_float;
	reg         [31:0] r_sys_tmp52_float;
	reg         [31:0] r_sys_tmp53_float;
	reg         [31:0] r_sys_tmp54_float;
	reg         [31:0] r_sys_tmp55_float;
	reg         [31:0] r_sys_tmp56_float;
	reg         [31:0] r_sys_tmp57_float;
	reg         [31:0] r_sys_tmp58_float;
	reg         [31:0] r_sys_tmp59_float;
	reg         [31:0] r_sys_tmp60_float;
	reg         [31:0] r_sys_tmp61_float;
	reg         [31:0] r_sys_tmp62_float;
	reg         [31:0] r_sys_tmp63_float;
	reg         [31:0] r_sys_tmp64_float;
	reg         [31:0] r_sys_tmp65_float;
	reg         [31:0] r_sys_tmp66_float;
	reg         [31:0] r_sys_tmp67_float;
	reg         [31:0] r_sys_tmp68_float;
	reg         [31:0] r_sys_tmp69_float;
	reg         [31:0] r_sys_tmp70_float;
	reg         [31:0] r_sys_tmp71_float;
	reg         [31:0] r_sys_tmp72_float;
	reg         [31:0] r_sys_tmp73_float;
	reg         [31:0] r_sys_tmp74_float;
	reg         [31:0] r_sys_tmp75_float;
	reg         [31:0] r_sys_tmp76_float;
	reg         [31:0] r_sys_tmp77_float;
	reg         [31:0] r_sys_tmp78_float;
	reg         [31:0] r_sys_tmp79_float;
	reg         [31:0] r_sys_tmp80_float;
	reg         [31:0] r_sys_tmp81_float;
	reg         [31:0] r_sys_tmp82_float;
	reg         [31:0] r_sys_tmp83_float;
	reg         [31:0] r_sys_tmp84_float;
	reg         [31:0] r_sys_tmp85_float;
	reg         [31:0] r_sys_tmp86_float;
	reg         [31:0] r_sys_tmp87_float;
	reg         [31:0] r_sys_tmp88_float;
	reg         [31:0] r_sys_tmp89_float;
	reg         [31:0] r_sys_tmp90_float;
	reg         [31:0] r_sys_tmp91_float;
	reg         [31:0] r_sys_tmp92_float;
	reg         [31:0] r_sys_tmp93_float;
	reg         [31:0] r_sys_tmp94_float;
	reg         [31:0] r_sys_tmp95_float;
	reg         [31:0] r_sys_tmp96_float;
	reg         [31:0] r_sys_tmp97_float;
	reg         [31:0] r_sys_tmp98_float;
	reg         [31:0] r_sys_tmp99_float;
	reg         [31:0] r_sys_tmp100_float;
	reg         [31:0] r_sys_tmp101_float;
	reg         [31:0] r_sys_tmp102_float;
	reg         [31:0] r_sys_tmp103_float;
	reg         [31:0] r_sys_tmp104_float;
	reg         [31:0] r_sys_tmp105_float;
	reg         [31:0] r_sys_tmp106_float;
	reg         [31:0] r_sys_tmp107_float;
	reg         [31:0] r_sys_tmp108_float;
	reg         [31:0] r_sys_tmp109_float;
	wire signed [31:0] w_sys_tmp1;
	wire signed [31:0] w_sys_tmp3;
	wire        [31:0] w_sys_tmp5;
	wire signed [31:0] w_sys_tmp6;
	wire        [31:0] w_sys_tmp7;
	wire        [31:0] w_sys_tmp8;
	wire        [31:0] w_sys_tmp9;
	wire        [31:0] w_sys_tmp10;
	wire        [31:0] w_sys_tmp11;
	wire        [31:0] w_sys_tmp12;
	wire               w_sys_tmp13;
	wire               w_sys_tmp14;
	wire signed [31:0] w_sys_tmp15;
	wire               w_sys_tmp16;
	wire               w_sys_tmp17;
	wire        [31:0] w_sys_tmp19;
	wire        [31:0] w_sys_tmp20;
	wire signed [31:0] w_sys_tmp21;
	wire signed [31:0] w_sys_tmp23;
	wire signed [31:0] w_sys_tmp24;
	wire signed [31:0] w_sys_tmp25;
	wire        [31:0] w_sys_tmp26;
	wire signed [31:0] w_sys_tmp28;
	wire signed [31:0] w_sys_tmp29;
	wire signed [31:0] w_sys_tmp33;
	wire signed [31:0] w_sys_tmp34;
	wire        [31:0] w_sys_tmp37;
	wire        [31:0] w_sys_tmp38;
	wire        [31:0] w_sys_tmp39;
	wire signed [31:0] w_sys_tmp42;
	wire signed [31:0] w_sys_tmp43;
	wire signed [31:0] w_sys_tmp46;
	wire signed [31:0] w_sys_tmp47;
	wire signed [31:0] w_sys_tmp48;
	wire signed [31:0] w_sys_tmp49;
	wire        [31:0] w_sys_tmp129;
	wire               w_sys_tmp227;
	wire               w_sys_tmp228;
	wire signed [31:0] w_sys_tmp229;
	wire signed [31:0] w_sys_tmp232;
	wire signed [31:0] w_sys_tmp233;
	wire        [31:0] w_sys_tmp234;
	wire        [31:0] w_sys_tmp240;
	wire signed [31:0] w_sys_tmp244;
	wire signed [31:0] w_sys_tmp245;
	wire signed [31:0] w_sys_tmp256;
	wire signed [31:0] w_sys_tmp257;
	wire signed [31:0] w_sys_tmp268;
	wire signed [31:0] w_sys_tmp269;
	wire signed [31:0] w_sys_tmp280;
	wire signed [31:0] w_sys_tmp281;
	wire signed [31:0] w_sys_tmp292;
	wire signed [31:0] w_sys_tmp293;
	wire signed [31:0] w_sys_tmp304;
	wire signed [31:0] w_sys_tmp305;
	wire signed [31:0] w_sys_tmp316;
	wire signed [31:0] w_sys_tmp317;
	wire signed [31:0] w_sys_tmp352;
	wire signed [31:0] w_sys_tmp353;
	wire signed [31:0] w_sys_tmp364;
	wire signed [31:0] w_sys_tmp365;
	wire signed [31:0] w_sys_tmp376;
	wire signed [31:0] w_sys_tmp377;
	wire signed [31:0] w_sys_tmp388;
	wire signed [31:0] w_sys_tmp389;
	wire signed [31:0] w_sys_tmp400;
	wire signed [31:0] w_sys_tmp401;
	wire signed [31:0] w_sys_tmp412;
	wire signed [31:0] w_sys_tmp413;
	wire signed [31:0] w_sys_tmp448;
	wire signed [31:0] w_sys_tmp449;
	wire signed [31:0] w_sys_tmp460;
	wire signed [31:0] w_sys_tmp461;
	wire signed [31:0] w_sys_tmp472;
	wire signed [31:0] w_sys_tmp473;
	wire signed [31:0] w_sys_tmp484;
	wire signed [31:0] w_sys_tmp485;
	wire signed [31:0] w_sys_tmp496;
	wire signed [31:0] w_sys_tmp497;
	wire signed [31:0] w_sys_tmp508;
	wire signed [31:0] w_sys_tmp509;
	wire signed [31:0] w_sys_tmp544;
	wire signed [31:0] w_sys_tmp545;
	wire signed [31:0] w_sys_tmp556;
	wire signed [31:0] w_sys_tmp557;
	wire signed [31:0] w_sys_tmp568;
	wire signed [31:0] w_sys_tmp569;
	wire signed [31:0] w_sys_tmp580;
	wire signed [31:0] w_sys_tmp581;
	wire signed [31:0] w_sys_tmp592;
	wire signed [31:0] w_sys_tmp593;
	wire signed [31:0] w_sys_tmp604;
	wire signed [31:0] w_sys_tmp605;
	wire signed [31:0] w_sys_tmp640;
	wire signed [31:0] w_sys_tmp641;
	wire signed [31:0] w_sys_tmp652;
	wire signed [31:0] w_sys_tmp653;
	wire signed [31:0] w_sys_tmp664;
	wire signed [31:0] w_sys_tmp665;
	wire signed [31:0] w_sys_tmp676;
	wire signed [31:0] w_sys_tmp677;
	wire signed [31:0] w_sys_tmp688;
	wire signed [31:0] w_sys_tmp689;
	wire signed [31:0] w_sys_tmp700;
	wire signed [31:0] w_sys_tmp701;
	wire signed [31:0] w_sys_tmp712;
	wire signed [31:0] w_sys_tmp713;
	wire signed [31:0] w_sys_tmp724;
	wire signed [31:0] w_sys_tmp725;
	wire signed [31:0] w_sys_tmp736;
	wire signed [31:0] w_sys_tmp737;
	wire signed [31:0] w_sys_tmp748;
	wire signed [31:0] w_sys_tmp749;
	wire signed [31:0] w_sys_tmp760;
	wire signed [31:0] w_sys_tmp761;
	wire signed [31:0] w_sys_tmp772;
	wire signed [31:0] w_sys_tmp773;
	wire signed [31:0] w_sys_tmp784;
	wire signed [31:0] w_sys_tmp785;
	wire signed [31:0] w_sys_tmp820;
	wire signed [31:0] w_sys_tmp821;
	wire signed [31:0] w_sys_tmp832;
	wire signed [31:0] w_sys_tmp833;
	wire signed [31:0] w_sys_tmp844;
	wire signed [31:0] w_sys_tmp845;
	wire signed [31:0] w_sys_tmp856;
	wire signed [31:0] w_sys_tmp857;
	wire signed [31:0] w_sys_tmp868;
	wire signed [31:0] w_sys_tmp869;
	wire signed [31:0] w_sys_tmp880;
	wire signed [31:0] w_sys_tmp881;
	wire signed [31:0] w_sys_tmp916;
	wire signed [31:0] w_sys_tmp917;
	wire signed [31:0] w_sys_tmp928;
	wire signed [31:0] w_sys_tmp929;
	wire signed [31:0] w_sys_tmp940;
	wire signed [31:0] w_sys_tmp941;
	wire signed [31:0] w_sys_tmp952;
	wire signed [31:0] w_sys_tmp953;
	wire signed [31:0] w_sys_tmp964;
	wire signed [31:0] w_sys_tmp965;
	wire signed [31:0] w_sys_tmp976;
	wire signed [31:0] w_sys_tmp977;
	wire signed [31:0] w_sys_tmp1012;
	wire signed [31:0] w_sys_tmp1013;
	wire signed [31:0] w_sys_tmp1024;
	wire signed [31:0] w_sys_tmp1025;
	wire signed [31:0] w_sys_tmp1036;
	wire signed [31:0] w_sys_tmp1037;
	wire signed [31:0] w_sys_tmp1048;
	wire signed [31:0] w_sys_tmp1049;
	wire signed [31:0] w_sys_tmp1060;
	wire signed [31:0] w_sys_tmp1061;
	wire signed [31:0] w_sys_tmp1072;
	wire signed [31:0] w_sys_tmp1073;
	wire signed [31:0] w_sys_tmp1108;
	wire signed [31:0] w_sys_tmp1109;
	wire signed [31:0] w_sys_tmp1120;
	wire signed [31:0] w_sys_tmp1121;
	wire signed [31:0] w_sys_tmp1132;
	wire signed [31:0] w_sys_tmp1133;
	wire signed [31:0] w_sys_tmp1144;
	wire signed [31:0] w_sys_tmp1145;
	wire signed [31:0] w_sys_tmp1156;
	wire signed [31:0] w_sys_tmp1157;
	wire signed [31:0] w_sys_tmp1168;
	wire signed [31:0] w_sys_tmp1169;
	wire signed [31:0] w_sys_tmp1180;
	wire signed [31:0] w_sys_tmp1181;
	wire signed [31:0] w_sys_tmp1192;
	wire signed [31:0] w_sys_tmp1193;
	wire signed [31:0] w_sys_tmp1204;
	wire signed [31:0] w_sys_tmp1205;
	wire signed [31:0] w_sys_tmp1216;
	wire signed [31:0] w_sys_tmp1217;
	wire signed [31:0] w_sys_tmp1228;
	wire signed [31:0] w_sys_tmp1229;
	wire signed [31:0] w_sys_tmp1240;
	wire signed [31:0] w_sys_tmp1241;
	wire signed [31:0] w_sys_tmp1252;
	wire signed [31:0] w_sys_tmp1253;
	wire signed [31:0] w_sys_tmp1288;
	wire signed [31:0] w_sys_tmp1289;
	wire signed [31:0] w_sys_tmp1300;
	wire signed [31:0] w_sys_tmp1301;
	wire signed [31:0] w_sys_tmp1312;
	wire signed [31:0] w_sys_tmp1313;
	wire signed [31:0] w_sys_tmp1324;
	wire signed [31:0] w_sys_tmp1325;
	wire signed [31:0] w_sys_tmp1336;
	wire signed [31:0] w_sys_tmp1337;
	wire signed [31:0] w_sys_tmp1348;
	wire signed [31:0] w_sys_tmp1349;
	wire signed [31:0] w_sys_tmp1384;
	wire signed [31:0] w_sys_tmp1385;
	wire signed [31:0] w_sys_tmp1396;
	wire signed [31:0] w_sys_tmp1397;
	wire signed [31:0] w_sys_tmp1408;
	wire signed [31:0] w_sys_tmp1409;
	wire signed [31:0] w_sys_tmp1420;
	wire signed [31:0] w_sys_tmp1421;
	wire signed [31:0] w_sys_tmp1432;
	wire signed [31:0] w_sys_tmp1433;
	wire signed [31:0] w_sys_tmp1444;
	wire signed [31:0] w_sys_tmp1445;
	wire signed [31:0] w_sys_tmp1480;
	wire signed [31:0] w_sys_tmp1481;
	wire signed [31:0] w_sys_tmp1492;
	wire signed [31:0] w_sys_tmp1493;
	wire signed [31:0] w_sys_tmp1504;
	wire signed [31:0] w_sys_tmp1505;
	wire signed [31:0] w_sys_tmp1516;
	wire signed [31:0] w_sys_tmp1517;
	wire signed [31:0] w_sys_tmp1528;
	wire signed [31:0] w_sys_tmp1529;
	wire signed [31:0] w_sys_tmp1540;
	wire signed [31:0] w_sys_tmp1541;
	wire signed [31:0] w_sys_tmp1576;
	wire signed [31:0] w_sys_tmp1577;
	wire signed [31:0] w_sys_tmp1588;
	wire signed [31:0] w_sys_tmp1589;
	wire signed [31:0] w_sys_tmp1600;
	wire signed [31:0] w_sys_tmp1601;
	wire signed [31:0] w_sys_tmp1612;
	wire signed [31:0] w_sys_tmp1613;
	wire signed [31:0] w_sys_tmp1624;
	wire signed [31:0] w_sys_tmp1625;
	wire signed [31:0] w_sys_tmp1636;
	wire signed [31:0] w_sys_tmp1637;
	wire signed [31:0] w_sys_tmp1648;
	wire signed [31:0] w_sys_tmp1649;
	wire signed [31:0] w_sys_tmp1660;
	wire signed [31:0] w_sys_tmp1661;
	wire signed [31:0] w_sys_tmp1672;
	wire signed [31:0] w_sys_tmp1673;
	wire signed [31:0] w_sys_tmp1684;
	wire signed [31:0] w_sys_tmp1685;
	wire signed [31:0] w_sys_tmp1696;
	wire signed [31:0] w_sys_tmp1697;
	wire signed [31:0] w_sys_tmp1708;
	wire signed [31:0] w_sys_tmp1709;
	wire signed [31:0] w_sys_tmp1720;
	wire signed [31:0] w_sys_tmp1721;
	wire signed [31:0] w_sys_tmp1756;
	wire signed [31:0] w_sys_tmp1757;
	wire signed [31:0] w_sys_tmp1768;
	wire signed [31:0] w_sys_tmp1769;
	wire signed [31:0] w_sys_tmp1780;
	wire signed [31:0] w_sys_tmp1781;
	wire signed [31:0] w_sys_tmp1792;
	wire signed [31:0] w_sys_tmp1793;
	wire signed [31:0] w_sys_tmp1804;
	wire signed [31:0] w_sys_tmp1805;
	wire signed [31:0] w_sys_tmp1816;
	wire signed [31:0] w_sys_tmp1817;
	wire signed [31:0] w_sys_tmp1852;
	wire signed [31:0] w_sys_tmp1853;
	wire signed [31:0] w_sys_tmp1864;
	wire signed [31:0] w_sys_tmp1865;
	wire signed [31:0] w_sys_tmp1876;
	wire signed [31:0] w_sys_tmp1877;
	wire signed [31:0] w_sys_tmp1888;
	wire signed [31:0] w_sys_tmp1889;
	wire signed [31:0] w_sys_tmp1900;
	wire signed [31:0] w_sys_tmp1901;
	wire signed [31:0] w_sys_tmp1912;
	wire signed [31:0] w_sys_tmp1913;
	wire signed [31:0] w_sys_tmp1948;
	wire signed [31:0] w_sys_tmp1949;
	wire signed [31:0] w_sys_tmp1960;
	wire signed [31:0] w_sys_tmp1961;
	wire signed [31:0] w_sys_tmp1972;
	wire signed [31:0] w_sys_tmp1973;
	wire signed [31:0] w_sys_tmp1984;
	wire signed [31:0] w_sys_tmp1985;
	wire signed [31:0] w_sys_tmp1996;
	wire signed [31:0] w_sys_tmp1997;
	wire signed [31:0] w_sys_tmp2008;
	wire signed [31:0] w_sys_tmp2009;
	wire signed [31:0] w_sys_tmp2044;
	wire signed [31:0] w_sys_tmp2045;
	wire signed [31:0] w_sys_tmp2056;
	wire signed [31:0] w_sys_tmp2057;
	wire signed [31:0] w_sys_tmp2068;
	wire signed [31:0] w_sys_tmp2069;
	wire signed [31:0] w_sys_tmp2080;
	wire signed [31:0] w_sys_tmp2081;
	wire signed [31:0] w_sys_tmp2092;
	wire signed [31:0] w_sys_tmp2093;
	wire signed [31:0] w_sys_tmp2103;
	wire signed [31:0] w_sys_tmp2104;
	wire               w_sys_tmp2105;
	wire               w_sys_tmp2106;
	wire signed [31:0] w_sys_tmp2107;
	wire signed [31:0] w_sys_tmp2110;
	wire signed [31:0] w_sys_tmp2111;
	wire        [31:0] w_sys_tmp2112;
	wire        [31:0] w_sys_tmp2118;
	wire signed [31:0] w_sys_tmp2122;
	wire signed [31:0] w_sys_tmp2123;
	wire signed [31:0] w_sys_tmp2134;
	wire signed [31:0] w_sys_tmp2135;
	wire signed [31:0] w_sys_tmp2146;
	wire signed [31:0] w_sys_tmp2147;
	wire signed [31:0] w_sys_tmp2158;
	wire signed [31:0] w_sys_tmp2159;
	wire signed [31:0] w_sys_tmp2170;
	wire signed [31:0] w_sys_tmp2171;
	wire signed [31:0] w_sys_tmp2182;
	wire signed [31:0] w_sys_tmp2183;
	wire signed [31:0] w_sys_tmp2194;
	wire signed [31:0] w_sys_tmp2195;
	wire signed [31:0] w_sys_tmp2230;
	wire signed [31:0] w_sys_tmp2231;
	wire signed [31:0] w_sys_tmp2242;
	wire signed [31:0] w_sys_tmp2243;
	wire signed [31:0] w_sys_tmp2254;
	wire signed [31:0] w_sys_tmp2255;
	wire signed [31:0] w_sys_tmp2266;
	wire signed [31:0] w_sys_tmp2267;
	wire signed [31:0] w_sys_tmp2278;
	wire signed [31:0] w_sys_tmp2279;
	wire signed [31:0] w_sys_tmp2290;
	wire signed [31:0] w_sys_tmp2291;
	wire signed [31:0] w_sys_tmp2326;
	wire signed [31:0] w_sys_tmp2327;
	wire signed [31:0] w_sys_tmp2338;
	wire signed [31:0] w_sys_tmp2339;
	wire signed [31:0] w_sys_tmp2350;
	wire signed [31:0] w_sys_tmp2351;
	wire signed [31:0] w_sys_tmp2362;
	wire signed [31:0] w_sys_tmp2363;
	wire signed [31:0] w_sys_tmp2374;
	wire signed [31:0] w_sys_tmp2375;
	wire signed [31:0] w_sys_tmp2386;
	wire signed [31:0] w_sys_tmp2387;
	wire signed [31:0] w_sys_tmp2422;
	wire signed [31:0] w_sys_tmp2423;
	wire signed [31:0] w_sys_tmp2434;
	wire signed [31:0] w_sys_tmp2435;
	wire signed [31:0] w_sys_tmp2446;
	wire signed [31:0] w_sys_tmp2447;
	wire signed [31:0] w_sys_tmp2458;
	wire signed [31:0] w_sys_tmp2459;
	wire signed [31:0] w_sys_tmp2470;
	wire signed [31:0] w_sys_tmp2471;
	wire signed [31:0] w_sys_tmp2482;
	wire signed [31:0] w_sys_tmp2483;
	wire signed [31:0] w_sys_tmp2518;
	wire signed [31:0] w_sys_tmp2519;
	wire signed [31:0] w_sys_tmp2530;
	wire signed [31:0] w_sys_tmp2531;
	wire signed [31:0] w_sys_tmp2542;
	wire signed [31:0] w_sys_tmp2543;
	wire signed [31:0] w_sys_tmp2554;
	wire signed [31:0] w_sys_tmp2555;
	wire signed [31:0] w_sys_tmp2566;
	wire signed [31:0] w_sys_tmp2567;
	wire signed [31:0] w_sys_tmp2577;
	wire               w_sys_tmp2578;
	wire               w_sys_tmp2579;
	wire signed [31:0] w_sys_tmp2580;
	wire               w_sys_tmp2581;
	wire               w_sys_tmp2582;
	wire signed [31:0] w_sys_tmp2585;
	wire signed [31:0] w_sys_tmp2586;
	wire        [31:0] w_sys_tmp2587;
	wire signed [31:0] w_sys_tmp2589;
	wire signed [31:0] w_sys_tmp2590;
	wire        [31:0] w_sys_tmp2592;
	wire signed [31:0] w_sys_tmp2593;
	wire signed [31:0] w_sys_tmp2594;
	wire signed [31:0] w_sys_tmp2595;
	wire signed [31:0] w_sys_tmp2597;
	wire               w_sys_tmp2598;
	wire               w_sys_tmp2599;
	wire signed [31:0] w_sys_tmp2602;
	wire signed [31:0] w_sys_tmp2603;
	wire signed [31:0] w_sys_tmp2604;
	wire        [31:0] w_sys_tmp2605;
	wire signed [31:0] w_sys_tmp2607;
	wire signed [31:0] w_sys_tmp2608;
	wire signed [31:0] w_sys_tmp2611;
	wire signed [31:0] w_sys_tmp2612;
	wire signed [31:0] w_sys_tmp2685;
	wire signed [31:0] w_sys_tmp2686;
	wire               w_sys_tmp2687;
	wire               w_sys_tmp2688;
	wire signed [31:0] w_sys_tmp2689;
	wire signed [31:0] w_sys_tmp2690;
	wire signed [31:0] w_sys_tmp2693;
	wire signed [31:0] w_sys_tmp2694;
	wire signed [31:0] w_sys_tmp2695;
	wire        [31:0] w_sys_tmp2696;
	wire signed [31:0] w_sys_tmp2697;
	wire               w_sys_tmp2734;
	wire               w_sys_tmp2735;
	wire signed [31:0] w_sys_tmp2736;
	wire signed [31:0] w_sys_tmp2739;
	wire signed [31:0] w_sys_tmp2740;
	wire        [31:0] w_sys_tmp2741;
	wire signed [31:0] w_sys_tmp2745;
	wire signed [31:0] w_sys_tmp2746;
	wire signed [31:0] w_sys_tmp2751;
	wire signed [31:0] w_sys_tmp2752;
	wire signed [31:0] w_sys_tmp2757;
	wire signed [31:0] w_sys_tmp2758;
	wire signed [31:0] w_sys_tmp2763;
	wire signed [31:0] w_sys_tmp2764;
	wire signed [31:0] w_sys_tmp2769;
	wire signed [31:0] w_sys_tmp2770;
	wire signed [31:0] w_sys_tmp2775;
	wire signed [31:0] w_sys_tmp2776;
	wire signed [31:0] w_sys_tmp2781;
	wire signed [31:0] w_sys_tmp2782;
	wire signed [31:0] w_sys_tmp2799;
	wire signed [31:0] w_sys_tmp2800;
	wire signed [31:0] w_sys_tmp2805;
	wire signed [31:0] w_sys_tmp2806;
	wire signed [31:0] w_sys_tmp2811;
	wire signed [31:0] w_sys_tmp2812;
	wire signed [31:0] w_sys_tmp2817;
	wire signed [31:0] w_sys_tmp2818;
	wire signed [31:0] w_sys_tmp2823;
	wire signed [31:0] w_sys_tmp2824;
	wire signed [31:0] w_sys_tmp2829;
	wire signed [31:0] w_sys_tmp2830;
	wire signed [31:0] w_sys_tmp2847;
	wire signed [31:0] w_sys_tmp2848;
	wire signed [31:0] w_sys_tmp2853;
	wire signed [31:0] w_sys_tmp2854;
	wire signed [31:0] w_sys_tmp2859;
	wire signed [31:0] w_sys_tmp2860;
	wire signed [31:0] w_sys_tmp2865;
	wire signed [31:0] w_sys_tmp2866;
	wire signed [31:0] w_sys_tmp2871;
	wire signed [31:0] w_sys_tmp2872;
	wire signed [31:0] w_sys_tmp2877;
	wire signed [31:0] w_sys_tmp2878;
	wire signed [31:0] w_sys_tmp2895;
	wire signed [31:0] w_sys_tmp2896;
	wire signed [31:0] w_sys_tmp2901;
	wire signed [31:0] w_sys_tmp2902;
	wire signed [31:0] w_sys_tmp2907;
	wire signed [31:0] w_sys_tmp2908;
	wire signed [31:0] w_sys_tmp2913;
	wire signed [31:0] w_sys_tmp2914;
	wire signed [31:0] w_sys_tmp2919;
	wire signed [31:0] w_sys_tmp2920;
	wire signed [31:0] w_sys_tmp2925;
	wire signed [31:0] w_sys_tmp2926;
	wire signed [31:0] w_sys_tmp2943;
	wire signed [31:0] w_sys_tmp2944;
	wire signed [31:0] w_sys_tmp2949;
	wire signed [31:0] w_sys_tmp2950;
	wire signed [31:0] w_sys_tmp2955;
	wire signed [31:0] w_sys_tmp2956;
	wire signed [31:0] w_sys_tmp2961;
	wire signed [31:0] w_sys_tmp2962;
	wire signed [31:0] w_sys_tmp2967;
	wire signed [31:0] w_sys_tmp2968;
	wire signed [31:0] w_sys_tmp2973;
	wire signed [31:0] w_sys_tmp2974;
	wire signed [31:0] w_sys_tmp2979;
	wire signed [31:0] w_sys_tmp2980;
	wire signed [31:0] w_sys_tmp2985;
	wire signed [31:0] w_sys_tmp2986;
	wire signed [31:0] w_sys_tmp2991;
	wire signed [31:0] w_sys_tmp2992;
	wire signed [31:0] w_sys_tmp2997;
	wire signed [31:0] w_sys_tmp2998;
	wire signed [31:0] w_sys_tmp3003;
	wire signed [31:0] w_sys_tmp3004;
	wire signed [31:0] w_sys_tmp3009;
	wire signed [31:0] w_sys_tmp3010;
	wire signed [31:0] w_sys_tmp3015;
	wire signed [31:0] w_sys_tmp3016;
	wire signed [31:0] w_sys_tmp3033;
	wire signed [31:0] w_sys_tmp3034;
	wire signed [31:0] w_sys_tmp3039;
	wire signed [31:0] w_sys_tmp3040;
	wire signed [31:0] w_sys_tmp3045;
	wire signed [31:0] w_sys_tmp3046;
	wire signed [31:0] w_sys_tmp3051;
	wire signed [31:0] w_sys_tmp3052;
	wire signed [31:0] w_sys_tmp3057;
	wire signed [31:0] w_sys_tmp3058;
	wire signed [31:0] w_sys_tmp3063;
	wire signed [31:0] w_sys_tmp3064;
	wire signed [31:0] w_sys_tmp3081;
	wire signed [31:0] w_sys_tmp3082;
	wire signed [31:0] w_sys_tmp3087;
	wire signed [31:0] w_sys_tmp3088;
	wire signed [31:0] w_sys_tmp3093;
	wire signed [31:0] w_sys_tmp3094;
	wire signed [31:0] w_sys_tmp3099;
	wire signed [31:0] w_sys_tmp3100;
	wire signed [31:0] w_sys_tmp3105;
	wire signed [31:0] w_sys_tmp3106;
	wire signed [31:0] w_sys_tmp3111;
	wire signed [31:0] w_sys_tmp3112;
	wire signed [31:0] w_sys_tmp3129;
	wire signed [31:0] w_sys_tmp3130;
	wire signed [31:0] w_sys_tmp3135;
	wire signed [31:0] w_sys_tmp3136;
	wire signed [31:0] w_sys_tmp3141;
	wire signed [31:0] w_sys_tmp3142;
	wire signed [31:0] w_sys_tmp3147;
	wire signed [31:0] w_sys_tmp3148;
	wire signed [31:0] w_sys_tmp3153;
	wire signed [31:0] w_sys_tmp3154;
	wire signed [31:0] w_sys_tmp3159;
	wire signed [31:0] w_sys_tmp3160;
	wire signed [31:0] w_sys_tmp3177;
	wire signed [31:0] w_sys_tmp3178;
	wire signed [31:0] w_sys_tmp3183;
	wire signed [31:0] w_sys_tmp3184;
	wire signed [31:0] w_sys_tmp3189;
	wire signed [31:0] w_sys_tmp3190;
	wire signed [31:0] w_sys_tmp3195;
	wire signed [31:0] w_sys_tmp3196;
	wire signed [31:0] w_sys_tmp3201;
	wire signed [31:0] w_sys_tmp3202;
	wire signed [31:0] w_sys_tmp3207;
	wire signed [31:0] w_sys_tmp3208;
	wire signed [31:0] w_sys_tmp3213;
	wire signed [31:0] w_sys_tmp3214;
	wire signed [31:0] w_sys_tmp3219;
	wire signed [31:0] w_sys_tmp3220;
	wire signed [31:0] w_sys_tmp3225;
	wire signed [31:0] w_sys_tmp3226;
	wire signed [31:0] w_sys_tmp3231;
	wire signed [31:0] w_sys_tmp3232;
	wire signed [31:0] w_sys_tmp3237;
	wire signed [31:0] w_sys_tmp3238;
	wire signed [31:0] w_sys_tmp3243;
	wire signed [31:0] w_sys_tmp3244;
	wire signed [31:0] w_sys_tmp3249;
	wire signed [31:0] w_sys_tmp3250;
	wire signed [31:0] w_sys_tmp3267;
	wire signed [31:0] w_sys_tmp3268;
	wire signed [31:0] w_sys_tmp3273;
	wire signed [31:0] w_sys_tmp3274;
	wire signed [31:0] w_sys_tmp3279;
	wire signed [31:0] w_sys_tmp3280;
	wire signed [31:0] w_sys_tmp3285;
	wire signed [31:0] w_sys_tmp3286;
	wire signed [31:0] w_sys_tmp3291;
	wire signed [31:0] w_sys_tmp3292;
	wire signed [31:0] w_sys_tmp3297;
	wire signed [31:0] w_sys_tmp3298;
	wire signed [31:0] w_sys_tmp3315;
	wire signed [31:0] w_sys_tmp3316;
	wire signed [31:0] w_sys_tmp3321;
	wire signed [31:0] w_sys_tmp3322;
	wire signed [31:0] w_sys_tmp3327;
	wire signed [31:0] w_sys_tmp3328;
	wire signed [31:0] w_sys_tmp3333;
	wire signed [31:0] w_sys_tmp3334;
	wire signed [31:0] w_sys_tmp3339;
	wire signed [31:0] w_sys_tmp3340;
	wire signed [31:0] w_sys_tmp3345;
	wire signed [31:0] w_sys_tmp3346;
	wire signed [31:0] w_sys_tmp3363;
	wire signed [31:0] w_sys_tmp3364;
	wire signed [31:0] w_sys_tmp3369;
	wire signed [31:0] w_sys_tmp3370;
	wire signed [31:0] w_sys_tmp3375;
	wire signed [31:0] w_sys_tmp3376;
	wire signed [31:0] w_sys_tmp3381;
	wire signed [31:0] w_sys_tmp3382;
	wire signed [31:0] w_sys_tmp3387;
	wire signed [31:0] w_sys_tmp3388;
	wire signed [31:0] w_sys_tmp3393;
	wire signed [31:0] w_sys_tmp3394;
	wire signed [31:0] w_sys_tmp3411;
	wire signed [31:0] w_sys_tmp3412;
	wire signed [31:0] w_sys_tmp3417;
	wire signed [31:0] w_sys_tmp3418;
	wire signed [31:0] w_sys_tmp3423;
	wire signed [31:0] w_sys_tmp3424;
	wire signed [31:0] w_sys_tmp3429;
	wire signed [31:0] w_sys_tmp3430;
	wire signed [31:0] w_sys_tmp3435;
	wire signed [31:0] w_sys_tmp3436;
	wire signed [31:0] w_sys_tmp3441;
	wire signed [31:0] w_sys_tmp3442;
	wire signed [31:0] w_sys_tmp3447;
	wire signed [31:0] w_sys_tmp3448;
	wire signed [31:0] w_sys_tmp3453;
	wire signed [31:0] w_sys_tmp3454;
	wire signed [31:0] w_sys_tmp3459;
	wire signed [31:0] w_sys_tmp3460;
	wire signed [31:0] w_sys_tmp3465;
	wire signed [31:0] w_sys_tmp3466;
	wire signed [31:0] w_sys_tmp3471;
	wire signed [31:0] w_sys_tmp3472;
	wire signed [31:0] w_sys_tmp3477;
	wire signed [31:0] w_sys_tmp3478;
	wire signed [31:0] w_sys_tmp3483;
	wire signed [31:0] w_sys_tmp3484;
	wire signed [31:0] w_sys_tmp3501;
	wire signed [31:0] w_sys_tmp3502;
	wire signed [31:0] w_sys_tmp3507;
	wire signed [31:0] w_sys_tmp3508;
	wire signed [31:0] w_sys_tmp3513;
	wire signed [31:0] w_sys_tmp3514;
	wire signed [31:0] w_sys_tmp3519;
	wire signed [31:0] w_sys_tmp3520;
	wire signed [31:0] w_sys_tmp3525;
	wire signed [31:0] w_sys_tmp3526;
	wire signed [31:0] w_sys_tmp3531;
	wire signed [31:0] w_sys_tmp3532;
	wire signed [31:0] w_sys_tmp3549;
	wire signed [31:0] w_sys_tmp3550;
	wire signed [31:0] w_sys_tmp3555;
	wire signed [31:0] w_sys_tmp3556;
	wire signed [31:0] w_sys_tmp3561;
	wire signed [31:0] w_sys_tmp3562;
	wire signed [31:0] w_sys_tmp3567;
	wire signed [31:0] w_sys_tmp3568;
	wire signed [31:0] w_sys_tmp3573;
	wire signed [31:0] w_sys_tmp3574;
	wire signed [31:0] w_sys_tmp3579;
	wire signed [31:0] w_sys_tmp3580;
	wire signed [31:0] w_sys_tmp3597;
	wire signed [31:0] w_sys_tmp3598;
	wire signed [31:0] w_sys_tmp3603;
	wire signed [31:0] w_sys_tmp3604;
	wire signed [31:0] w_sys_tmp3609;
	wire signed [31:0] w_sys_tmp3610;
	wire signed [31:0] w_sys_tmp3615;
	wire signed [31:0] w_sys_tmp3616;
	wire signed [31:0] w_sys_tmp3621;
	wire signed [31:0] w_sys_tmp3622;
	wire signed [31:0] w_sys_tmp3627;
	wire signed [31:0] w_sys_tmp3628;
	wire signed [31:0] w_sys_tmp3645;
	wire signed [31:0] w_sys_tmp3646;
	wire signed [31:0] w_sys_tmp3651;
	wire signed [31:0] w_sys_tmp3652;
	wire signed [31:0] w_sys_tmp3657;
	wire signed [31:0] w_sys_tmp3658;
	wire signed [31:0] w_sys_tmp3663;
	wire signed [31:0] w_sys_tmp3664;
	wire signed [31:0] w_sys_tmp3669;
	wire signed [31:0] w_sys_tmp3670;
	wire signed [31:0] w_sys_tmp3674;
	wire signed [31:0] w_sys_tmp3675;
	wire               w_sys_tmp3676;
	wire               w_sys_tmp3677;
	wire signed [31:0] w_sys_tmp3678;
	wire signed [31:0] w_sys_tmp3681;
	wire signed [31:0] w_sys_tmp3682;
	wire        [31:0] w_sys_tmp3683;
	wire signed [31:0] w_sys_tmp3687;
	wire signed [31:0] w_sys_tmp3688;
	wire signed [31:0] w_sys_tmp3693;
	wire signed [31:0] w_sys_tmp3694;
	wire signed [31:0] w_sys_tmp3699;
	wire signed [31:0] w_sys_tmp3700;
	wire signed [31:0] w_sys_tmp3705;
	wire signed [31:0] w_sys_tmp3706;
	wire signed [31:0] w_sys_tmp3711;
	wire signed [31:0] w_sys_tmp3712;
	wire signed [31:0] w_sys_tmp3717;
	wire signed [31:0] w_sys_tmp3718;
	wire signed [31:0] w_sys_tmp3723;
	wire signed [31:0] w_sys_tmp3724;
	wire signed [31:0] w_sys_tmp3741;
	wire signed [31:0] w_sys_tmp3742;
	wire signed [31:0] w_sys_tmp3747;
	wire signed [31:0] w_sys_tmp3748;
	wire signed [31:0] w_sys_tmp3753;
	wire signed [31:0] w_sys_tmp3754;
	wire signed [31:0] w_sys_tmp3759;
	wire signed [31:0] w_sys_tmp3760;
	wire signed [31:0] w_sys_tmp3765;
	wire signed [31:0] w_sys_tmp3766;
	wire signed [31:0] w_sys_tmp3771;
	wire signed [31:0] w_sys_tmp3772;
	wire signed [31:0] w_sys_tmp3789;
	wire signed [31:0] w_sys_tmp3790;
	wire signed [31:0] w_sys_tmp3795;
	wire signed [31:0] w_sys_tmp3796;
	wire signed [31:0] w_sys_tmp3801;
	wire signed [31:0] w_sys_tmp3802;
	wire signed [31:0] w_sys_tmp3807;
	wire signed [31:0] w_sys_tmp3808;
	wire signed [31:0] w_sys_tmp3813;
	wire signed [31:0] w_sys_tmp3814;
	wire signed [31:0] w_sys_tmp3819;
	wire signed [31:0] w_sys_tmp3820;
	wire signed [31:0] w_sys_tmp3837;
	wire signed [31:0] w_sys_tmp3838;
	wire signed [31:0] w_sys_tmp3843;
	wire signed [31:0] w_sys_tmp3844;
	wire signed [31:0] w_sys_tmp3849;
	wire signed [31:0] w_sys_tmp3850;
	wire signed [31:0] w_sys_tmp3855;
	wire signed [31:0] w_sys_tmp3856;
	wire signed [31:0] w_sys_tmp3861;
	wire signed [31:0] w_sys_tmp3862;
	wire signed [31:0] w_sys_tmp3867;
	wire signed [31:0] w_sys_tmp3868;
	wire signed [31:0] w_sys_tmp3885;
	wire signed [31:0] w_sys_tmp3886;
	wire signed [31:0] w_sys_tmp3891;
	wire signed [31:0] w_sys_tmp3892;
	wire signed [31:0] w_sys_tmp3897;
	wire signed [31:0] w_sys_tmp3898;
	wire signed [31:0] w_sys_tmp3903;
	wire signed [31:0] w_sys_tmp3904;
	wire signed [31:0] w_sys_tmp3909;
	wire signed [31:0] w_sys_tmp3910;
	wire signed [31:0] w_sys_tmp3914;
	wire signed [31:0] w_sys_tmp3915;
	wire               w_sys_tmp3916;
	wire               w_sys_tmp3917;
	wire signed [31:0] w_sys_tmp3918;
	wire signed [31:0] w_sys_tmp3921;
	wire signed [31:0] w_sys_tmp3922;
	wire        [31:0] w_sys_tmp3923;
	wire signed [31:0] w_sys_tmp3927;
	wire signed [31:0] w_sys_tmp3928;
	wire signed [31:0] w_sys_tmp3933;
	wire signed [31:0] w_sys_tmp3934;
	wire signed [31:0] w_sys_tmp3939;
	wire signed [31:0] w_sys_tmp3940;
	wire signed [31:0] w_sys_tmp3945;
	wire signed [31:0] w_sys_tmp3946;
	wire signed [31:0] w_sys_tmp3951;
	wire signed [31:0] w_sys_tmp3952;
	wire signed [31:0] w_sys_tmp3957;
	wire signed [31:0] w_sys_tmp3958;
	wire signed [31:0] w_sys_tmp3962;
	wire signed [31:0] w_sys_tmp3963;
	wire signed [31:0] w_sys_tmp3967;
	wire signed [31:0] w_sys_tmp3968;
	wire signed [31:0] w_sys_tmp3972;
	wire signed [31:0] w_sys_tmp3973;
	wire signed [31:0] w_sys_tmp3977;
	wire signed [31:0] w_sys_tmp3978;
	wire signed [31:0] w_sys_tmp3982;
	wire signed [31:0] w_sys_tmp3983;
	wire signed [31:0] w_sys_tmp3987;
	wire signed [31:0] w_sys_tmp3988;
	wire signed [31:0] w_sys_tmp3992;
	wire signed [31:0] w_sys_tmp3993;
	wire signed [31:0] w_sys_tmp3997;
	wire signed [31:0] w_sys_tmp3998;
	wire signed [31:0] w_sys_tmp4002;
	wire signed [31:0] w_sys_tmp4003;
	wire signed [31:0] w_sys_tmp4007;
	wire signed [31:0] w_sys_tmp4008;
	wire signed [31:0] w_sys_tmp4012;
	wire signed [31:0] w_sys_tmp4013;
	wire signed [31:0] w_sys_tmp4017;
	wire signed [31:0] w_sys_tmp4018;
	wire signed [31:0] w_sys_tmp4022;
	wire signed [31:0] w_sys_tmp4023;
	wire signed [31:0] w_sys_tmp4027;
	wire signed [31:0] w_sys_tmp4028;
	wire signed [31:0] w_sys_tmp4032;
	wire signed [31:0] w_sys_tmp4033;
	wire signed [31:0] w_sys_tmp4037;
	wire signed [31:0] w_sys_tmp4038;
	wire signed [31:0] w_sys_tmp4042;
	wire signed [31:0] w_sys_tmp4043;
	wire signed [31:0] w_sys_tmp4047;
	wire signed [31:0] w_sys_tmp4048;
	wire signed [31:0] w_sys_tmp4052;
	wire signed [31:0] w_sys_tmp4053;
	wire signed [31:0] w_sys_tmp4057;
	wire signed [31:0] w_sys_tmp4058;
	wire signed [31:0] w_sys_tmp4062;
	wire signed [31:0] w_sys_tmp4063;
	wire signed [31:0] w_sys_tmp4067;
	wire signed [31:0] w_sys_tmp4068;
	wire signed [31:0] w_sys_tmp4072;
	wire signed [31:0] w_sys_tmp4073;
	wire signed [31:0] w_sys_tmp4077;
	wire signed [31:0] w_sys_tmp4078;
	wire signed [31:0] w_sys_tmp4082;
	wire signed [31:0] w_sys_tmp4083;
	wire signed [31:0] w_sys_tmp4087;
	wire signed [31:0] w_sys_tmp4088;
	wire signed [31:0] w_sys_tmp4092;
	wire signed [31:0] w_sys_tmp4093;
	wire signed [31:0] w_sys_tmp4097;
	wire signed [31:0] w_sys_tmp4098;
	wire signed [31:0] w_sys_tmp4102;
	wire signed [31:0] w_sys_tmp4103;
	wire signed [31:0] w_sys_tmp4107;
	wire signed [31:0] w_sys_tmp4108;
	wire signed [31:0] w_sys_tmp4112;
	wire signed [31:0] w_sys_tmp4113;
	wire signed [31:0] w_sys_tmp4117;
	wire signed [31:0] w_sys_tmp4118;
	wire signed [31:0] w_sys_tmp4122;
	wire signed [31:0] w_sys_tmp4123;
	wire signed [31:0] w_sys_tmp4127;
	wire signed [31:0] w_sys_tmp4128;
	wire signed [31:0] w_sys_tmp4132;
	wire signed [31:0] w_sys_tmp4133;
	wire signed [31:0] w_sys_tmp4137;
	wire signed [31:0] w_sys_tmp4138;
	wire signed [31:0] w_sys_tmp4142;
	wire signed [31:0] w_sys_tmp4143;
	wire signed [31:0] w_sys_tmp4147;
	wire signed [31:0] w_sys_tmp4148;
	wire signed [31:0] w_sys_tmp4152;
	wire signed [31:0] w_sys_tmp4153;
	wire signed [31:0] w_sys_tmp4157;
	wire signed [31:0] w_sys_tmp4158;
	wire signed [31:0] w_sys_tmp4162;
	wire signed [31:0] w_sys_tmp4163;
	wire signed [31:0] w_sys_tmp4167;
	wire signed [31:0] w_sys_tmp4168;
	wire signed [31:0] w_sys_tmp4172;
	wire signed [31:0] w_sys_tmp4173;
	wire signed [31:0] w_sys_tmp4177;
	wire signed [31:0] w_sys_tmp4178;
	wire signed [31:0] w_sys_tmp4182;
	wire signed [31:0] w_sys_tmp4183;
	wire signed [31:0] w_sys_tmp4187;
	wire signed [31:0] w_sys_tmp4188;
	wire signed [31:0] w_sys_tmp4192;
	wire signed [31:0] w_sys_tmp4193;
	wire signed [31:0] w_sys_tmp4197;
	wire signed [31:0] w_sys_tmp4198;
	wire signed [31:0] w_sys_tmp4202;
	wire signed [31:0] w_sys_tmp4203;
	wire signed [31:0] w_sys_tmp4207;
	wire signed [31:0] w_sys_tmp4208;
	wire signed [31:0] w_sys_tmp4212;
	wire signed [31:0] w_sys_tmp4213;
	wire signed [31:0] w_sys_tmp4217;
	wire signed [31:0] w_sys_tmp4218;
	wire signed [31:0] w_sys_tmp4222;
	wire signed [31:0] w_sys_tmp4223;
	wire signed [31:0] w_sys_tmp4227;
	wire signed [31:0] w_sys_tmp4228;
	wire signed [31:0] w_sys_tmp4232;
	wire signed [31:0] w_sys_tmp4233;
	wire signed [31:0] w_sys_tmp4237;
	wire signed [31:0] w_sys_tmp4238;
	wire signed [31:0] w_sys_tmp4242;
	wire signed [31:0] w_sys_tmp4243;
	wire signed [31:0] w_sys_tmp4247;
	wire signed [31:0] w_sys_tmp4248;
	wire signed [31:0] w_sys_tmp4252;
	wire signed [31:0] w_sys_tmp4253;
	wire signed [31:0] w_sys_tmp4257;
	wire signed [31:0] w_sys_tmp4258;
	wire signed [31:0] w_sys_tmp4262;
	wire signed [31:0] w_sys_tmp4263;
	wire signed [31:0] w_sys_tmp4267;
	wire signed [31:0] w_sys_tmp4268;
	wire signed [31:0] w_sys_tmp4272;
	wire signed [31:0] w_sys_tmp4273;
	wire signed [31:0] w_sys_tmp4277;
	wire signed [31:0] w_sys_tmp4278;
	wire signed [31:0] w_sys_tmp4282;
	wire signed [31:0] w_sys_tmp4283;
	wire signed [31:0] w_sys_tmp4287;
	wire signed [31:0] w_sys_tmp4288;
	wire signed [31:0] w_sys_tmp4292;
	wire signed [31:0] w_sys_tmp4293;
	wire signed [31:0] w_sys_tmp4297;
	wire signed [31:0] w_sys_tmp4298;
	wire signed [31:0] w_sys_tmp4302;
	wire signed [31:0] w_sys_tmp4303;
	wire signed [31:0] w_sys_tmp4307;
	wire signed [31:0] w_sys_tmp4308;
	wire signed [31:0] w_sys_tmp4312;
	wire signed [31:0] w_sys_tmp4313;
	wire signed [31:0] w_sys_tmp4317;
	wire signed [31:0] w_sys_tmp4318;
	wire signed [31:0] w_sys_tmp4322;
	wire signed [31:0] w_sys_tmp4323;
	wire signed [31:0] w_sys_tmp4327;
	wire signed [31:0] w_sys_tmp4328;
	wire signed [31:0] w_sys_tmp4332;
	wire signed [31:0] w_sys_tmp4333;
	wire signed [31:0] w_sys_tmp4337;
	wire signed [31:0] w_sys_tmp4338;
	wire signed [31:0] w_sys_tmp4342;
	wire signed [31:0] w_sys_tmp4343;
	wire signed [31:0] w_sys_tmp4347;
	wire signed [31:0] w_sys_tmp4348;
	wire signed [31:0] w_sys_tmp4352;
	wire signed [31:0] w_sys_tmp4353;
	wire signed [31:0] w_sys_tmp4357;
	wire signed [31:0] w_sys_tmp4358;
	wire signed [31:0] w_sys_tmp4362;
	wire signed [31:0] w_sys_tmp4363;
	wire signed [31:0] w_sys_tmp4367;
	wire signed [31:0] w_sys_tmp4368;
	wire signed [31:0] w_sys_tmp4372;
	wire signed [31:0] w_sys_tmp4373;
	wire signed [31:0] w_sys_tmp4377;
	wire signed [31:0] w_sys_tmp4378;
	wire signed [31:0] w_sys_tmp4382;
	wire signed [31:0] w_sys_tmp4383;
	wire signed [31:0] w_sys_tmp4387;
	wire signed [31:0] w_sys_tmp4388;
	wire signed [31:0] w_sys_tmp4392;
	wire signed [31:0] w_sys_tmp4393;
	wire signed [31:0] w_sys_tmp4397;
	wire signed [31:0] w_sys_tmp4398;
	wire signed [31:0] w_sys_tmp4402;
	wire signed [31:0] w_sys_tmp4403;
	wire signed [31:0] w_sys_tmp4407;
	wire signed [31:0] w_sys_tmp4408;
	wire signed [31:0] w_sys_tmp4412;
	wire signed [31:0] w_sys_tmp4413;
	wire signed [31:0] w_sys_tmp4417;
	wire signed [31:0] w_sys_tmp4418;
	wire signed [31:0] w_sys_tmp4422;
	wire signed [31:0] w_sys_tmp4423;
	wire signed [31:0] w_sys_tmp4427;
	wire signed [31:0] w_sys_tmp4428;
	wire signed [31:0] w_sys_tmp4432;
	wire signed [31:0] w_sys_tmp4433;
	wire signed [31:0] w_sys_tmp4437;
	wire signed [31:0] w_sys_tmp4438;
	wire signed [31:0] w_sys_tmp4442;
	wire signed [31:0] w_sys_tmp4443;
	wire signed [31:0] w_sys_tmp4447;
	wire signed [31:0] w_sys_tmp4448;
	wire signed [31:0] w_sys_tmp4452;
	wire signed [31:0] w_sys_tmp4453;
	wire signed [31:0] w_sys_tmp4457;
	wire signed [31:0] w_sys_tmp4458;
	wire signed [31:0] w_sys_tmp4462;
	wire signed [31:0] w_sys_tmp4463;
	wire signed [31:0] w_sys_tmp4467;
	wire signed [31:0] w_sys_tmp4468;
	wire signed [31:0] w_sys_tmp4472;
	wire signed [31:0] w_sys_tmp4473;
	wire signed [31:0] w_sys_tmp4477;
	wire signed [31:0] w_sys_tmp4478;
	wire signed [31:0] w_sys_tmp4482;
	wire signed [31:0] w_sys_tmp4483;
	wire signed [31:0] w_sys_tmp4487;
	wire signed [31:0] w_sys_tmp4488;
	wire signed [31:0] w_sys_tmp4492;
	wire signed [31:0] w_sys_tmp4493;
	wire signed [31:0] w_sys_tmp4497;
	wire signed [31:0] w_sys_tmp4498;
	wire signed [31:0] w_sys_tmp4502;
	wire signed [31:0] w_sys_tmp4503;
	wire signed [31:0] w_sys_tmp4506;
	wire signed [31:0] w_sys_tmp4507;
	wire               w_sys_tmp4508;
	wire               w_sys_tmp4509;
	wire signed [31:0] w_sys_tmp4510;
	wire signed [31:0] w_sys_tmp4513;
	wire signed [31:0] w_sys_tmp4514;
	wire        [31:0] w_sys_tmp4515;
	wire signed [31:0] w_sys_tmp4519;
	wire signed [31:0] w_sys_tmp4520;
	wire signed [31:0] w_sys_tmp4525;
	wire signed [31:0] w_sys_tmp4526;
	wire signed [31:0] w_sys_tmp4531;
	wire signed [31:0] w_sys_tmp4532;
	wire signed [31:0] w_sys_tmp4537;
	wire signed [31:0] w_sys_tmp4538;
	wire signed [31:0] w_sys_tmp4543;
	wire signed [31:0] w_sys_tmp4544;
	wire signed [31:0] w_sys_tmp4549;
	wire signed [31:0] w_sys_tmp4550;
	wire signed [31:0] w_sys_tmp4554;
	wire signed [31:0] w_sys_tmp4555;
	wire signed [31:0] w_sys_tmp4559;
	wire signed [31:0] w_sys_tmp4560;
	wire signed [31:0] w_sys_tmp4564;
	wire signed [31:0] w_sys_tmp4565;
	wire signed [31:0] w_sys_tmp4569;
	wire signed [31:0] w_sys_tmp4570;
	wire signed [31:0] w_sys_tmp4574;
	wire signed [31:0] w_sys_tmp4575;
	wire signed [31:0] w_sys_tmp4579;
	wire signed [31:0] w_sys_tmp4580;
	wire signed [31:0] w_sys_tmp4584;
	wire signed [31:0] w_sys_tmp4585;
	wire signed [31:0] w_sys_tmp4589;
	wire signed [31:0] w_sys_tmp4590;
	wire signed [31:0] w_sys_tmp4594;
	wire signed [31:0] w_sys_tmp4595;
	wire signed [31:0] w_sys_tmp4599;
	wire signed [31:0] w_sys_tmp4600;
	wire signed [31:0] w_sys_tmp4604;
	wire signed [31:0] w_sys_tmp4605;
	wire signed [31:0] w_sys_tmp4609;
	wire signed [31:0] w_sys_tmp4610;
	wire signed [31:0] w_sys_tmp4614;
	wire signed [31:0] w_sys_tmp4615;
	wire signed [31:0] w_sys_tmp4619;
	wire signed [31:0] w_sys_tmp4620;
	wire signed [31:0] w_sys_tmp4624;
	wire signed [31:0] w_sys_tmp4625;
	wire signed [31:0] w_sys_tmp4629;
	wire signed [31:0] w_sys_tmp4630;
	wire signed [31:0] w_sys_tmp4634;
	wire signed [31:0] w_sys_tmp4635;
	wire signed [31:0] w_sys_tmp4639;
	wire signed [31:0] w_sys_tmp4640;
	wire signed [31:0] w_sys_tmp4644;
	wire signed [31:0] w_sys_tmp4645;
	wire signed [31:0] w_sys_tmp4649;
	wire signed [31:0] w_sys_tmp4650;
	wire signed [31:0] w_sys_tmp4654;
	wire signed [31:0] w_sys_tmp4655;
	wire signed [31:0] w_sys_tmp4659;
	wire signed [31:0] w_sys_tmp4660;
	wire signed [31:0] w_sys_tmp4663;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 5'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 8'h1);
	assign w_fld_T_0_addr_0 = 10'sh0;
	assign w_fld_T_0_datain_0 = 32'h0;
	assign w_fld_T_0_r_w_0 = 1'h0;
	assign w_fld_T_0_ce_0 = w_sys_ce;
	assign w_fld_T_0_ce_1 = w_sys_ce;
	assign w_fld_TT_1_addr_0 = 10'sh0;
	assign w_fld_TT_1_datain_0 = 32'h0;
	assign w_fld_TT_1_r_w_0 = 1'h0;
	assign w_fld_TT_1_ce_0 = w_sys_ce;
	assign w_fld_TT_1_ce_1 = w_sys_ce;
	assign w_fld_U_2_addr_0 = 10'sh0;
	assign w_fld_U_2_datain_0 = 32'h0;
	assign w_fld_U_2_r_w_0 = 1'h0;
	assign w_fld_U_2_ce_0 = w_sys_ce;
	assign w_fld_U_2_ce_1 = w_sys_ce;
	assign w_fld_V_3_addr_0 = 10'sh0;
	assign w_fld_V_3_datain_0 = 32'h0;
	assign w_fld_V_3_r_w_0 = 1'h0;
	assign w_fld_V_3_ce_0 = w_sys_ce;
	assign w_fld_V_3_ce_1 = w_sys_ce;
	assign w_sub19_T_addr = ( (|r_sys_processing_methodID) ? r_sub19_T_addr : 10'sh0 ) ;
	assign w_sub19_T_datain = ( (|r_sys_processing_methodID) ? r_sub19_T_datain : 32'h0 ) ;
	assign w_sub19_T_r_w = ( (|r_sys_processing_methodID) ? r_sub19_T_r_w : 1'h0 ) ;
	assign w_sub19_V_addr = ( (|r_sys_processing_methodID) ? r_sub19_V_addr : 10'sh0 ) ;
	assign w_sub19_V_datain = ( (|r_sys_processing_methodID) ? r_sub19_V_datain : 32'h0 ) ;
	assign w_sub19_V_r_w = ( (|r_sys_processing_methodID) ? r_sub19_V_r_w : 1'h0 ) ;
	assign w_sub19_U_addr = ( (|r_sys_processing_methodID) ? r_sub19_U_addr : 10'sh0 ) ;
	assign w_sub19_U_datain = ( (|r_sys_processing_methodID) ? r_sub19_U_datain : 32'h0 ) ;
	assign w_sub19_U_r_w = ( (|r_sys_processing_methodID) ? r_sub19_U_r_w : 1'h0 ) ;
	assign w_sub19_result_addr = ( (|r_sys_processing_methodID) ? r_sub19_result_addr : 10'sh0 ) ;
	assign w_sub19_result_datain = ( (|r_sys_processing_methodID) ? r_sub19_result_datain : 32'h0 ) ;
	assign w_sub19_result_r_w = ( (|r_sys_processing_methodID) ? r_sub19_result_r_w : 1'h0 ) ;
	assign w_sub09_T_addr = ( (|r_sys_processing_methodID) ? r_sub09_T_addr : 10'sh0 ) ;
	assign w_sub09_T_datain = ( (|r_sys_processing_methodID) ? r_sub09_T_datain : 32'h0 ) ;
	assign w_sub09_T_r_w = ( (|r_sys_processing_methodID) ? r_sub09_T_r_w : 1'h0 ) ;
	assign w_sub09_V_addr = ( (|r_sys_processing_methodID) ? r_sub09_V_addr : 10'sh0 ) ;
	assign w_sub09_V_datain = ( (|r_sys_processing_methodID) ? r_sub09_V_datain : 32'h0 ) ;
	assign w_sub09_V_r_w = ( (|r_sys_processing_methodID) ? r_sub09_V_r_w : 1'h0 ) ;
	assign w_sub09_U_addr = ( (|r_sys_processing_methodID) ? r_sub09_U_addr : 10'sh0 ) ;
	assign w_sub09_U_datain = ( (|r_sys_processing_methodID) ? r_sub09_U_datain : 32'h0 ) ;
	assign w_sub09_U_r_w = ( (|r_sys_processing_methodID) ? r_sub09_U_r_w : 1'h0 ) ;
	assign w_sub09_result_addr = ( (|r_sys_processing_methodID) ? r_sub09_result_addr : 10'sh0 ) ;
	assign w_sub09_result_datain = ( (|r_sys_processing_methodID) ? r_sub09_result_datain : 32'h0 ) ;
	assign w_sub09_result_r_w = ( (|r_sys_processing_methodID) ? r_sub09_result_r_w : 1'h0 ) ;
	assign w_sub08_T_addr = ( (|r_sys_processing_methodID) ? r_sub08_T_addr : 10'sh0 ) ;
	assign w_sub08_T_datain = ( (|r_sys_processing_methodID) ? r_sub08_T_datain : 32'h0 ) ;
	assign w_sub08_T_r_w = ( (|r_sys_processing_methodID) ? r_sub08_T_r_w : 1'h0 ) ;
	assign w_sub08_V_addr = ( (|r_sys_processing_methodID) ? r_sub08_V_addr : 10'sh0 ) ;
	assign w_sub08_V_datain = ( (|r_sys_processing_methodID) ? r_sub08_V_datain : 32'h0 ) ;
	assign w_sub08_V_r_w = ( (|r_sys_processing_methodID) ? r_sub08_V_r_w : 1'h0 ) ;
	assign w_sub08_U_addr = ( (|r_sys_processing_methodID) ? r_sub08_U_addr : 10'sh0 ) ;
	assign w_sub08_U_datain = ( (|r_sys_processing_methodID) ? r_sub08_U_datain : 32'h0 ) ;
	assign w_sub08_U_r_w = ( (|r_sys_processing_methodID) ? r_sub08_U_r_w : 1'h0 ) ;
	assign w_sub08_result_addr = ( (|r_sys_processing_methodID) ? r_sub08_result_addr : 10'sh0 ) ;
	assign w_sub08_result_datain = ( (|r_sys_processing_methodID) ? r_sub08_result_datain : 32'h0 ) ;
	assign w_sub08_result_r_w = ( (|r_sys_processing_methodID) ? r_sub08_result_r_w : 1'h0 ) ;
	assign w_sub24_T_addr = ( (|r_sys_processing_methodID) ? r_sub24_T_addr : 10'sh0 ) ;
	assign w_sub24_T_datain = ( (|r_sys_processing_methodID) ? r_sub24_T_datain : 32'h0 ) ;
	assign w_sub24_T_r_w = ( (|r_sys_processing_methodID) ? r_sub24_T_r_w : 1'h0 ) ;
	assign w_sub24_V_addr = ( (|r_sys_processing_methodID) ? r_sub24_V_addr : 10'sh0 ) ;
	assign w_sub24_V_datain = ( (|r_sys_processing_methodID) ? r_sub24_V_datain : 32'h0 ) ;
	assign w_sub24_V_r_w = ( (|r_sys_processing_methodID) ? r_sub24_V_r_w : 1'h0 ) ;
	assign w_sub24_U_addr = ( (|r_sys_processing_methodID) ? r_sub24_U_addr : 10'sh0 ) ;
	assign w_sub24_U_datain = ( (|r_sys_processing_methodID) ? r_sub24_U_datain : 32'h0 ) ;
	assign w_sub24_U_r_w = ( (|r_sys_processing_methodID) ? r_sub24_U_r_w : 1'h0 ) ;
	assign w_sub24_result_addr = ( (|r_sys_processing_methodID) ? r_sub24_result_addr : 10'sh0 ) ;
	assign w_sub24_result_datain = ( (|r_sys_processing_methodID) ? r_sub24_result_datain : 32'h0 ) ;
	assign w_sub24_result_r_w = ( (|r_sys_processing_methodID) ? r_sub24_result_r_w : 1'h0 ) ;
	assign w_sub22_T_addr = ( (|r_sys_processing_methodID) ? r_sub22_T_addr : 10'sh0 ) ;
	assign w_sub22_T_datain = ( (|r_sys_processing_methodID) ? r_sub22_T_datain : 32'h0 ) ;
	assign w_sub22_T_r_w = ( (|r_sys_processing_methodID) ? r_sub22_T_r_w : 1'h0 ) ;
	assign w_sub22_V_addr = ( (|r_sys_processing_methodID) ? r_sub22_V_addr : 10'sh0 ) ;
	assign w_sub22_V_datain = ( (|r_sys_processing_methodID) ? r_sub22_V_datain : 32'h0 ) ;
	assign w_sub22_V_r_w = ( (|r_sys_processing_methodID) ? r_sub22_V_r_w : 1'h0 ) ;
	assign w_sub22_U_addr = ( (|r_sys_processing_methodID) ? r_sub22_U_addr : 10'sh0 ) ;
	assign w_sub22_U_datain = ( (|r_sys_processing_methodID) ? r_sub22_U_datain : 32'h0 ) ;
	assign w_sub22_U_r_w = ( (|r_sys_processing_methodID) ? r_sub22_U_r_w : 1'h0 ) ;
	assign w_sub22_result_addr = ( (|r_sys_processing_methodID) ? r_sub22_result_addr : 10'sh0 ) ;
	assign w_sub22_result_datain = ( (|r_sys_processing_methodID) ? r_sub22_result_datain : 32'h0 ) ;
	assign w_sub22_result_r_w = ( (|r_sys_processing_methodID) ? r_sub22_result_r_w : 1'h0 ) ;
	assign w_sub23_T_addr = ( (|r_sys_processing_methodID) ? r_sub23_T_addr : 10'sh0 ) ;
	assign w_sub23_T_datain = ( (|r_sys_processing_methodID) ? r_sub23_T_datain : 32'h0 ) ;
	assign w_sub23_T_r_w = ( (|r_sys_processing_methodID) ? r_sub23_T_r_w : 1'h0 ) ;
	assign w_sub23_V_addr = ( (|r_sys_processing_methodID) ? r_sub23_V_addr : 10'sh0 ) ;
	assign w_sub23_V_datain = ( (|r_sys_processing_methodID) ? r_sub23_V_datain : 32'h0 ) ;
	assign w_sub23_V_r_w = ( (|r_sys_processing_methodID) ? r_sub23_V_r_w : 1'h0 ) ;
	assign w_sub23_U_addr = ( (|r_sys_processing_methodID) ? r_sub23_U_addr : 10'sh0 ) ;
	assign w_sub23_U_datain = ( (|r_sys_processing_methodID) ? r_sub23_U_datain : 32'h0 ) ;
	assign w_sub23_U_r_w = ( (|r_sys_processing_methodID) ? r_sub23_U_r_w : 1'h0 ) ;
	assign w_sub23_result_addr = ( (|r_sys_processing_methodID) ? r_sub23_result_addr : 10'sh0 ) ;
	assign w_sub23_result_datain = ( (|r_sys_processing_methodID) ? r_sub23_result_datain : 32'h0 ) ;
	assign w_sub23_result_r_w = ( (|r_sys_processing_methodID) ? r_sub23_result_r_w : 1'h0 ) ;
	assign w_sub12_T_addr = ( (|r_sys_processing_methodID) ? r_sub12_T_addr : 10'sh0 ) ;
	assign w_sub12_T_datain = ( (|r_sys_processing_methodID) ? r_sub12_T_datain : 32'h0 ) ;
	assign w_sub12_T_r_w = ( (|r_sys_processing_methodID) ? r_sub12_T_r_w : 1'h0 ) ;
	assign w_sub12_V_addr = ( (|r_sys_processing_methodID) ? r_sub12_V_addr : 10'sh0 ) ;
	assign w_sub12_V_datain = ( (|r_sys_processing_methodID) ? r_sub12_V_datain : 32'h0 ) ;
	assign w_sub12_V_r_w = ( (|r_sys_processing_methodID) ? r_sub12_V_r_w : 1'h0 ) ;
	assign w_sub12_U_addr = ( (|r_sys_processing_methodID) ? r_sub12_U_addr : 10'sh0 ) ;
	assign w_sub12_U_datain = ( (|r_sys_processing_methodID) ? r_sub12_U_datain : 32'h0 ) ;
	assign w_sub12_U_r_w = ( (|r_sys_processing_methodID) ? r_sub12_U_r_w : 1'h0 ) ;
	assign w_sub12_result_addr = ( (|r_sys_processing_methodID) ? r_sub12_result_addr : 10'sh0 ) ;
	assign w_sub12_result_datain = ( (|r_sys_processing_methodID) ? r_sub12_result_datain : 32'h0 ) ;
	assign w_sub12_result_r_w = ( (|r_sys_processing_methodID) ? r_sub12_result_r_w : 1'h0 ) ;
	assign w_sub03_T_addr = ( (|r_sys_processing_methodID) ? r_sub03_T_addr : 10'sh0 ) ;
	assign w_sub03_T_datain = ( (|r_sys_processing_methodID) ? r_sub03_T_datain : 32'h0 ) ;
	assign w_sub03_T_r_w = ( (|r_sys_processing_methodID) ? r_sub03_T_r_w : 1'h0 ) ;
	assign w_sub03_V_addr = ( (|r_sys_processing_methodID) ? r_sub03_V_addr : 10'sh0 ) ;
	assign w_sub03_V_datain = ( (|r_sys_processing_methodID) ? r_sub03_V_datain : 32'h0 ) ;
	assign w_sub03_V_r_w = ( (|r_sys_processing_methodID) ? r_sub03_V_r_w : 1'h0 ) ;
	assign w_sub03_U_addr = ( (|r_sys_processing_methodID) ? r_sub03_U_addr : 10'sh0 ) ;
	assign w_sub03_U_datain = ( (|r_sys_processing_methodID) ? r_sub03_U_datain : 32'h0 ) ;
	assign w_sub03_U_r_w = ( (|r_sys_processing_methodID) ? r_sub03_U_r_w : 1'h0 ) ;
	assign w_sub03_result_addr = ( (|r_sys_processing_methodID) ? r_sub03_result_addr : 10'sh0 ) ;
	assign w_sub03_result_datain = ( (|r_sys_processing_methodID) ? r_sub03_result_datain : 32'h0 ) ;
	assign w_sub03_result_r_w = ( (|r_sys_processing_methodID) ? r_sub03_result_r_w : 1'h0 ) ;
	assign w_sub02_T_addr = ( (|r_sys_processing_methodID) ? r_sub02_T_addr : 10'sh0 ) ;
	assign w_sub02_T_datain = ( (|r_sys_processing_methodID) ? r_sub02_T_datain : 32'h0 ) ;
	assign w_sub02_T_r_w = ( (|r_sys_processing_methodID) ? r_sub02_T_r_w : 1'h0 ) ;
	assign w_sub02_V_addr = ( (|r_sys_processing_methodID) ? r_sub02_V_addr : 10'sh0 ) ;
	assign w_sub02_V_datain = ( (|r_sys_processing_methodID) ? r_sub02_V_datain : 32'h0 ) ;
	assign w_sub02_V_r_w = ( (|r_sys_processing_methodID) ? r_sub02_V_r_w : 1'h0 ) ;
	assign w_sub02_U_addr = ( (|r_sys_processing_methodID) ? r_sub02_U_addr : 10'sh0 ) ;
	assign w_sub02_U_datain = ( (|r_sys_processing_methodID) ? r_sub02_U_datain : 32'h0 ) ;
	assign w_sub02_U_r_w = ( (|r_sys_processing_methodID) ? r_sub02_U_r_w : 1'h0 ) ;
	assign w_sub02_result_addr = ( (|r_sys_processing_methodID) ? r_sub02_result_addr : 10'sh0 ) ;
	assign w_sub02_result_datain = ( (|r_sys_processing_methodID) ? r_sub02_result_datain : 32'h0 ) ;
	assign w_sub02_result_r_w = ( (|r_sys_processing_methodID) ? r_sub02_result_r_w : 1'h0 ) ;
	assign w_sub11_T_addr = ( (|r_sys_processing_methodID) ? r_sub11_T_addr : 10'sh0 ) ;
	assign w_sub11_T_datain = ( (|r_sys_processing_methodID) ? r_sub11_T_datain : 32'h0 ) ;
	assign w_sub11_T_r_w = ( (|r_sys_processing_methodID) ? r_sub11_T_r_w : 1'h0 ) ;
	assign w_sub11_V_addr = ( (|r_sys_processing_methodID) ? r_sub11_V_addr : 10'sh0 ) ;
	assign w_sub11_V_datain = ( (|r_sys_processing_methodID) ? r_sub11_V_datain : 32'h0 ) ;
	assign w_sub11_V_r_w = ( (|r_sys_processing_methodID) ? r_sub11_V_r_w : 1'h0 ) ;
	assign w_sub11_U_addr = ( (|r_sys_processing_methodID) ? r_sub11_U_addr : 10'sh0 ) ;
	assign w_sub11_U_datain = ( (|r_sys_processing_methodID) ? r_sub11_U_datain : 32'h0 ) ;
	assign w_sub11_U_r_w = ( (|r_sys_processing_methodID) ? r_sub11_U_r_w : 1'h0 ) ;
	assign w_sub11_result_addr = ( (|r_sys_processing_methodID) ? r_sub11_result_addr : 10'sh0 ) ;
	assign w_sub11_result_datain = ( (|r_sys_processing_methodID) ? r_sub11_result_datain : 32'h0 ) ;
	assign w_sub11_result_r_w = ( (|r_sys_processing_methodID) ? r_sub11_result_r_w : 1'h0 ) ;
	assign w_sub14_T_addr = ( (|r_sys_processing_methodID) ? r_sub14_T_addr : 10'sh0 ) ;
	assign w_sub14_T_datain = ( (|r_sys_processing_methodID) ? r_sub14_T_datain : 32'h0 ) ;
	assign w_sub14_T_r_w = ( (|r_sys_processing_methodID) ? r_sub14_T_r_w : 1'h0 ) ;
	assign w_sub14_V_addr = ( (|r_sys_processing_methodID) ? r_sub14_V_addr : 10'sh0 ) ;
	assign w_sub14_V_datain = ( (|r_sys_processing_methodID) ? r_sub14_V_datain : 32'h0 ) ;
	assign w_sub14_V_r_w = ( (|r_sys_processing_methodID) ? r_sub14_V_r_w : 1'h0 ) ;
	assign w_sub14_U_addr = ( (|r_sys_processing_methodID) ? r_sub14_U_addr : 10'sh0 ) ;
	assign w_sub14_U_datain = ( (|r_sys_processing_methodID) ? r_sub14_U_datain : 32'h0 ) ;
	assign w_sub14_U_r_w = ( (|r_sys_processing_methodID) ? r_sub14_U_r_w : 1'h0 ) ;
	assign w_sub14_result_addr = ( (|r_sys_processing_methodID) ? r_sub14_result_addr : 10'sh0 ) ;
	assign w_sub14_result_datain = ( (|r_sys_processing_methodID) ? r_sub14_result_datain : 32'h0 ) ;
	assign w_sub14_result_r_w = ( (|r_sys_processing_methodID) ? r_sub14_result_r_w : 1'h0 ) ;
	assign w_sub01_T_addr = ( (|r_sys_processing_methodID) ? r_sub01_T_addr : 10'sh0 ) ;
	assign w_sub01_T_datain = ( (|r_sys_processing_methodID) ? r_sub01_T_datain : 32'h0 ) ;
	assign w_sub01_T_r_w = ( (|r_sys_processing_methodID) ? r_sub01_T_r_w : 1'h0 ) ;
	assign w_sub01_V_addr = ( (|r_sys_processing_methodID) ? r_sub01_V_addr : 10'sh0 ) ;
	assign w_sub01_V_datain = ( (|r_sys_processing_methodID) ? r_sub01_V_datain : 32'h0 ) ;
	assign w_sub01_V_r_w = ( (|r_sys_processing_methodID) ? r_sub01_V_r_w : 1'h0 ) ;
	assign w_sub01_U_addr = ( (|r_sys_processing_methodID) ? r_sub01_U_addr : 10'sh0 ) ;
	assign w_sub01_U_datain = ( (|r_sys_processing_methodID) ? r_sub01_U_datain : 32'h0 ) ;
	assign w_sub01_U_r_w = ( (|r_sys_processing_methodID) ? r_sub01_U_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 10'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub00_T_addr = ( (|r_sys_processing_methodID) ? r_sub00_T_addr : 10'sh0 ) ;
	assign w_sub00_T_datain = ( (|r_sys_processing_methodID) ? r_sub00_T_datain : 32'h0 ) ;
	assign w_sub00_T_r_w = ( (|r_sys_processing_methodID) ? r_sub00_T_r_w : 1'h0 ) ;
	assign w_sub00_V_addr = ( (|r_sys_processing_methodID) ? r_sub00_V_addr : 10'sh0 ) ;
	assign w_sub00_V_datain = ( (|r_sys_processing_methodID) ? r_sub00_V_datain : 32'h0 ) ;
	assign w_sub00_V_r_w = ( (|r_sys_processing_methodID) ? r_sub00_V_r_w : 1'h0 ) ;
	assign w_sub00_U_addr = ( (|r_sys_processing_methodID) ? r_sub00_U_addr : 10'sh0 ) ;
	assign w_sub00_U_datain = ( (|r_sys_processing_methodID) ? r_sub00_U_datain : 32'h0 ) ;
	assign w_sub00_U_r_w = ( (|r_sys_processing_methodID) ? r_sub00_U_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 10'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sub13_T_addr = ( (|r_sys_processing_methodID) ? r_sub13_T_addr : 10'sh0 ) ;
	assign w_sub13_T_datain = ( (|r_sys_processing_methodID) ? r_sub13_T_datain : 32'h0 ) ;
	assign w_sub13_T_r_w = ( (|r_sys_processing_methodID) ? r_sub13_T_r_w : 1'h0 ) ;
	assign w_sub13_V_addr = ( (|r_sys_processing_methodID) ? r_sub13_V_addr : 10'sh0 ) ;
	assign w_sub13_V_datain = ( (|r_sys_processing_methodID) ? r_sub13_V_datain : 32'h0 ) ;
	assign w_sub13_V_r_w = ( (|r_sys_processing_methodID) ? r_sub13_V_r_w : 1'h0 ) ;
	assign w_sub13_U_addr = ( (|r_sys_processing_methodID) ? r_sub13_U_addr : 10'sh0 ) ;
	assign w_sub13_U_datain = ( (|r_sys_processing_methodID) ? r_sub13_U_datain : 32'h0 ) ;
	assign w_sub13_U_r_w = ( (|r_sys_processing_methodID) ? r_sub13_U_r_w : 1'h0 ) ;
	assign w_sub13_result_addr = ( (|r_sys_processing_methodID) ? r_sub13_result_addr : 10'sh0 ) ;
	assign w_sub13_result_datain = ( (|r_sys_processing_methodID) ? r_sub13_result_datain : 32'h0 ) ;
	assign w_sub13_result_r_w = ( (|r_sys_processing_methodID) ? r_sub13_result_r_w : 1'h0 ) ;
	assign w_sub07_T_addr = ( (|r_sys_processing_methodID) ? r_sub07_T_addr : 10'sh0 ) ;
	assign w_sub07_T_datain = ( (|r_sys_processing_methodID) ? r_sub07_T_datain : 32'h0 ) ;
	assign w_sub07_T_r_w = ( (|r_sys_processing_methodID) ? r_sub07_T_r_w : 1'h0 ) ;
	assign w_sub07_V_addr = ( (|r_sys_processing_methodID) ? r_sub07_V_addr : 10'sh0 ) ;
	assign w_sub07_V_datain = ( (|r_sys_processing_methodID) ? r_sub07_V_datain : 32'h0 ) ;
	assign w_sub07_V_r_w = ( (|r_sys_processing_methodID) ? r_sub07_V_r_w : 1'h0 ) ;
	assign w_sub07_U_addr = ( (|r_sys_processing_methodID) ? r_sub07_U_addr : 10'sh0 ) ;
	assign w_sub07_U_datain = ( (|r_sys_processing_methodID) ? r_sub07_U_datain : 32'h0 ) ;
	assign w_sub07_U_r_w = ( (|r_sys_processing_methodID) ? r_sub07_U_r_w : 1'h0 ) ;
	assign w_sub07_result_addr = ( (|r_sys_processing_methodID) ? r_sub07_result_addr : 10'sh0 ) ;
	assign w_sub07_result_datain = ( (|r_sys_processing_methodID) ? r_sub07_result_datain : 32'h0 ) ;
	assign w_sub07_result_r_w = ( (|r_sys_processing_methodID) ? r_sub07_result_r_w : 1'h0 ) ;
	assign w_sub16_T_addr = ( (|r_sys_processing_methodID) ? r_sub16_T_addr : 10'sh0 ) ;
	assign w_sub16_T_datain = ( (|r_sys_processing_methodID) ? r_sub16_T_datain : 32'h0 ) ;
	assign w_sub16_T_r_w = ( (|r_sys_processing_methodID) ? r_sub16_T_r_w : 1'h0 ) ;
	assign w_sub16_V_addr = ( (|r_sys_processing_methodID) ? r_sub16_V_addr : 10'sh0 ) ;
	assign w_sub16_V_datain = ( (|r_sys_processing_methodID) ? r_sub16_V_datain : 32'h0 ) ;
	assign w_sub16_V_r_w = ( (|r_sys_processing_methodID) ? r_sub16_V_r_w : 1'h0 ) ;
	assign w_sub16_U_addr = ( (|r_sys_processing_methodID) ? r_sub16_U_addr : 10'sh0 ) ;
	assign w_sub16_U_datain = ( (|r_sys_processing_methodID) ? r_sub16_U_datain : 32'h0 ) ;
	assign w_sub16_U_r_w = ( (|r_sys_processing_methodID) ? r_sub16_U_r_w : 1'h0 ) ;
	assign w_sub16_result_addr = ( (|r_sys_processing_methodID) ? r_sub16_result_addr : 10'sh0 ) ;
	assign w_sub16_result_datain = ( (|r_sys_processing_methodID) ? r_sub16_result_datain : 32'h0 ) ;
	assign w_sub16_result_r_w = ( (|r_sys_processing_methodID) ? r_sub16_result_r_w : 1'h0 ) ;
	assign w_sub06_T_addr = ( (|r_sys_processing_methodID) ? r_sub06_T_addr : 10'sh0 ) ;
	assign w_sub06_T_datain = ( (|r_sys_processing_methodID) ? r_sub06_T_datain : 32'h0 ) ;
	assign w_sub06_T_r_w = ( (|r_sys_processing_methodID) ? r_sub06_T_r_w : 1'h0 ) ;
	assign w_sub06_V_addr = ( (|r_sys_processing_methodID) ? r_sub06_V_addr : 10'sh0 ) ;
	assign w_sub06_V_datain = ( (|r_sys_processing_methodID) ? r_sub06_V_datain : 32'h0 ) ;
	assign w_sub06_V_r_w = ( (|r_sys_processing_methodID) ? r_sub06_V_r_w : 1'h0 ) ;
	assign w_sub06_U_addr = ( (|r_sys_processing_methodID) ? r_sub06_U_addr : 10'sh0 ) ;
	assign w_sub06_U_datain = ( (|r_sys_processing_methodID) ? r_sub06_U_datain : 32'h0 ) ;
	assign w_sub06_U_r_w = ( (|r_sys_processing_methodID) ? r_sub06_U_r_w : 1'h0 ) ;
	assign w_sub06_result_addr = ( (|r_sys_processing_methodID) ? r_sub06_result_addr : 10'sh0 ) ;
	assign w_sub06_result_datain = ( (|r_sys_processing_methodID) ? r_sub06_result_datain : 32'h0 ) ;
	assign w_sub06_result_r_w = ( (|r_sys_processing_methodID) ? r_sub06_result_r_w : 1'h0 ) ;
	assign w_sub15_T_addr = ( (|r_sys_processing_methodID) ? r_sub15_T_addr : 10'sh0 ) ;
	assign w_sub15_T_datain = ( (|r_sys_processing_methodID) ? r_sub15_T_datain : 32'h0 ) ;
	assign w_sub15_T_r_w = ( (|r_sys_processing_methodID) ? r_sub15_T_r_w : 1'h0 ) ;
	assign w_sub15_V_addr = ( (|r_sys_processing_methodID) ? r_sub15_V_addr : 10'sh0 ) ;
	assign w_sub15_V_datain = ( (|r_sys_processing_methodID) ? r_sub15_V_datain : 32'h0 ) ;
	assign w_sub15_V_r_w = ( (|r_sys_processing_methodID) ? r_sub15_V_r_w : 1'h0 ) ;
	assign w_sub15_U_addr = ( (|r_sys_processing_methodID) ? r_sub15_U_addr : 10'sh0 ) ;
	assign w_sub15_U_datain = ( (|r_sys_processing_methodID) ? r_sub15_U_datain : 32'h0 ) ;
	assign w_sub15_U_r_w = ( (|r_sys_processing_methodID) ? r_sub15_U_r_w : 1'h0 ) ;
	assign w_sub15_result_addr = ( (|r_sys_processing_methodID) ? r_sub15_result_addr : 10'sh0 ) ;
	assign w_sub15_result_datain = ( (|r_sys_processing_methodID) ? r_sub15_result_datain : 32'h0 ) ;
	assign w_sub15_result_r_w = ( (|r_sys_processing_methodID) ? r_sub15_result_r_w : 1'h0 ) ;
	assign w_sub05_T_addr = ( (|r_sys_processing_methodID) ? r_sub05_T_addr : 10'sh0 ) ;
	assign w_sub05_T_datain = ( (|r_sys_processing_methodID) ? r_sub05_T_datain : 32'h0 ) ;
	assign w_sub05_T_r_w = ( (|r_sys_processing_methodID) ? r_sub05_T_r_w : 1'h0 ) ;
	assign w_sub05_V_addr = ( (|r_sys_processing_methodID) ? r_sub05_V_addr : 10'sh0 ) ;
	assign w_sub05_V_datain = ( (|r_sys_processing_methodID) ? r_sub05_V_datain : 32'h0 ) ;
	assign w_sub05_V_r_w = ( (|r_sys_processing_methodID) ? r_sub05_V_r_w : 1'h0 ) ;
	assign w_sub05_U_addr = ( (|r_sys_processing_methodID) ? r_sub05_U_addr : 10'sh0 ) ;
	assign w_sub05_U_datain = ( (|r_sys_processing_methodID) ? r_sub05_U_datain : 32'h0 ) ;
	assign w_sub05_U_r_w = ( (|r_sys_processing_methodID) ? r_sub05_U_r_w : 1'h0 ) ;
	assign w_sub05_result_addr = ( (|r_sys_processing_methodID) ? r_sub05_result_addr : 10'sh0 ) ;
	assign w_sub05_result_datain = ( (|r_sys_processing_methodID) ? r_sub05_result_datain : 32'h0 ) ;
	assign w_sub05_result_r_w = ( (|r_sys_processing_methodID) ? r_sub05_result_r_w : 1'h0 ) ;
	assign w_sub18_T_addr = ( (|r_sys_processing_methodID) ? r_sub18_T_addr : 10'sh0 ) ;
	assign w_sub18_T_datain = ( (|r_sys_processing_methodID) ? r_sub18_T_datain : 32'h0 ) ;
	assign w_sub18_T_r_w = ( (|r_sys_processing_methodID) ? r_sub18_T_r_w : 1'h0 ) ;
	assign w_sub18_V_addr = ( (|r_sys_processing_methodID) ? r_sub18_V_addr : 10'sh0 ) ;
	assign w_sub18_V_datain = ( (|r_sys_processing_methodID) ? r_sub18_V_datain : 32'h0 ) ;
	assign w_sub18_V_r_w = ( (|r_sys_processing_methodID) ? r_sub18_V_r_w : 1'h0 ) ;
	assign w_sub18_U_addr = ( (|r_sys_processing_methodID) ? r_sub18_U_addr : 10'sh0 ) ;
	assign w_sub18_U_datain = ( (|r_sys_processing_methodID) ? r_sub18_U_datain : 32'h0 ) ;
	assign w_sub18_U_r_w = ( (|r_sys_processing_methodID) ? r_sub18_U_r_w : 1'h0 ) ;
	assign w_sub18_result_addr = ( (|r_sys_processing_methodID) ? r_sub18_result_addr : 10'sh0 ) ;
	assign w_sub18_result_datain = ( (|r_sys_processing_methodID) ? r_sub18_result_datain : 32'h0 ) ;
	assign w_sub18_result_r_w = ( (|r_sys_processing_methodID) ? r_sub18_result_r_w : 1'h0 ) ;
	assign w_sub04_T_addr = ( (|r_sys_processing_methodID) ? r_sub04_T_addr : 10'sh0 ) ;
	assign w_sub04_T_datain = ( (|r_sys_processing_methodID) ? r_sub04_T_datain : 32'h0 ) ;
	assign w_sub04_T_r_w = ( (|r_sys_processing_methodID) ? r_sub04_T_r_w : 1'h0 ) ;
	assign w_sub04_V_addr = ( (|r_sys_processing_methodID) ? r_sub04_V_addr : 10'sh0 ) ;
	assign w_sub04_V_datain = ( (|r_sys_processing_methodID) ? r_sub04_V_datain : 32'h0 ) ;
	assign w_sub04_V_r_w = ( (|r_sys_processing_methodID) ? r_sub04_V_r_w : 1'h0 ) ;
	assign w_sub04_U_addr = ( (|r_sys_processing_methodID) ? r_sub04_U_addr : 10'sh0 ) ;
	assign w_sub04_U_datain = ( (|r_sys_processing_methodID) ? r_sub04_U_datain : 32'h0 ) ;
	assign w_sub04_U_r_w = ( (|r_sys_processing_methodID) ? r_sub04_U_r_w : 1'h0 ) ;
	assign w_sub04_result_addr = ( (|r_sys_processing_methodID) ? r_sub04_result_addr : 10'sh0 ) ;
	assign w_sub04_result_datain = ( (|r_sys_processing_methodID) ? r_sub04_result_datain : 32'h0 ) ;
	assign w_sub04_result_r_w = ( (|r_sys_processing_methodID) ? r_sub04_result_r_w : 1'h0 ) ;
	assign w_sub17_T_addr = ( (|r_sys_processing_methodID) ? r_sub17_T_addr : 10'sh0 ) ;
	assign w_sub17_T_datain = ( (|r_sys_processing_methodID) ? r_sub17_T_datain : 32'h0 ) ;
	assign w_sub17_T_r_w = ( (|r_sys_processing_methodID) ? r_sub17_T_r_w : 1'h0 ) ;
	assign w_sub17_V_addr = ( (|r_sys_processing_methodID) ? r_sub17_V_addr : 10'sh0 ) ;
	assign w_sub17_V_datain = ( (|r_sys_processing_methodID) ? r_sub17_V_datain : 32'h0 ) ;
	assign w_sub17_V_r_w = ( (|r_sys_processing_methodID) ? r_sub17_V_r_w : 1'h0 ) ;
	assign w_sub17_U_addr = ( (|r_sys_processing_methodID) ? r_sub17_U_addr : 10'sh0 ) ;
	assign w_sub17_U_datain = ( (|r_sys_processing_methodID) ? r_sub17_U_datain : 32'h0 ) ;
	assign w_sub17_U_r_w = ( (|r_sys_processing_methodID) ? r_sub17_U_r_w : 1'h0 ) ;
	assign w_sub17_result_addr = ( (|r_sys_processing_methodID) ? r_sub17_result_addr : 10'sh0 ) ;
	assign w_sub17_result_datain = ( (|r_sys_processing_methodID) ? r_sub17_result_datain : 32'h0 ) ;
	assign w_sub17_result_r_w = ( (|r_sys_processing_methodID) ? r_sub17_result_r_w : 1'h0 ) ;
	assign w_sub10_T_addr = ( (|r_sys_processing_methodID) ? r_sub10_T_addr : 10'sh0 ) ;
	assign w_sub10_T_datain = ( (|r_sys_processing_methodID) ? r_sub10_T_datain : 32'h0 ) ;
	assign w_sub10_T_r_w = ( (|r_sys_processing_methodID) ? r_sub10_T_r_w : 1'h0 ) ;
	assign w_sub10_V_addr = ( (|r_sys_processing_methodID) ? r_sub10_V_addr : 10'sh0 ) ;
	assign w_sub10_V_datain = ( (|r_sys_processing_methodID) ? r_sub10_V_datain : 32'h0 ) ;
	assign w_sub10_V_r_w = ( (|r_sys_processing_methodID) ? r_sub10_V_r_w : 1'h0 ) ;
	assign w_sub10_U_addr = ( (|r_sys_processing_methodID) ? r_sub10_U_addr : 10'sh0 ) ;
	assign w_sub10_U_datain = ( (|r_sys_processing_methodID) ? r_sub10_U_datain : 32'h0 ) ;
	assign w_sub10_U_r_w = ( (|r_sys_processing_methodID) ? r_sub10_U_r_w : 1'h0 ) ;
	assign w_sub10_result_addr = ( (|r_sys_processing_methodID) ? r_sub10_result_addr : 10'sh0 ) ;
	assign w_sub10_result_datain = ( (|r_sys_processing_methodID) ? r_sub10_result_datain : 32'h0 ) ;
	assign w_sub10_result_r_w = ( (|r_sys_processing_methodID) ? r_sub10_result_r_w : 1'h0 ) ;
	assign w_sub20_T_addr = ( (|r_sys_processing_methodID) ? r_sub20_T_addr : 10'sh0 ) ;
	assign w_sub20_T_datain = ( (|r_sys_processing_methodID) ? r_sub20_T_datain : 32'h0 ) ;
	assign w_sub20_T_r_w = ( (|r_sys_processing_methodID) ? r_sub20_T_r_w : 1'h0 ) ;
	assign w_sub20_V_addr = ( (|r_sys_processing_methodID) ? r_sub20_V_addr : 10'sh0 ) ;
	assign w_sub20_V_datain = ( (|r_sys_processing_methodID) ? r_sub20_V_datain : 32'h0 ) ;
	assign w_sub20_V_r_w = ( (|r_sys_processing_methodID) ? r_sub20_V_r_w : 1'h0 ) ;
	assign w_sub20_U_addr = ( (|r_sys_processing_methodID) ? r_sub20_U_addr : 10'sh0 ) ;
	assign w_sub20_U_datain = ( (|r_sys_processing_methodID) ? r_sub20_U_datain : 32'h0 ) ;
	assign w_sub20_U_r_w = ( (|r_sys_processing_methodID) ? r_sub20_U_r_w : 1'h0 ) ;
	assign w_sub20_result_addr = ( (|r_sys_processing_methodID) ? r_sub20_result_addr : 10'sh0 ) ;
	assign w_sub20_result_datain = ( (|r_sys_processing_methodID) ? r_sub20_result_datain : 32'h0 ) ;
	assign w_sub20_result_r_w = ( (|r_sys_processing_methodID) ? r_sub20_result_r_w : 1'h0 ) ;
	assign w_sub21_T_addr = ( (|r_sys_processing_methodID) ? r_sub21_T_addr : 10'sh0 ) ;
	assign w_sub21_T_datain = ( (|r_sys_processing_methodID) ? r_sub21_T_datain : 32'h0 ) ;
	assign w_sub21_T_r_w = ( (|r_sys_processing_methodID) ? r_sub21_T_r_w : 1'h0 ) ;
	assign w_sub21_V_addr = ( (|r_sys_processing_methodID) ? r_sub21_V_addr : 10'sh0 ) ;
	assign w_sub21_V_datain = ( (|r_sys_processing_methodID) ? r_sub21_V_datain : 32'h0 ) ;
	assign w_sub21_V_r_w = ( (|r_sys_processing_methodID) ? r_sub21_V_r_w : 1'h0 ) ;
	assign w_sub21_U_addr = ( (|r_sys_processing_methodID) ? r_sub21_U_addr : 10'sh0 ) ;
	assign w_sub21_U_datain = ( (|r_sys_processing_methodID) ? r_sub21_U_datain : 32'h0 ) ;
	assign w_sub21_U_r_w = ( (|r_sys_processing_methodID) ? r_sub21_U_r_w : 1'h0 ) ;
	assign w_sub21_result_addr = ( (|r_sys_processing_methodID) ? r_sub21_result_addr : 10'sh0 ) ;
	assign w_sub21_result_datain = ( (|r_sys_processing_methodID) ? r_sub21_result_datain : 32'h0 ) ;
	assign w_sub21_result_r_w = ( (|r_sys_processing_methodID) ? r_sub21_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh0000001e;
	assign w_sys_tmp3 = 32'sh0000001f;
	assign w_sys_tmp5 = 32'h3a03126f;
	assign w_sys_tmp6 = 32'sh00000002;
	assign w_sys_tmp7 = 32'h3e088889;
	assign w_sys_tmp8 = 32'h3d088889;
	assign w_sys_tmp9 = 32'h3af5c28f;
	assign w_sys_tmp10 = 32'h3bf5c28f;
	assign w_sys_tmp11 = 32'h3ce66665;
	assign w_sys_tmp12 = 32'h3ee66665;
	assign w_sys_tmp13 = ( !w_sys_tmp14 );
	assign w_sys_tmp14 = (r_run_my_33 < r_run_k_29);
	assign w_sys_tmp15 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp16 = ( !w_sys_tmp17 );
	assign w_sys_tmp17 = (r_run_mx_32 < r_run_j_30);
	assign w_sys_tmp19 = w_ip_MultFloat_product_0;
	assign w_sys_tmp20 = w_ip_FixedToFloat_floating_0;
	assign w_sys_tmp21 = (r_run_k_29 - w_sys_intOne);
	assign w_sys_tmp23 = (w_sys_tmp24 + r_run_k_29);
	assign w_sys_tmp24 = (r_run_j_30 * w_sys_tmp25);
	assign w_sys_tmp25 = 32'sh0000001f;
	assign w_sys_tmp26 = 32'h0;
	assign w_sys_tmp28 = (w_sys_tmp29 + r_run_k_29);
	assign w_sys_tmp29 = (r_run_copy2_j_47 * w_sys_tmp25);
	assign w_sys_tmp33 = (w_sys_tmp34 + r_run_k_29);
	assign w_sys_tmp34 = (r_run_copy1_j_46 * w_sys_tmp25);
	assign w_sys_tmp37 = 32'h42200000;
	assign w_sys_tmp38 = w_sys_tmp19;
	assign w_sys_tmp39 = 32'h3f800000;
	assign w_sys_tmp42 = (w_sys_tmp43 + r_run_k_29);
	assign w_sys_tmp43 = (r_run_copy0_j_45 * w_sys_tmp25);
	assign w_sys_tmp46 = (r_run_copy0_j_45 + w_sys_intOne);
	assign w_sys_tmp47 = (r_run_copy1_j_46 + w_sys_intOne);
	assign w_sys_tmp48 = (r_run_copy2_j_47 + w_sys_intOne);
	assign w_sys_tmp49 = (r_run_j_30 + w_sys_intOne);
	assign w_sys_tmp129 = r_sys_tmp4_float;
	assign w_sys_tmp227 = ( !w_sys_tmp228 );
	assign w_sys_tmp228 = (w_sys_tmp229 < r_run_k_29);
	assign w_sys_tmp229 = 32'sh00000008;
	assign w_sys_tmp232 = (w_sys_tmp233 + r_run_k_29);
	assign w_sys_tmp233 = 32'sh0000001f;
	assign w_sys_tmp234 = w_fld_U_2_dataout_1;
	assign w_sys_tmp240 = w_fld_V_3_dataout_1;
	assign w_sys_tmp244 = (w_sys_tmp245 + r_run_k_29);
	assign w_sys_tmp245 = 32'sh0000003e;
	assign w_sys_tmp256 = (w_sys_tmp257 + r_run_k_29);
	assign w_sys_tmp257 = 32'sh0000005d;
	assign w_sys_tmp268 = (w_sys_tmp269 + r_run_k_29);
	assign w_sys_tmp269 = 32'sh0000007c;
	assign w_sys_tmp280 = (w_sys_tmp281 + r_run_k_29);
	assign w_sys_tmp281 = 32'sh0000009b;
	assign w_sys_tmp292 = (w_sys_tmp293 + r_run_k_29);
	assign w_sys_tmp293 = 32'sh000000ba;
	assign w_sys_tmp304 = (w_sys_tmp305 + r_run_k_29);
	assign w_sys_tmp305 = 32'sh000000d9;
	assign w_sys_tmp316 = (w_sys_tmp317 + r_run_k_29);
	assign w_sys_tmp317 = 32'sh000000f8;
	assign w_sys_tmp352 = (w_sys_tmp353 + r_run_k_29);
	assign w_sys_tmp353 = 32'sh00000117;
	assign w_sys_tmp364 = (w_sys_tmp365 + r_run_k_29);
	assign w_sys_tmp365 = 32'sh00000136;
	assign w_sys_tmp376 = (w_sys_tmp377 + r_run_k_29);
	assign w_sys_tmp377 = 32'sh00000155;
	assign w_sys_tmp388 = (w_sys_tmp389 + r_run_k_29);
	assign w_sys_tmp389 = 32'sh00000174;
	assign w_sys_tmp400 = (w_sys_tmp401 + r_run_k_29);
	assign w_sys_tmp401 = 32'sh00000193;
	assign w_sys_tmp412 = (w_sys_tmp413 + r_run_k_29);
	assign w_sys_tmp413 = 32'sh000001b2;
	assign w_sys_tmp448 = (w_sys_tmp449 + r_run_k_29);
	assign w_sys_tmp449 = 32'sh000001d1;
	assign w_sys_tmp460 = (w_sys_tmp461 + r_run_k_29);
	assign w_sys_tmp461 = 32'sh000001f0;
	assign w_sys_tmp472 = (w_sys_tmp473 + r_run_k_29);
	assign w_sys_tmp473 = 32'sh0000020f;
	assign w_sys_tmp484 = (w_sys_tmp485 + r_run_k_29);
	assign w_sys_tmp485 = 32'sh0000022e;
	assign w_sys_tmp496 = (w_sys_tmp497 + r_run_k_29);
	assign w_sys_tmp497 = 32'sh0000024d;
	assign w_sys_tmp508 = (w_sys_tmp509 + r_run_k_29);
	assign w_sys_tmp509 = 32'sh0000026c;
	assign w_sys_tmp544 = (w_sys_tmp545 + r_run_k_29);
	assign w_sys_tmp545 = 32'sh0000028b;
	assign w_sys_tmp556 = (w_sys_tmp557 + r_run_k_29);
	assign w_sys_tmp557 = 32'sh000002aa;
	assign w_sys_tmp568 = (w_sys_tmp569 + r_run_k_29);
	assign w_sys_tmp569 = 32'sh000002c9;
	assign w_sys_tmp580 = (w_sys_tmp581 + r_run_k_29);
	assign w_sys_tmp581 = 32'sh000002e8;
	assign w_sys_tmp592 = (w_sys_tmp593 + r_run_k_29);
	assign w_sys_tmp593 = 32'sh00000307;
	assign w_sys_tmp604 = (w_sys_tmp605 + r_run_k_29);
	assign w_sys_tmp605 = 32'sh00000326;
	assign w_sys_tmp640 = (w_sys_tmp641 + r_run_k_29);
	assign w_sys_tmp641 = 32'sh00000345;
	assign w_sys_tmp652 = (w_sys_tmp653 + r_run_k_29);
	assign w_sys_tmp653 = 32'sh00000364;
	assign w_sys_tmp664 = (w_sys_tmp665 + r_run_k_29);
	assign w_sys_tmp665 = 32'sh00000383;
	assign w_sys_tmp676 = (w_sys_tmp677 + r_run_k_29);
	assign w_sys_tmp677 = 32'sh000003a2;
	assign w_sys_tmp688 = (w_sys_tmp689 + r_run_k_29);
	assign w_sys_tmp689 = 32'sh000003c1;
	assign w_sys_tmp700 = (w_sys_tmp701 + r_run_k_29);
	assign w_sys_tmp701 = 32'sh00000025;
	assign w_sys_tmp712 = (w_sys_tmp713 + r_run_k_29);
	assign w_sys_tmp713 = 32'sh00000044;
	assign w_sys_tmp724 = (w_sys_tmp725 + r_run_k_29);
	assign w_sys_tmp725 = 32'sh00000063;
	assign w_sys_tmp736 = (w_sys_tmp737 + r_run_k_29);
	assign w_sys_tmp737 = 32'sh00000082;
	assign w_sys_tmp748 = (w_sys_tmp749 + r_run_k_29);
	assign w_sys_tmp749 = 32'sh000000a1;
	assign w_sys_tmp760 = (w_sys_tmp761 + r_run_k_29);
	assign w_sys_tmp761 = 32'sh000000c0;
	assign w_sys_tmp772 = (w_sys_tmp773 + r_run_k_29);
	assign w_sys_tmp773 = 32'sh000000df;
	assign w_sys_tmp784 = (w_sys_tmp785 + r_run_k_29);
	assign w_sys_tmp785 = 32'sh000000fe;
	assign w_sys_tmp820 = (w_sys_tmp821 + r_run_k_29);
	assign w_sys_tmp821 = 32'sh0000011d;
	assign w_sys_tmp832 = (w_sys_tmp833 + r_run_k_29);
	assign w_sys_tmp833 = 32'sh0000013c;
	assign w_sys_tmp844 = (w_sys_tmp845 + r_run_k_29);
	assign w_sys_tmp845 = 32'sh0000015b;
	assign w_sys_tmp856 = (w_sys_tmp857 + r_run_k_29);
	assign w_sys_tmp857 = 32'sh0000017a;
	assign w_sys_tmp868 = (w_sys_tmp869 + r_run_k_29);
	assign w_sys_tmp869 = 32'sh00000199;
	assign w_sys_tmp880 = (w_sys_tmp881 + r_run_k_29);
	assign w_sys_tmp881 = 32'sh000001b8;
	assign w_sys_tmp916 = (w_sys_tmp917 + r_run_k_29);
	assign w_sys_tmp917 = 32'sh000001d7;
	assign w_sys_tmp928 = (w_sys_tmp929 + r_run_k_29);
	assign w_sys_tmp929 = 32'sh000001f6;
	assign w_sys_tmp940 = (w_sys_tmp941 + r_run_k_29);
	assign w_sys_tmp941 = 32'sh00000215;
	assign w_sys_tmp952 = (w_sys_tmp953 + r_run_k_29);
	assign w_sys_tmp953 = 32'sh00000234;
	assign w_sys_tmp964 = (w_sys_tmp965 + r_run_k_29);
	assign w_sys_tmp965 = 32'sh00000253;
	assign w_sys_tmp976 = (w_sys_tmp977 + r_run_k_29);
	assign w_sys_tmp977 = 32'sh00000272;
	assign w_sys_tmp1012 = (w_sys_tmp1013 + r_run_k_29);
	assign w_sys_tmp1013 = 32'sh00000291;
	assign w_sys_tmp1024 = (w_sys_tmp1025 + r_run_k_29);
	assign w_sys_tmp1025 = 32'sh000002b0;
	assign w_sys_tmp1036 = (w_sys_tmp1037 + r_run_k_29);
	assign w_sys_tmp1037 = 32'sh000002cf;
	assign w_sys_tmp1048 = (w_sys_tmp1049 + r_run_k_29);
	assign w_sys_tmp1049 = 32'sh000002ee;
	assign w_sys_tmp1060 = (w_sys_tmp1061 + r_run_k_29);
	assign w_sys_tmp1061 = 32'sh0000030d;
	assign w_sys_tmp1072 = (w_sys_tmp1073 + r_run_k_29);
	assign w_sys_tmp1073 = 32'sh0000032c;
	assign w_sys_tmp1108 = (w_sys_tmp1109 + r_run_k_29);
	assign w_sys_tmp1109 = 32'sh0000034b;
	assign w_sys_tmp1120 = (w_sys_tmp1121 + r_run_k_29);
	assign w_sys_tmp1121 = 32'sh0000036a;
	assign w_sys_tmp1132 = (w_sys_tmp1133 + r_run_k_29);
	assign w_sys_tmp1133 = 32'sh00000389;
	assign w_sys_tmp1144 = (w_sys_tmp1145 + r_run_k_29);
	assign w_sys_tmp1145 = 32'sh000003a8;
	assign w_sys_tmp1156 = (w_sys_tmp1157 + r_run_k_29);
	assign w_sys_tmp1157 = 32'sh000003c7;
	assign w_sys_tmp1168 = (w_sys_tmp1169 + r_run_k_29);
	assign w_sys_tmp1169 = 32'sh0000002b;
	assign w_sys_tmp1180 = (w_sys_tmp1181 + r_run_k_29);
	assign w_sys_tmp1181 = 32'sh0000004a;
	assign w_sys_tmp1192 = (w_sys_tmp1193 + r_run_k_29);
	assign w_sys_tmp1193 = 32'sh00000069;
	assign w_sys_tmp1204 = (w_sys_tmp1205 + r_run_k_29);
	assign w_sys_tmp1205 = 32'sh00000088;
	assign w_sys_tmp1216 = (w_sys_tmp1217 + r_run_k_29);
	assign w_sys_tmp1217 = 32'sh000000a7;
	assign w_sys_tmp1228 = (w_sys_tmp1229 + r_run_k_29);
	assign w_sys_tmp1229 = 32'sh000000c6;
	assign w_sys_tmp1240 = (w_sys_tmp1241 + r_run_k_29);
	assign w_sys_tmp1241 = 32'sh000000e5;
	assign w_sys_tmp1252 = (w_sys_tmp1253 + r_run_k_29);
	assign w_sys_tmp1253 = 32'sh00000104;
	assign w_sys_tmp1288 = (w_sys_tmp1289 + r_run_k_29);
	assign w_sys_tmp1289 = 32'sh00000123;
	assign w_sys_tmp1300 = (w_sys_tmp1301 + r_run_k_29);
	assign w_sys_tmp1301 = 32'sh00000142;
	assign w_sys_tmp1312 = (w_sys_tmp1313 + r_run_k_29);
	assign w_sys_tmp1313 = 32'sh00000161;
	assign w_sys_tmp1324 = (w_sys_tmp1325 + r_run_k_29);
	assign w_sys_tmp1325 = 32'sh00000180;
	assign w_sys_tmp1336 = (w_sys_tmp1337 + r_run_k_29);
	assign w_sys_tmp1337 = 32'sh0000019f;
	assign w_sys_tmp1348 = (w_sys_tmp1349 + r_run_k_29);
	assign w_sys_tmp1349 = 32'sh000001be;
	assign w_sys_tmp1384 = (w_sys_tmp1385 + r_run_k_29);
	assign w_sys_tmp1385 = 32'sh000001dd;
	assign w_sys_tmp1396 = (w_sys_tmp1397 + r_run_k_29);
	assign w_sys_tmp1397 = 32'sh000001fc;
	assign w_sys_tmp1408 = (w_sys_tmp1409 + r_run_k_29);
	assign w_sys_tmp1409 = 32'sh0000021b;
	assign w_sys_tmp1420 = (w_sys_tmp1421 + r_run_k_29);
	assign w_sys_tmp1421 = 32'sh0000023a;
	assign w_sys_tmp1432 = (w_sys_tmp1433 + r_run_k_29);
	assign w_sys_tmp1433 = 32'sh00000259;
	assign w_sys_tmp1444 = (w_sys_tmp1445 + r_run_k_29);
	assign w_sys_tmp1445 = 32'sh00000278;
	assign w_sys_tmp1480 = (w_sys_tmp1481 + r_run_k_29);
	assign w_sys_tmp1481 = 32'sh00000297;
	assign w_sys_tmp1492 = (w_sys_tmp1493 + r_run_k_29);
	assign w_sys_tmp1493 = 32'sh000002b6;
	assign w_sys_tmp1504 = (w_sys_tmp1505 + r_run_k_29);
	assign w_sys_tmp1505 = 32'sh000002d5;
	assign w_sys_tmp1516 = (w_sys_tmp1517 + r_run_k_29);
	assign w_sys_tmp1517 = 32'sh000002f4;
	assign w_sys_tmp1528 = (w_sys_tmp1529 + r_run_k_29);
	assign w_sys_tmp1529 = 32'sh00000313;
	assign w_sys_tmp1540 = (w_sys_tmp1541 + r_run_k_29);
	assign w_sys_tmp1541 = 32'sh00000332;
	assign w_sys_tmp1576 = (w_sys_tmp1577 + r_run_k_29);
	assign w_sys_tmp1577 = 32'sh00000351;
	assign w_sys_tmp1588 = (w_sys_tmp1589 + r_run_k_29);
	assign w_sys_tmp1589 = 32'sh00000370;
	assign w_sys_tmp1600 = (w_sys_tmp1601 + r_run_k_29);
	assign w_sys_tmp1601 = 32'sh0000038f;
	assign w_sys_tmp1612 = (w_sys_tmp1613 + r_run_k_29);
	assign w_sys_tmp1613 = 32'sh000003ae;
	assign w_sys_tmp1624 = (w_sys_tmp1625 + r_run_k_29);
	assign w_sys_tmp1625 = 32'sh000003cd;
	assign w_sys_tmp1636 = (w_sys_tmp1637 + r_run_k_29);
	assign w_sys_tmp1637 = 32'sh00000031;
	assign w_sys_tmp1648 = (w_sys_tmp1649 + r_run_k_29);
	assign w_sys_tmp1649 = 32'sh00000050;
	assign w_sys_tmp1660 = (w_sys_tmp1661 + r_run_k_29);
	assign w_sys_tmp1661 = 32'sh0000006f;
	assign w_sys_tmp1672 = (w_sys_tmp1673 + r_run_k_29);
	assign w_sys_tmp1673 = 32'sh0000008e;
	assign w_sys_tmp1684 = (w_sys_tmp1685 + r_run_k_29);
	assign w_sys_tmp1685 = 32'sh000000ad;
	assign w_sys_tmp1696 = (w_sys_tmp1697 + r_run_k_29);
	assign w_sys_tmp1697 = 32'sh000000cc;
	assign w_sys_tmp1708 = (w_sys_tmp1709 + r_run_k_29);
	assign w_sys_tmp1709 = 32'sh000000eb;
	assign w_sys_tmp1720 = (w_sys_tmp1721 + r_run_k_29);
	assign w_sys_tmp1721 = 32'sh0000010a;
	assign w_sys_tmp1756 = (w_sys_tmp1757 + r_run_k_29);
	assign w_sys_tmp1757 = 32'sh00000129;
	assign w_sys_tmp1768 = (w_sys_tmp1769 + r_run_k_29);
	assign w_sys_tmp1769 = 32'sh00000148;
	assign w_sys_tmp1780 = (w_sys_tmp1781 + r_run_k_29);
	assign w_sys_tmp1781 = 32'sh00000167;
	assign w_sys_tmp1792 = (w_sys_tmp1793 + r_run_k_29);
	assign w_sys_tmp1793 = 32'sh00000186;
	assign w_sys_tmp1804 = (w_sys_tmp1805 + r_run_k_29);
	assign w_sys_tmp1805 = 32'sh000001a5;
	assign w_sys_tmp1816 = (w_sys_tmp1817 + r_run_k_29);
	assign w_sys_tmp1817 = 32'sh000001c4;
	assign w_sys_tmp1852 = (w_sys_tmp1853 + r_run_k_29);
	assign w_sys_tmp1853 = 32'sh000001e3;
	assign w_sys_tmp1864 = (w_sys_tmp1865 + r_run_k_29);
	assign w_sys_tmp1865 = 32'sh00000202;
	assign w_sys_tmp1876 = (w_sys_tmp1877 + r_run_k_29);
	assign w_sys_tmp1877 = 32'sh00000221;
	assign w_sys_tmp1888 = (w_sys_tmp1889 + r_run_k_29);
	assign w_sys_tmp1889 = 32'sh00000240;
	assign w_sys_tmp1900 = (w_sys_tmp1901 + r_run_k_29);
	assign w_sys_tmp1901 = 32'sh0000025f;
	assign w_sys_tmp1912 = (w_sys_tmp1913 + r_run_k_29);
	assign w_sys_tmp1913 = 32'sh0000027e;
	assign w_sys_tmp1948 = (w_sys_tmp1949 + r_run_k_29);
	assign w_sys_tmp1949 = 32'sh0000029d;
	assign w_sys_tmp1960 = (w_sys_tmp1961 + r_run_k_29);
	assign w_sys_tmp1961 = 32'sh000002bc;
	assign w_sys_tmp1972 = (w_sys_tmp1973 + r_run_k_29);
	assign w_sys_tmp1973 = 32'sh000002db;
	assign w_sys_tmp1984 = (w_sys_tmp1985 + r_run_k_29);
	assign w_sys_tmp1985 = 32'sh000002fa;
	assign w_sys_tmp1996 = (w_sys_tmp1997 + r_run_k_29);
	assign w_sys_tmp1997 = 32'sh00000319;
	assign w_sys_tmp2008 = (w_sys_tmp2009 + r_run_k_29);
	assign w_sys_tmp2009 = 32'sh00000338;
	assign w_sys_tmp2044 = (w_sys_tmp2045 + r_run_k_29);
	assign w_sys_tmp2045 = 32'sh00000357;
	assign w_sys_tmp2056 = (w_sys_tmp2057 + r_run_k_29);
	assign w_sys_tmp2057 = 32'sh00000376;
	assign w_sys_tmp2068 = (w_sys_tmp2069 + r_run_k_29);
	assign w_sys_tmp2069 = 32'sh00000395;
	assign w_sys_tmp2080 = (w_sys_tmp2081 + r_run_k_29);
	assign w_sys_tmp2081 = 32'sh000003b4;
	assign w_sys_tmp2092 = (w_sys_tmp2093 + r_run_k_29);
	assign w_sys_tmp2093 = 32'sh000003d3;
	assign w_sys_tmp2103 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp2104 = 32'sh00000019;
	assign w_sys_tmp2105 = ( !w_sys_tmp2106 );
	assign w_sys_tmp2106 = (w_sys_tmp2107 < r_run_k_29);
	assign w_sys_tmp2107 = 32'sh0000001f;
	assign w_sys_tmp2110 = (w_sys_tmp2111 + r_run_k_29);
	assign w_sys_tmp2111 = 32'sh0000001f;
	assign w_sys_tmp2112 = w_fld_U_2_dataout_1;
	assign w_sys_tmp2118 = w_fld_V_3_dataout_1;
	assign w_sys_tmp2122 = (w_sys_tmp2123 + r_run_k_29);
	assign w_sys_tmp2123 = 32'sh0000003e;
	assign w_sys_tmp2134 = (w_sys_tmp2135 + r_run_k_29);
	assign w_sys_tmp2135 = 32'sh0000005d;
	assign w_sys_tmp2146 = (w_sys_tmp2147 + r_run_k_29);
	assign w_sys_tmp2147 = 32'sh0000007c;
	assign w_sys_tmp2158 = (w_sys_tmp2159 + r_run_k_29);
	assign w_sys_tmp2159 = 32'sh0000009b;
	assign w_sys_tmp2170 = (w_sys_tmp2171 + r_run_k_29);
	assign w_sys_tmp2171 = 32'sh000000ba;
	assign w_sys_tmp2182 = (w_sys_tmp2183 + r_run_k_29);
	assign w_sys_tmp2183 = 32'sh000000d9;
	assign w_sys_tmp2194 = (w_sys_tmp2195 + r_run_k_29);
	assign w_sys_tmp2195 = 32'sh000000f8;
	assign w_sys_tmp2230 = (w_sys_tmp2231 + r_run_k_29);
	assign w_sys_tmp2231 = 32'sh00000117;
	assign w_sys_tmp2242 = (w_sys_tmp2243 + r_run_k_29);
	assign w_sys_tmp2243 = 32'sh00000136;
	assign w_sys_tmp2254 = (w_sys_tmp2255 + r_run_k_29);
	assign w_sys_tmp2255 = 32'sh00000155;
	assign w_sys_tmp2266 = (w_sys_tmp2267 + r_run_k_29);
	assign w_sys_tmp2267 = 32'sh00000174;
	assign w_sys_tmp2278 = (w_sys_tmp2279 + r_run_k_29);
	assign w_sys_tmp2279 = 32'sh00000193;
	assign w_sys_tmp2290 = (w_sys_tmp2291 + r_run_k_29);
	assign w_sys_tmp2291 = 32'sh000001b2;
	assign w_sys_tmp2326 = (w_sys_tmp2327 + r_run_k_29);
	assign w_sys_tmp2327 = 32'sh000001d1;
	assign w_sys_tmp2338 = (w_sys_tmp2339 + r_run_k_29);
	assign w_sys_tmp2339 = 32'sh000001f0;
	assign w_sys_tmp2350 = (w_sys_tmp2351 + r_run_k_29);
	assign w_sys_tmp2351 = 32'sh0000020f;
	assign w_sys_tmp2362 = (w_sys_tmp2363 + r_run_k_29);
	assign w_sys_tmp2363 = 32'sh0000022e;
	assign w_sys_tmp2374 = (w_sys_tmp2375 + r_run_k_29);
	assign w_sys_tmp2375 = 32'sh0000024d;
	assign w_sys_tmp2386 = (w_sys_tmp2387 + r_run_k_29);
	assign w_sys_tmp2387 = 32'sh0000026c;
	assign w_sys_tmp2422 = (w_sys_tmp2423 + r_run_k_29);
	assign w_sys_tmp2423 = 32'sh0000028b;
	assign w_sys_tmp2434 = (w_sys_tmp2435 + r_run_k_29);
	assign w_sys_tmp2435 = 32'sh000002aa;
	assign w_sys_tmp2446 = (w_sys_tmp2447 + r_run_k_29);
	assign w_sys_tmp2447 = 32'sh000002c9;
	assign w_sys_tmp2458 = (w_sys_tmp2459 + r_run_k_29);
	assign w_sys_tmp2459 = 32'sh000002e8;
	assign w_sys_tmp2470 = (w_sys_tmp2471 + r_run_k_29);
	assign w_sys_tmp2471 = 32'sh00000307;
	assign w_sys_tmp2482 = (w_sys_tmp2483 + r_run_k_29);
	assign w_sys_tmp2483 = 32'sh00000326;
	assign w_sys_tmp2518 = (w_sys_tmp2519 + r_run_k_29);
	assign w_sys_tmp2519 = 32'sh00000345;
	assign w_sys_tmp2530 = (w_sys_tmp2531 + r_run_k_29);
	assign w_sys_tmp2531 = 32'sh00000364;
	assign w_sys_tmp2542 = (w_sys_tmp2543 + r_run_k_29);
	assign w_sys_tmp2543 = 32'sh00000383;
	assign w_sys_tmp2554 = (w_sys_tmp2555 + r_run_k_29);
	assign w_sys_tmp2555 = 32'sh000003a2;
	assign w_sys_tmp2566 = (w_sys_tmp2567 + r_run_k_29);
	assign w_sys_tmp2567 = 32'sh000003c1;
	assign w_sys_tmp2577 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp2578 = ( !w_sys_tmp2579 );
	assign w_sys_tmp2579 = (r_run_nlast_44 < r_run_n_31);
	assign w_sys_tmp2580 = (r_run_n_31 + w_sys_intOne);
	assign w_sys_tmp2581 = ( !w_sys_tmp2582 );
	assign w_sys_tmp2582 = (r_run_my_33 < r_run_k_29);
	assign w_sys_tmp2585 = (w_sys_tmp2586 + r_run_k_29);
	assign w_sys_tmp2586 = 32'sh0000001f;
	assign w_sys_tmp2587 = 32'h0;
	assign w_sys_tmp2589 = (w_sys_tmp2590 + r_run_k_29);
	assign w_sys_tmp2590 = (r_run_mx_32 * w_sys_tmp2586);
	assign w_sys_tmp2592 = w_fld_T_0_dataout_1;
	assign w_sys_tmp2593 = (w_sys_tmp2594 + r_run_k_29);
	assign w_sys_tmp2594 = (w_sys_tmp2595 * w_sys_tmp2586);
	assign w_sys_tmp2595 = (r_run_mx_32 - w_sys_intOne);
	assign w_sys_tmp2597 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp2598 = ( !w_sys_tmp2599 );
	assign w_sys_tmp2599 = (r_run_mx_32 < r_run_j_30);
	assign w_sys_tmp2602 = (w_sys_tmp2603 + w_sys_intOne);
	assign w_sys_tmp2603 = (r_run_j_30 * w_sys_tmp2604);
	assign w_sys_tmp2604 = 32'sh0000001f;
	assign w_sys_tmp2605 = 32'h0;
	assign w_sys_tmp2607 = (w_sys_tmp2608 + r_run_my_33);
	assign w_sys_tmp2608 = (r_run_copy0_j_48 * w_sys_tmp2604);
	assign w_sys_tmp2611 = (r_run_copy0_j_48 + w_sys_intOne);
	assign w_sys_tmp2612 = (r_run_j_30 + w_sys_intOne);
	assign w_sys_tmp2685 = w_ip_DivInt_quotient_0;
	assign w_sys_tmp2686 = 32'sh00000004;
	assign w_sys_tmp2687 = ( !w_sys_tmp2688 );
	assign w_sys_tmp2688 = (w_sys_tmp2689 < r_run_j_30);
	assign w_sys_tmp2689 = w_ip_DivInt_quotient_1;
	assign w_sys_tmp2690 = 32'sh00000002;
	assign w_sys_tmp2693 = (w_sys_tmp2694 + w_sys_intOne);
	assign w_sys_tmp2694 = (r_run_j_30 * w_sys_tmp2695);
	assign w_sys_tmp2695 = 32'sh0000001f;
	assign w_sys_tmp2696 = 32'h3f800000;
	assign w_sys_tmp2697 = (r_run_j_30 + w_sys_intOne);
	assign w_sys_tmp2734 = ( !w_sys_tmp2735 );
	assign w_sys_tmp2735 = (w_sys_tmp2736 < r_run_k_29);
	assign w_sys_tmp2736 = 32'sh00000008;
	assign w_sys_tmp2739 = (w_sys_tmp2740 + r_run_k_29);
	assign w_sys_tmp2740 = 32'sh0000001f;
	assign w_sys_tmp2741 = w_fld_T_0_dataout_1;
	assign w_sys_tmp2745 = (w_sys_tmp2746 + r_run_k_29);
	assign w_sys_tmp2746 = 32'sh0000003e;
	assign w_sys_tmp2751 = (w_sys_tmp2752 + r_run_k_29);
	assign w_sys_tmp2752 = 32'sh0000005d;
	assign w_sys_tmp2757 = (w_sys_tmp2758 + r_run_k_29);
	assign w_sys_tmp2758 = 32'sh0000007c;
	assign w_sys_tmp2763 = (w_sys_tmp2764 + r_run_k_29);
	assign w_sys_tmp2764 = 32'sh0000009b;
	assign w_sys_tmp2769 = (w_sys_tmp2770 + r_run_k_29);
	assign w_sys_tmp2770 = 32'sh000000ba;
	assign w_sys_tmp2775 = (w_sys_tmp2776 + r_run_k_29);
	assign w_sys_tmp2776 = 32'sh000000d9;
	assign w_sys_tmp2781 = (w_sys_tmp2782 + r_run_k_29);
	assign w_sys_tmp2782 = 32'sh000000f8;
	assign w_sys_tmp2799 = (w_sys_tmp2800 + r_run_k_29);
	assign w_sys_tmp2800 = 32'sh00000117;
	assign w_sys_tmp2805 = (w_sys_tmp2806 + r_run_k_29);
	assign w_sys_tmp2806 = 32'sh00000136;
	assign w_sys_tmp2811 = (w_sys_tmp2812 + r_run_k_29);
	assign w_sys_tmp2812 = 32'sh00000155;
	assign w_sys_tmp2817 = (w_sys_tmp2818 + r_run_k_29);
	assign w_sys_tmp2818 = 32'sh00000174;
	assign w_sys_tmp2823 = (w_sys_tmp2824 + r_run_k_29);
	assign w_sys_tmp2824 = 32'sh00000193;
	assign w_sys_tmp2829 = (w_sys_tmp2830 + r_run_k_29);
	assign w_sys_tmp2830 = 32'sh000001b2;
	assign w_sys_tmp2847 = (w_sys_tmp2848 + r_run_k_29);
	assign w_sys_tmp2848 = 32'sh000001d1;
	assign w_sys_tmp2853 = (w_sys_tmp2854 + r_run_k_29);
	assign w_sys_tmp2854 = 32'sh000001f0;
	assign w_sys_tmp2859 = (w_sys_tmp2860 + r_run_k_29);
	assign w_sys_tmp2860 = 32'sh0000020f;
	assign w_sys_tmp2865 = (w_sys_tmp2866 + r_run_k_29);
	assign w_sys_tmp2866 = 32'sh0000022e;
	assign w_sys_tmp2871 = (w_sys_tmp2872 + r_run_k_29);
	assign w_sys_tmp2872 = 32'sh0000024d;
	assign w_sys_tmp2877 = (w_sys_tmp2878 + r_run_k_29);
	assign w_sys_tmp2878 = 32'sh0000026c;
	assign w_sys_tmp2895 = (w_sys_tmp2896 + r_run_k_29);
	assign w_sys_tmp2896 = 32'sh0000028b;
	assign w_sys_tmp2901 = (w_sys_tmp2902 + r_run_k_29);
	assign w_sys_tmp2902 = 32'sh000002aa;
	assign w_sys_tmp2907 = (w_sys_tmp2908 + r_run_k_29);
	assign w_sys_tmp2908 = 32'sh000002c9;
	assign w_sys_tmp2913 = (w_sys_tmp2914 + r_run_k_29);
	assign w_sys_tmp2914 = 32'sh000002e8;
	assign w_sys_tmp2919 = (w_sys_tmp2920 + r_run_k_29);
	assign w_sys_tmp2920 = 32'sh00000307;
	assign w_sys_tmp2925 = (w_sys_tmp2926 + r_run_k_29);
	assign w_sys_tmp2926 = 32'sh00000326;
	assign w_sys_tmp2943 = (w_sys_tmp2944 + r_run_k_29);
	assign w_sys_tmp2944 = 32'sh00000345;
	assign w_sys_tmp2949 = (w_sys_tmp2950 + r_run_k_29);
	assign w_sys_tmp2950 = 32'sh00000364;
	assign w_sys_tmp2955 = (w_sys_tmp2956 + r_run_k_29);
	assign w_sys_tmp2956 = 32'sh00000383;
	assign w_sys_tmp2961 = (w_sys_tmp2962 + r_run_k_29);
	assign w_sys_tmp2962 = 32'sh000003a2;
	assign w_sys_tmp2967 = (w_sys_tmp2968 + r_run_k_29);
	assign w_sys_tmp2968 = 32'sh000003c1;
	assign w_sys_tmp2973 = (w_sys_tmp2974 + r_run_k_29);
	assign w_sys_tmp2974 = 32'sh00000025;
	assign w_sys_tmp2979 = (w_sys_tmp2980 + r_run_k_29);
	assign w_sys_tmp2980 = 32'sh00000044;
	assign w_sys_tmp2985 = (w_sys_tmp2986 + r_run_k_29);
	assign w_sys_tmp2986 = 32'sh00000063;
	assign w_sys_tmp2991 = (w_sys_tmp2992 + r_run_k_29);
	assign w_sys_tmp2992 = 32'sh00000082;
	assign w_sys_tmp2997 = (w_sys_tmp2998 + r_run_k_29);
	assign w_sys_tmp2998 = 32'sh000000a1;
	assign w_sys_tmp3003 = (w_sys_tmp3004 + r_run_k_29);
	assign w_sys_tmp3004 = 32'sh000000c0;
	assign w_sys_tmp3009 = (w_sys_tmp3010 + r_run_k_29);
	assign w_sys_tmp3010 = 32'sh000000df;
	assign w_sys_tmp3015 = (w_sys_tmp3016 + r_run_k_29);
	assign w_sys_tmp3016 = 32'sh000000fe;
	assign w_sys_tmp3033 = (w_sys_tmp3034 + r_run_k_29);
	assign w_sys_tmp3034 = 32'sh0000011d;
	assign w_sys_tmp3039 = (w_sys_tmp3040 + r_run_k_29);
	assign w_sys_tmp3040 = 32'sh0000013c;
	assign w_sys_tmp3045 = (w_sys_tmp3046 + r_run_k_29);
	assign w_sys_tmp3046 = 32'sh0000015b;
	assign w_sys_tmp3051 = (w_sys_tmp3052 + r_run_k_29);
	assign w_sys_tmp3052 = 32'sh0000017a;
	assign w_sys_tmp3057 = (w_sys_tmp3058 + r_run_k_29);
	assign w_sys_tmp3058 = 32'sh00000199;
	assign w_sys_tmp3063 = (w_sys_tmp3064 + r_run_k_29);
	assign w_sys_tmp3064 = 32'sh000001b8;
	assign w_sys_tmp3081 = (w_sys_tmp3082 + r_run_k_29);
	assign w_sys_tmp3082 = 32'sh000001d7;
	assign w_sys_tmp3087 = (w_sys_tmp3088 + r_run_k_29);
	assign w_sys_tmp3088 = 32'sh000001f6;
	assign w_sys_tmp3093 = (w_sys_tmp3094 + r_run_k_29);
	assign w_sys_tmp3094 = 32'sh00000215;
	assign w_sys_tmp3099 = (w_sys_tmp3100 + r_run_k_29);
	assign w_sys_tmp3100 = 32'sh00000234;
	assign w_sys_tmp3105 = (w_sys_tmp3106 + r_run_k_29);
	assign w_sys_tmp3106 = 32'sh00000253;
	assign w_sys_tmp3111 = (w_sys_tmp3112 + r_run_k_29);
	assign w_sys_tmp3112 = 32'sh00000272;
	assign w_sys_tmp3129 = (w_sys_tmp3130 + r_run_k_29);
	assign w_sys_tmp3130 = 32'sh00000291;
	assign w_sys_tmp3135 = (w_sys_tmp3136 + r_run_k_29);
	assign w_sys_tmp3136 = 32'sh000002b0;
	assign w_sys_tmp3141 = (w_sys_tmp3142 + r_run_k_29);
	assign w_sys_tmp3142 = 32'sh000002cf;
	assign w_sys_tmp3147 = (w_sys_tmp3148 + r_run_k_29);
	assign w_sys_tmp3148 = 32'sh000002ee;
	assign w_sys_tmp3153 = (w_sys_tmp3154 + r_run_k_29);
	assign w_sys_tmp3154 = 32'sh0000030d;
	assign w_sys_tmp3159 = (w_sys_tmp3160 + r_run_k_29);
	assign w_sys_tmp3160 = 32'sh0000032c;
	assign w_sys_tmp3177 = (w_sys_tmp3178 + r_run_k_29);
	assign w_sys_tmp3178 = 32'sh0000034b;
	assign w_sys_tmp3183 = (w_sys_tmp3184 + r_run_k_29);
	assign w_sys_tmp3184 = 32'sh0000036a;
	assign w_sys_tmp3189 = (w_sys_tmp3190 + r_run_k_29);
	assign w_sys_tmp3190 = 32'sh00000389;
	assign w_sys_tmp3195 = (w_sys_tmp3196 + r_run_k_29);
	assign w_sys_tmp3196 = 32'sh000003a8;
	assign w_sys_tmp3201 = (w_sys_tmp3202 + r_run_k_29);
	assign w_sys_tmp3202 = 32'sh000003c7;
	assign w_sys_tmp3207 = (w_sys_tmp3208 + r_run_k_29);
	assign w_sys_tmp3208 = 32'sh0000002b;
	assign w_sys_tmp3213 = (w_sys_tmp3214 + r_run_k_29);
	assign w_sys_tmp3214 = 32'sh0000004a;
	assign w_sys_tmp3219 = (w_sys_tmp3220 + r_run_k_29);
	assign w_sys_tmp3220 = 32'sh00000069;
	assign w_sys_tmp3225 = (w_sys_tmp3226 + r_run_k_29);
	assign w_sys_tmp3226 = 32'sh00000088;
	assign w_sys_tmp3231 = (w_sys_tmp3232 + r_run_k_29);
	assign w_sys_tmp3232 = 32'sh000000a7;
	assign w_sys_tmp3237 = (w_sys_tmp3238 + r_run_k_29);
	assign w_sys_tmp3238 = 32'sh000000c6;
	assign w_sys_tmp3243 = (w_sys_tmp3244 + r_run_k_29);
	assign w_sys_tmp3244 = 32'sh000000e5;
	assign w_sys_tmp3249 = (w_sys_tmp3250 + r_run_k_29);
	assign w_sys_tmp3250 = 32'sh00000104;
	assign w_sys_tmp3267 = (w_sys_tmp3268 + r_run_k_29);
	assign w_sys_tmp3268 = 32'sh00000123;
	assign w_sys_tmp3273 = (w_sys_tmp3274 + r_run_k_29);
	assign w_sys_tmp3274 = 32'sh00000142;
	assign w_sys_tmp3279 = (w_sys_tmp3280 + r_run_k_29);
	assign w_sys_tmp3280 = 32'sh00000161;
	assign w_sys_tmp3285 = (w_sys_tmp3286 + r_run_k_29);
	assign w_sys_tmp3286 = 32'sh00000180;
	assign w_sys_tmp3291 = (w_sys_tmp3292 + r_run_k_29);
	assign w_sys_tmp3292 = 32'sh0000019f;
	assign w_sys_tmp3297 = (w_sys_tmp3298 + r_run_k_29);
	assign w_sys_tmp3298 = 32'sh000001be;
	assign w_sys_tmp3315 = (w_sys_tmp3316 + r_run_k_29);
	assign w_sys_tmp3316 = 32'sh000001dd;
	assign w_sys_tmp3321 = (w_sys_tmp3322 + r_run_k_29);
	assign w_sys_tmp3322 = 32'sh000001fc;
	assign w_sys_tmp3327 = (w_sys_tmp3328 + r_run_k_29);
	assign w_sys_tmp3328 = 32'sh0000021b;
	assign w_sys_tmp3333 = (w_sys_tmp3334 + r_run_k_29);
	assign w_sys_tmp3334 = 32'sh0000023a;
	assign w_sys_tmp3339 = (w_sys_tmp3340 + r_run_k_29);
	assign w_sys_tmp3340 = 32'sh00000259;
	assign w_sys_tmp3345 = (w_sys_tmp3346 + r_run_k_29);
	assign w_sys_tmp3346 = 32'sh00000278;
	assign w_sys_tmp3363 = (w_sys_tmp3364 + r_run_k_29);
	assign w_sys_tmp3364 = 32'sh00000297;
	assign w_sys_tmp3369 = (w_sys_tmp3370 + r_run_k_29);
	assign w_sys_tmp3370 = 32'sh000002b6;
	assign w_sys_tmp3375 = (w_sys_tmp3376 + r_run_k_29);
	assign w_sys_tmp3376 = 32'sh000002d5;
	assign w_sys_tmp3381 = (w_sys_tmp3382 + r_run_k_29);
	assign w_sys_tmp3382 = 32'sh000002f4;
	assign w_sys_tmp3387 = (w_sys_tmp3388 + r_run_k_29);
	assign w_sys_tmp3388 = 32'sh00000313;
	assign w_sys_tmp3393 = (w_sys_tmp3394 + r_run_k_29);
	assign w_sys_tmp3394 = 32'sh00000332;
	assign w_sys_tmp3411 = (w_sys_tmp3412 + r_run_k_29);
	assign w_sys_tmp3412 = 32'sh00000351;
	assign w_sys_tmp3417 = (w_sys_tmp3418 + r_run_k_29);
	assign w_sys_tmp3418 = 32'sh00000370;
	assign w_sys_tmp3423 = (w_sys_tmp3424 + r_run_k_29);
	assign w_sys_tmp3424 = 32'sh0000038f;
	assign w_sys_tmp3429 = (w_sys_tmp3430 + r_run_k_29);
	assign w_sys_tmp3430 = 32'sh000003ae;
	assign w_sys_tmp3435 = (w_sys_tmp3436 + r_run_k_29);
	assign w_sys_tmp3436 = 32'sh000003cd;
	assign w_sys_tmp3441 = (w_sys_tmp3442 + r_run_k_29);
	assign w_sys_tmp3442 = 32'sh00000031;
	assign w_sys_tmp3447 = (w_sys_tmp3448 + r_run_k_29);
	assign w_sys_tmp3448 = 32'sh00000050;
	assign w_sys_tmp3453 = (w_sys_tmp3454 + r_run_k_29);
	assign w_sys_tmp3454 = 32'sh0000006f;
	assign w_sys_tmp3459 = (w_sys_tmp3460 + r_run_k_29);
	assign w_sys_tmp3460 = 32'sh0000008e;
	assign w_sys_tmp3465 = (w_sys_tmp3466 + r_run_k_29);
	assign w_sys_tmp3466 = 32'sh000000ad;
	assign w_sys_tmp3471 = (w_sys_tmp3472 + r_run_k_29);
	assign w_sys_tmp3472 = 32'sh000000cc;
	assign w_sys_tmp3477 = (w_sys_tmp3478 + r_run_k_29);
	assign w_sys_tmp3478 = 32'sh000000eb;
	assign w_sys_tmp3483 = (w_sys_tmp3484 + r_run_k_29);
	assign w_sys_tmp3484 = 32'sh0000010a;
	assign w_sys_tmp3501 = (w_sys_tmp3502 + r_run_k_29);
	assign w_sys_tmp3502 = 32'sh00000129;
	assign w_sys_tmp3507 = (w_sys_tmp3508 + r_run_k_29);
	assign w_sys_tmp3508 = 32'sh00000148;
	assign w_sys_tmp3513 = (w_sys_tmp3514 + r_run_k_29);
	assign w_sys_tmp3514 = 32'sh00000167;
	assign w_sys_tmp3519 = (w_sys_tmp3520 + r_run_k_29);
	assign w_sys_tmp3520 = 32'sh00000186;
	assign w_sys_tmp3525 = (w_sys_tmp3526 + r_run_k_29);
	assign w_sys_tmp3526 = 32'sh000001a5;
	assign w_sys_tmp3531 = (w_sys_tmp3532 + r_run_k_29);
	assign w_sys_tmp3532 = 32'sh000001c4;
	assign w_sys_tmp3549 = (w_sys_tmp3550 + r_run_k_29);
	assign w_sys_tmp3550 = 32'sh000001e3;
	assign w_sys_tmp3555 = (w_sys_tmp3556 + r_run_k_29);
	assign w_sys_tmp3556 = 32'sh00000202;
	assign w_sys_tmp3561 = (w_sys_tmp3562 + r_run_k_29);
	assign w_sys_tmp3562 = 32'sh00000221;
	assign w_sys_tmp3567 = (w_sys_tmp3568 + r_run_k_29);
	assign w_sys_tmp3568 = 32'sh00000240;
	assign w_sys_tmp3573 = (w_sys_tmp3574 + r_run_k_29);
	assign w_sys_tmp3574 = 32'sh0000025f;
	assign w_sys_tmp3579 = (w_sys_tmp3580 + r_run_k_29);
	assign w_sys_tmp3580 = 32'sh0000027e;
	assign w_sys_tmp3597 = (w_sys_tmp3598 + r_run_k_29);
	assign w_sys_tmp3598 = 32'sh0000029d;
	assign w_sys_tmp3603 = (w_sys_tmp3604 + r_run_k_29);
	assign w_sys_tmp3604 = 32'sh000002bc;
	assign w_sys_tmp3609 = (w_sys_tmp3610 + r_run_k_29);
	assign w_sys_tmp3610 = 32'sh000002db;
	assign w_sys_tmp3615 = (w_sys_tmp3616 + r_run_k_29);
	assign w_sys_tmp3616 = 32'sh000002fa;
	assign w_sys_tmp3621 = (w_sys_tmp3622 + r_run_k_29);
	assign w_sys_tmp3622 = 32'sh00000319;
	assign w_sys_tmp3627 = (w_sys_tmp3628 + r_run_k_29);
	assign w_sys_tmp3628 = 32'sh00000338;
	assign w_sys_tmp3645 = (w_sys_tmp3646 + r_run_k_29);
	assign w_sys_tmp3646 = 32'sh00000357;
	assign w_sys_tmp3651 = (w_sys_tmp3652 + r_run_k_29);
	assign w_sys_tmp3652 = 32'sh00000376;
	assign w_sys_tmp3657 = (w_sys_tmp3658 + r_run_k_29);
	assign w_sys_tmp3658 = 32'sh00000395;
	assign w_sys_tmp3663 = (w_sys_tmp3664 + r_run_k_29);
	assign w_sys_tmp3664 = 32'sh000003b4;
	assign w_sys_tmp3669 = (w_sys_tmp3670 + r_run_k_29);
	assign w_sys_tmp3670 = 32'sh000003d3;
	assign w_sys_tmp3674 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp3675 = 32'sh00000019;
	assign w_sys_tmp3676 = ( !w_sys_tmp3677 );
	assign w_sys_tmp3677 = (w_sys_tmp3678 < r_run_k_29);
	assign w_sys_tmp3678 = 32'sh0000001f;
	assign w_sys_tmp3681 = (w_sys_tmp3682 + r_run_k_29);
	assign w_sys_tmp3682 = 32'sh0000001f;
	assign w_sys_tmp3683 = w_fld_T_0_dataout_1;
	assign w_sys_tmp3687 = (w_sys_tmp3688 + r_run_k_29);
	assign w_sys_tmp3688 = 32'sh0000003e;
	assign w_sys_tmp3693 = (w_sys_tmp3694 + r_run_k_29);
	assign w_sys_tmp3694 = 32'sh0000005d;
	assign w_sys_tmp3699 = (w_sys_tmp3700 + r_run_k_29);
	assign w_sys_tmp3700 = 32'sh0000007c;
	assign w_sys_tmp3705 = (w_sys_tmp3706 + r_run_k_29);
	assign w_sys_tmp3706 = 32'sh0000009b;
	assign w_sys_tmp3711 = (w_sys_tmp3712 + r_run_k_29);
	assign w_sys_tmp3712 = 32'sh000000ba;
	assign w_sys_tmp3717 = (w_sys_tmp3718 + r_run_k_29);
	assign w_sys_tmp3718 = 32'sh000000d9;
	assign w_sys_tmp3723 = (w_sys_tmp3724 + r_run_k_29);
	assign w_sys_tmp3724 = 32'sh000000f8;
	assign w_sys_tmp3741 = (w_sys_tmp3742 + r_run_k_29);
	assign w_sys_tmp3742 = 32'sh00000117;
	assign w_sys_tmp3747 = (w_sys_tmp3748 + r_run_k_29);
	assign w_sys_tmp3748 = 32'sh00000136;
	assign w_sys_tmp3753 = (w_sys_tmp3754 + r_run_k_29);
	assign w_sys_tmp3754 = 32'sh00000155;
	assign w_sys_tmp3759 = (w_sys_tmp3760 + r_run_k_29);
	assign w_sys_tmp3760 = 32'sh00000174;
	assign w_sys_tmp3765 = (w_sys_tmp3766 + r_run_k_29);
	assign w_sys_tmp3766 = 32'sh00000193;
	assign w_sys_tmp3771 = (w_sys_tmp3772 + r_run_k_29);
	assign w_sys_tmp3772 = 32'sh000001b2;
	assign w_sys_tmp3789 = (w_sys_tmp3790 + r_run_k_29);
	assign w_sys_tmp3790 = 32'sh000001d1;
	assign w_sys_tmp3795 = (w_sys_tmp3796 + r_run_k_29);
	assign w_sys_tmp3796 = 32'sh000001f0;
	assign w_sys_tmp3801 = (w_sys_tmp3802 + r_run_k_29);
	assign w_sys_tmp3802 = 32'sh0000020f;
	assign w_sys_tmp3807 = (w_sys_tmp3808 + r_run_k_29);
	assign w_sys_tmp3808 = 32'sh0000022e;
	assign w_sys_tmp3813 = (w_sys_tmp3814 + r_run_k_29);
	assign w_sys_tmp3814 = 32'sh0000024d;
	assign w_sys_tmp3819 = (w_sys_tmp3820 + r_run_k_29);
	assign w_sys_tmp3820 = 32'sh0000026c;
	assign w_sys_tmp3837 = (w_sys_tmp3838 + r_run_k_29);
	assign w_sys_tmp3838 = 32'sh0000028b;
	assign w_sys_tmp3843 = (w_sys_tmp3844 + r_run_k_29);
	assign w_sys_tmp3844 = 32'sh000002aa;
	assign w_sys_tmp3849 = (w_sys_tmp3850 + r_run_k_29);
	assign w_sys_tmp3850 = 32'sh000002c9;
	assign w_sys_tmp3855 = (w_sys_tmp3856 + r_run_k_29);
	assign w_sys_tmp3856 = 32'sh000002e8;
	assign w_sys_tmp3861 = (w_sys_tmp3862 + r_run_k_29);
	assign w_sys_tmp3862 = 32'sh00000307;
	assign w_sys_tmp3867 = (w_sys_tmp3868 + r_run_k_29);
	assign w_sys_tmp3868 = 32'sh00000326;
	assign w_sys_tmp3885 = (w_sys_tmp3886 + r_run_k_29);
	assign w_sys_tmp3886 = 32'sh00000345;
	assign w_sys_tmp3891 = (w_sys_tmp3892 + r_run_k_29);
	assign w_sys_tmp3892 = 32'sh00000364;
	assign w_sys_tmp3897 = (w_sys_tmp3898 + r_run_k_29);
	assign w_sys_tmp3898 = 32'sh00000383;
	assign w_sys_tmp3903 = (w_sys_tmp3904 + r_run_k_29);
	assign w_sys_tmp3904 = 32'sh000003a2;
	assign w_sys_tmp3909 = (w_sys_tmp3910 + r_run_k_29);
	assign w_sys_tmp3910 = 32'sh000003c1;
	assign w_sys_tmp3914 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp3915 = 32'sh00000002;
	assign w_sys_tmp3916 = ( !w_sys_tmp3917 );
	assign w_sys_tmp3917 = (w_sys_tmp3918 < r_run_k_29);
	assign w_sys_tmp3918 = 32'sh00000007;
	assign w_sys_tmp3921 = (w_sys_tmp3922 + r_run_k_29);
	assign w_sys_tmp3922 = 32'sh0000003e;
	assign w_sys_tmp3923 = w_sub00_result_dataout;
	assign w_sys_tmp3927 = (w_sys_tmp3928 + r_run_k_29);
	assign w_sys_tmp3928 = 32'sh0000005d;
	assign w_sys_tmp3933 = (w_sys_tmp3934 + r_run_k_29);
	assign w_sys_tmp3934 = 32'sh0000007c;
	assign w_sys_tmp3939 = (w_sys_tmp3940 + r_run_k_29);
	assign w_sys_tmp3940 = 32'sh0000009b;
	assign w_sys_tmp3945 = (w_sys_tmp3946 + r_run_k_29);
	assign w_sys_tmp3946 = 32'sh000000ba;
	assign w_sys_tmp3951 = (w_sys_tmp3952 + r_run_k_29);
	assign w_sys_tmp3952 = 32'sh000000d9;
	assign w_sys_tmp3957 = (w_sys_tmp3958 + r_run_k_29);
	assign w_sys_tmp3958 = 32'sh000000f8;
	assign w_sys_tmp3962 = (w_sys_tmp3963 + r_run_k_29);
	assign w_sys_tmp3963 = 32'sh00000117;
	assign w_sys_tmp3967 = (w_sys_tmp3968 + r_run_k_29);
	assign w_sys_tmp3968 = 32'sh00000136;
	assign w_sys_tmp3972 = (w_sys_tmp3973 + r_run_k_29);
	assign w_sys_tmp3973 = 32'sh00000155;
	assign w_sys_tmp3977 = (w_sys_tmp3978 + r_run_k_29);
	assign w_sys_tmp3978 = 32'sh00000174;
	assign w_sys_tmp3982 = (w_sys_tmp3983 + r_run_k_29);
	assign w_sys_tmp3983 = 32'sh00000193;
	assign w_sys_tmp3987 = (w_sys_tmp3988 + r_run_k_29);
	assign w_sys_tmp3988 = 32'sh000001b2;
	assign w_sys_tmp3992 = (w_sys_tmp3993 + r_run_k_29);
	assign w_sys_tmp3993 = 32'sh000001d1;
	assign w_sys_tmp3997 = (w_sys_tmp3998 + r_run_k_29);
	assign w_sys_tmp3998 = 32'sh000001f0;
	assign w_sys_tmp4002 = (w_sys_tmp4003 + r_run_k_29);
	assign w_sys_tmp4003 = 32'sh0000020f;
	assign w_sys_tmp4007 = (w_sys_tmp4008 + r_run_k_29);
	assign w_sys_tmp4008 = 32'sh0000022e;
	assign w_sys_tmp4012 = (w_sys_tmp4013 + r_run_k_29);
	assign w_sys_tmp4013 = 32'sh0000024d;
	assign w_sys_tmp4017 = (w_sys_tmp4018 + r_run_k_29);
	assign w_sys_tmp4018 = 32'sh0000026c;
	assign w_sys_tmp4022 = (w_sys_tmp4023 + r_run_k_29);
	assign w_sys_tmp4023 = 32'sh0000028b;
	assign w_sys_tmp4027 = (w_sys_tmp4028 + r_run_k_29);
	assign w_sys_tmp4028 = 32'sh000002aa;
	assign w_sys_tmp4032 = (w_sys_tmp4033 + r_run_k_29);
	assign w_sys_tmp4033 = 32'sh000002c9;
	assign w_sys_tmp4037 = (w_sys_tmp4038 + r_run_k_29);
	assign w_sys_tmp4038 = 32'sh000002e8;
	assign w_sys_tmp4042 = (w_sys_tmp4043 + r_run_k_29);
	assign w_sys_tmp4043 = 32'sh00000307;
	assign w_sys_tmp4047 = (w_sys_tmp4048 + r_run_k_29);
	assign w_sys_tmp4048 = 32'sh00000326;
	assign w_sys_tmp4052 = (w_sys_tmp4053 + r_run_k_29);
	assign w_sys_tmp4053 = 32'sh00000345;
	assign w_sys_tmp4057 = (w_sys_tmp4058 + r_run_k_29);
	assign w_sys_tmp4058 = 32'sh00000364;
	assign w_sys_tmp4062 = (w_sys_tmp4063 + r_run_k_29);
	assign w_sys_tmp4063 = 32'sh00000383;
	assign w_sys_tmp4067 = (w_sys_tmp4068 + r_run_k_29);
	assign w_sys_tmp4068 = 32'sh000003a2;
	assign w_sys_tmp4072 = (w_sys_tmp4073 + r_run_k_29);
	assign w_sys_tmp4073 = 32'sh00000044;
	assign w_sys_tmp4077 = (w_sys_tmp4078 + r_run_k_29);
	assign w_sys_tmp4078 = 32'sh00000063;
	assign w_sys_tmp4082 = (w_sys_tmp4083 + r_run_k_29);
	assign w_sys_tmp4083 = 32'sh00000082;
	assign w_sys_tmp4087 = (w_sys_tmp4088 + r_run_k_29);
	assign w_sys_tmp4088 = 32'sh000000a1;
	assign w_sys_tmp4092 = (w_sys_tmp4093 + r_run_k_29);
	assign w_sys_tmp4093 = 32'sh000000c0;
	assign w_sys_tmp4097 = (w_sys_tmp4098 + r_run_k_29);
	assign w_sys_tmp4098 = 32'sh000000df;
	assign w_sys_tmp4102 = (w_sys_tmp4103 + r_run_k_29);
	assign w_sys_tmp4103 = 32'sh000000fe;
	assign w_sys_tmp4107 = (w_sys_tmp4108 + r_run_k_29);
	assign w_sys_tmp4108 = 32'sh0000011d;
	assign w_sys_tmp4112 = (w_sys_tmp4113 + r_run_k_29);
	assign w_sys_tmp4113 = 32'sh0000013c;
	assign w_sys_tmp4117 = (w_sys_tmp4118 + r_run_k_29);
	assign w_sys_tmp4118 = 32'sh0000015b;
	assign w_sys_tmp4122 = (w_sys_tmp4123 + r_run_k_29);
	assign w_sys_tmp4123 = 32'sh0000017a;
	assign w_sys_tmp4127 = (w_sys_tmp4128 + r_run_k_29);
	assign w_sys_tmp4128 = 32'sh00000199;
	assign w_sys_tmp4132 = (w_sys_tmp4133 + r_run_k_29);
	assign w_sys_tmp4133 = 32'sh000001b8;
	assign w_sys_tmp4137 = (w_sys_tmp4138 + r_run_k_29);
	assign w_sys_tmp4138 = 32'sh000001d7;
	assign w_sys_tmp4142 = (w_sys_tmp4143 + r_run_k_29);
	assign w_sys_tmp4143 = 32'sh000001f6;
	assign w_sys_tmp4147 = (w_sys_tmp4148 + r_run_k_29);
	assign w_sys_tmp4148 = 32'sh00000215;
	assign w_sys_tmp4152 = (w_sys_tmp4153 + r_run_k_29);
	assign w_sys_tmp4153 = 32'sh00000234;
	assign w_sys_tmp4157 = (w_sys_tmp4158 + r_run_k_29);
	assign w_sys_tmp4158 = 32'sh00000253;
	assign w_sys_tmp4162 = (w_sys_tmp4163 + r_run_k_29);
	assign w_sys_tmp4163 = 32'sh00000272;
	assign w_sys_tmp4167 = (w_sys_tmp4168 + r_run_k_29);
	assign w_sys_tmp4168 = 32'sh00000291;
	assign w_sys_tmp4172 = (w_sys_tmp4173 + r_run_k_29);
	assign w_sys_tmp4173 = 32'sh000002b0;
	assign w_sys_tmp4177 = (w_sys_tmp4178 + r_run_k_29);
	assign w_sys_tmp4178 = 32'sh000002cf;
	assign w_sys_tmp4182 = (w_sys_tmp4183 + r_run_k_29);
	assign w_sys_tmp4183 = 32'sh000002ee;
	assign w_sys_tmp4187 = (w_sys_tmp4188 + r_run_k_29);
	assign w_sys_tmp4188 = 32'sh0000030d;
	assign w_sys_tmp4192 = (w_sys_tmp4193 + r_run_k_29);
	assign w_sys_tmp4193 = 32'sh0000032c;
	assign w_sys_tmp4197 = (w_sys_tmp4198 + r_run_k_29);
	assign w_sys_tmp4198 = 32'sh0000034b;
	assign w_sys_tmp4202 = (w_sys_tmp4203 + r_run_k_29);
	assign w_sys_tmp4203 = 32'sh0000036a;
	assign w_sys_tmp4207 = (w_sys_tmp4208 + r_run_k_29);
	assign w_sys_tmp4208 = 32'sh00000389;
	assign w_sys_tmp4212 = (w_sys_tmp4213 + r_run_k_29);
	assign w_sys_tmp4213 = 32'sh000003a8;
	assign w_sys_tmp4217 = (w_sys_tmp4218 + r_run_k_29);
	assign w_sys_tmp4218 = 32'sh0000004a;
	assign w_sys_tmp4222 = (w_sys_tmp4223 + r_run_k_29);
	assign w_sys_tmp4223 = 32'sh00000069;
	assign w_sys_tmp4227 = (w_sys_tmp4228 + r_run_k_29);
	assign w_sys_tmp4228 = 32'sh00000088;
	assign w_sys_tmp4232 = (w_sys_tmp4233 + r_run_k_29);
	assign w_sys_tmp4233 = 32'sh000000a7;
	assign w_sys_tmp4237 = (w_sys_tmp4238 + r_run_k_29);
	assign w_sys_tmp4238 = 32'sh000000c6;
	assign w_sys_tmp4242 = (w_sys_tmp4243 + r_run_k_29);
	assign w_sys_tmp4243 = 32'sh000000e5;
	assign w_sys_tmp4247 = (w_sys_tmp4248 + r_run_k_29);
	assign w_sys_tmp4248 = 32'sh00000104;
	assign w_sys_tmp4252 = (w_sys_tmp4253 + r_run_k_29);
	assign w_sys_tmp4253 = 32'sh00000123;
	assign w_sys_tmp4257 = (w_sys_tmp4258 + r_run_k_29);
	assign w_sys_tmp4258 = 32'sh00000142;
	assign w_sys_tmp4262 = (w_sys_tmp4263 + r_run_k_29);
	assign w_sys_tmp4263 = 32'sh00000161;
	assign w_sys_tmp4267 = (w_sys_tmp4268 + r_run_k_29);
	assign w_sys_tmp4268 = 32'sh00000180;
	assign w_sys_tmp4272 = (w_sys_tmp4273 + r_run_k_29);
	assign w_sys_tmp4273 = 32'sh0000019f;
	assign w_sys_tmp4277 = (w_sys_tmp4278 + r_run_k_29);
	assign w_sys_tmp4278 = 32'sh000001be;
	assign w_sys_tmp4282 = (w_sys_tmp4283 + r_run_k_29);
	assign w_sys_tmp4283 = 32'sh000001dd;
	assign w_sys_tmp4287 = (w_sys_tmp4288 + r_run_k_29);
	assign w_sys_tmp4288 = 32'sh000001fc;
	assign w_sys_tmp4292 = (w_sys_tmp4293 + r_run_k_29);
	assign w_sys_tmp4293 = 32'sh0000021b;
	assign w_sys_tmp4297 = (w_sys_tmp4298 + r_run_k_29);
	assign w_sys_tmp4298 = 32'sh0000023a;
	assign w_sys_tmp4302 = (w_sys_tmp4303 + r_run_k_29);
	assign w_sys_tmp4303 = 32'sh00000259;
	assign w_sys_tmp4307 = (w_sys_tmp4308 + r_run_k_29);
	assign w_sys_tmp4308 = 32'sh00000278;
	assign w_sys_tmp4312 = (w_sys_tmp4313 + r_run_k_29);
	assign w_sys_tmp4313 = 32'sh00000297;
	assign w_sys_tmp4317 = (w_sys_tmp4318 + r_run_k_29);
	assign w_sys_tmp4318 = 32'sh000002b6;
	assign w_sys_tmp4322 = (w_sys_tmp4323 + r_run_k_29);
	assign w_sys_tmp4323 = 32'sh000002d5;
	assign w_sys_tmp4327 = (w_sys_tmp4328 + r_run_k_29);
	assign w_sys_tmp4328 = 32'sh000002f4;
	assign w_sys_tmp4332 = (w_sys_tmp4333 + r_run_k_29);
	assign w_sys_tmp4333 = 32'sh00000313;
	assign w_sys_tmp4337 = (w_sys_tmp4338 + r_run_k_29);
	assign w_sys_tmp4338 = 32'sh00000332;
	assign w_sys_tmp4342 = (w_sys_tmp4343 + r_run_k_29);
	assign w_sys_tmp4343 = 32'sh00000351;
	assign w_sys_tmp4347 = (w_sys_tmp4348 + r_run_k_29);
	assign w_sys_tmp4348 = 32'sh00000370;
	assign w_sys_tmp4352 = (w_sys_tmp4353 + r_run_k_29);
	assign w_sys_tmp4353 = 32'sh0000038f;
	assign w_sys_tmp4357 = (w_sys_tmp4358 + r_run_k_29);
	assign w_sys_tmp4358 = 32'sh000003ae;
	assign w_sys_tmp4362 = (w_sys_tmp4363 + r_run_k_29);
	assign w_sys_tmp4363 = 32'sh00000050;
	assign w_sys_tmp4367 = (w_sys_tmp4368 + r_run_k_29);
	assign w_sys_tmp4368 = 32'sh0000006f;
	assign w_sys_tmp4372 = (w_sys_tmp4373 + r_run_k_29);
	assign w_sys_tmp4373 = 32'sh0000008e;
	assign w_sys_tmp4377 = (w_sys_tmp4378 + r_run_k_29);
	assign w_sys_tmp4378 = 32'sh000000ad;
	assign w_sys_tmp4382 = (w_sys_tmp4383 + r_run_k_29);
	assign w_sys_tmp4383 = 32'sh000000cc;
	assign w_sys_tmp4387 = (w_sys_tmp4388 + r_run_k_29);
	assign w_sys_tmp4388 = 32'sh000000eb;
	assign w_sys_tmp4392 = (w_sys_tmp4393 + r_run_k_29);
	assign w_sys_tmp4393 = 32'sh0000010a;
	assign w_sys_tmp4397 = (w_sys_tmp4398 + r_run_k_29);
	assign w_sys_tmp4398 = 32'sh00000129;
	assign w_sys_tmp4402 = (w_sys_tmp4403 + r_run_k_29);
	assign w_sys_tmp4403 = 32'sh00000148;
	assign w_sys_tmp4407 = (w_sys_tmp4408 + r_run_k_29);
	assign w_sys_tmp4408 = 32'sh00000167;
	assign w_sys_tmp4412 = (w_sys_tmp4413 + r_run_k_29);
	assign w_sys_tmp4413 = 32'sh00000186;
	assign w_sys_tmp4417 = (w_sys_tmp4418 + r_run_k_29);
	assign w_sys_tmp4418 = 32'sh000001a5;
	assign w_sys_tmp4422 = (w_sys_tmp4423 + r_run_k_29);
	assign w_sys_tmp4423 = 32'sh000001c4;
	assign w_sys_tmp4427 = (w_sys_tmp4428 + r_run_k_29);
	assign w_sys_tmp4428 = 32'sh000001e3;
	assign w_sys_tmp4432 = (w_sys_tmp4433 + r_run_k_29);
	assign w_sys_tmp4433 = 32'sh00000202;
	assign w_sys_tmp4437 = (w_sys_tmp4438 + r_run_k_29);
	assign w_sys_tmp4438 = 32'sh00000221;
	assign w_sys_tmp4442 = (w_sys_tmp4443 + r_run_k_29);
	assign w_sys_tmp4443 = 32'sh00000240;
	assign w_sys_tmp4447 = (w_sys_tmp4448 + r_run_k_29);
	assign w_sys_tmp4448 = 32'sh0000025f;
	assign w_sys_tmp4452 = (w_sys_tmp4453 + r_run_k_29);
	assign w_sys_tmp4453 = 32'sh0000027e;
	assign w_sys_tmp4457 = (w_sys_tmp4458 + r_run_k_29);
	assign w_sys_tmp4458 = 32'sh0000029d;
	assign w_sys_tmp4462 = (w_sys_tmp4463 + r_run_k_29);
	assign w_sys_tmp4463 = 32'sh000002bc;
	assign w_sys_tmp4467 = (w_sys_tmp4468 + r_run_k_29);
	assign w_sys_tmp4468 = 32'sh000002db;
	assign w_sys_tmp4472 = (w_sys_tmp4473 + r_run_k_29);
	assign w_sys_tmp4473 = 32'sh000002fa;
	assign w_sys_tmp4477 = (w_sys_tmp4478 + r_run_k_29);
	assign w_sys_tmp4478 = 32'sh00000319;
	assign w_sys_tmp4482 = (w_sys_tmp4483 + r_run_k_29);
	assign w_sys_tmp4483 = 32'sh00000338;
	assign w_sys_tmp4487 = (w_sys_tmp4488 + r_run_k_29);
	assign w_sys_tmp4488 = 32'sh00000357;
	assign w_sys_tmp4492 = (w_sys_tmp4493 + r_run_k_29);
	assign w_sys_tmp4493 = 32'sh00000376;
	assign w_sys_tmp4497 = (w_sys_tmp4498 + r_run_k_29);
	assign w_sys_tmp4498 = 32'sh00000395;
	assign w_sys_tmp4502 = (w_sys_tmp4503 + r_run_k_29);
	assign w_sys_tmp4503 = 32'sh000003b4;
	assign w_sys_tmp4506 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp4507 = 32'sh0000001a;
	assign w_sys_tmp4508 = ( !w_sys_tmp4509 );
	assign w_sys_tmp4509 = (w_sys_tmp4510 < r_run_k_29);
	assign w_sys_tmp4510 = 32'sh0000001e;
	assign w_sys_tmp4513 = (w_sys_tmp4514 + r_run_k_29);
	assign w_sys_tmp4514 = 32'sh0000003e;
	assign w_sys_tmp4515 = w_sub20_result_dataout;
	assign w_sys_tmp4519 = (w_sys_tmp4520 + r_run_k_29);
	assign w_sys_tmp4520 = 32'sh0000005d;
	assign w_sys_tmp4525 = (w_sys_tmp4526 + r_run_k_29);
	assign w_sys_tmp4526 = 32'sh0000007c;
	assign w_sys_tmp4531 = (w_sys_tmp4532 + r_run_k_29);
	assign w_sys_tmp4532 = 32'sh0000009b;
	assign w_sys_tmp4537 = (w_sys_tmp4538 + r_run_k_29);
	assign w_sys_tmp4538 = 32'sh000000ba;
	assign w_sys_tmp4543 = (w_sys_tmp4544 + r_run_k_29);
	assign w_sys_tmp4544 = 32'sh000000d9;
	assign w_sys_tmp4549 = (w_sys_tmp4550 + r_run_k_29);
	assign w_sys_tmp4550 = 32'sh000000f8;
	assign w_sys_tmp4554 = (w_sys_tmp4555 + r_run_k_29);
	assign w_sys_tmp4555 = 32'sh00000117;
	assign w_sys_tmp4559 = (w_sys_tmp4560 + r_run_k_29);
	assign w_sys_tmp4560 = 32'sh00000136;
	assign w_sys_tmp4564 = (w_sys_tmp4565 + r_run_k_29);
	assign w_sys_tmp4565 = 32'sh00000155;
	assign w_sys_tmp4569 = (w_sys_tmp4570 + r_run_k_29);
	assign w_sys_tmp4570 = 32'sh00000174;
	assign w_sys_tmp4574 = (w_sys_tmp4575 + r_run_k_29);
	assign w_sys_tmp4575 = 32'sh00000193;
	assign w_sys_tmp4579 = (w_sys_tmp4580 + r_run_k_29);
	assign w_sys_tmp4580 = 32'sh000001b2;
	assign w_sys_tmp4584 = (w_sys_tmp4585 + r_run_k_29);
	assign w_sys_tmp4585 = 32'sh000001d1;
	assign w_sys_tmp4589 = (w_sys_tmp4590 + r_run_k_29);
	assign w_sys_tmp4590 = 32'sh000001f0;
	assign w_sys_tmp4594 = (w_sys_tmp4595 + r_run_k_29);
	assign w_sys_tmp4595 = 32'sh0000020f;
	assign w_sys_tmp4599 = (w_sys_tmp4600 + r_run_k_29);
	assign w_sys_tmp4600 = 32'sh0000022e;
	assign w_sys_tmp4604 = (w_sys_tmp4605 + r_run_k_29);
	assign w_sys_tmp4605 = 32'sh0000024d;
	assign w_sys_tmp4609 = (w_sys_tmp4610 + r_run_k_29);
	assign w_sys_tmp4610 = 32'sh0000026c;
	assign w_sys_tmp4614 = (w_sys_tmp4615 + r_run_k_29);
	assign w_sys_tmp4615 = 32'sh0000028b;
	assign w_sys_tmp4619 = (w_sys_tmp4620 + r_run_k_29);
	assign w_sys_tmp4620 = 32'sh000002aa;
	assign w_sys_tmp4624 = (w_sys_tmp4625 + r_run_k_29);
	assign w_sys_tmp4625 = 32'sh000002c9;
	assign w_sys_tmp4629 = (w_sys_tmp4630 + r_run_k_29);
	assign w_sys_tmp4630 = 32'sh000002e8;
	assign w_sys_tmp4634 = (w_sys_tmp4635 + r_run_k_29);
	assign w_sys_tmp4635 = 32'sh00000307;
	assign w_sys_tmp4639 = (w_sys_tmp4640 + r_run_k_29);
	assign w_sys_tmp4640 = 32'sh00000326;
	assign w_sys_tmp4644 = (w_sys_tmp4645 + r_run_k_29);
	assign w_sys_tmp4645 = 32'sh00000345;
	assign w_sys_tmp4649 = (w_sys_tmp4650 + r_run_k_29);
	assign w_sys_tmp4650 = 32'sh00000364;
	assign w_sys_tmp4654 = (w_sys_tmp4655 + r_run_k_29);
	assign w_sys_tmp4655 = 32'sh00000383;
	assign w_sys_tmp4659 = (w_sys_tmp4660 + r_run_k_29);
	assign w_sys_tmp4660 = 32'sh000003a2;
	assign w_sys_tmp4663 = (r_run_k_29 + w_sys_intOne);


	sub19
		sub19_inst(
			.i_fld_T_0_addr_0 (w_sub19_T_addr),
			.i_fld_T_0_datain_0 (w_sub19_T_datain),
			.o_fld_T_0_dataout_0 (w_sub19_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub19_T_r_w),
			.i_fld_U_2_addr_0 (w_sub19_U_addr),
			.i_fld_U_2_datain_0 (w_sub19_U_datain),
			.o_fld_U_2_dataout_0 (w_sub19_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub19_U_r_w),
			.i_fld_V_1_addr_0 (w_sub19_V_addr),
			.i_fld_V_1_datain_0 (w_sub19_V_datain),
			.o_fld_V_1_dataout_0 (w_sub19_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub19_V_r_w),
			.i_fld_result_3_addr_0 (w_sub19_result_addr),
			.i_fld_result_3_datain_0 (w_sub19_result_datain),
			.o_fld_result_3_dataout_0 (w_sub19_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub19_result_r_w),
			.o_run_busy (w_sub19_run_busy),
			.i_run_req (r_sub19_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub09
		sub09_inst(
			.i_fld_T_0_addr_0 (w_sub09_T_addr),
			.i_fld_T_0_datain_0 (w_sub09_T_datain),
			.o_fld_T_0_dataout_0 (w_sub09_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub09_T_r_w),
			.i_fld_U_2_addr_0 (w_sub09_U_addr),
			.i_fld_U_2_datain_0 (w_sub09_U_datain),
			.o_fld_U_2_dataout_0 (w_sub09_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub09_U_r_w),
			.i_fld_V_1_addr_0 (w_sub09_V_addr),
			.i_fld_V_1_datain_0 (w_sub09_V_datain),
			.o_fld_V_1_dataout_0 (w_sub09_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub09_V_r_w),
			.i_fld_result_3_addr_0 (w_sub09_result_addr),
			.i_fld_result_3_datain_0 (w_sub09_result_datain),
			.o_fld_result_3_dataout_0 (w_sub09_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub09_result_r_w),
			.o_run_busy (w_sub09_run_busy),
			.i_run_req (r_sub09_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub08
		sub08_inst(
			.i_fld_T_0_addr_0 (w_sub08_T_addr),
			.i_fld_T_0_datain_0 (w_sub08_T_datain),
			.o_fld_T_0_dataout_0 (w_sub08_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub08_T_r_w),
			.i_fld_U_2_addr_0 (w_sub08_U_addr),
			.i_fld_U_2_datain_0 (w_sub08_U_datain),
			.o_fld_U_2_dataout_0 (w_sub08_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub08_U_r_w),
			.i_fld_V_1_addr_0 (w_sub08_V_addr),
			.i_fld_V_1_datain_0 (w_sub08_V_datain),
			.o_fld_V_1_dataout_0 (w_sub08_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub08_V_r_w),
			.i_fld_result_3_addr_0 (w_sub08_result_addr),
			.i_fld_result_3_datain_0 (w_sub08_result_datain),
			.o_fld_result_3_dataout_0 (w_sub08_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub08_result_r_w),
			.o_run_busy (w_sub08_run_busy),
			.i_run_req (r_sub08_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub24
		sub24_inst(
			.i_fld_T_0_addr_0 (w_sub24_T_addr),
			.i_fld_T_0_datain_0 (w_sub24_T_datain),
			.o_fld_T_0_dataout_0 (w_sub24_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub24_T_r_w),
			.i_fld_U_2_addr_0 (w_sub24_U_addr),
			.i_fld_U_2_datain_0 (w_sub24_U_datain),
			.o_fld_U_2_dataout_0 (w_sub24_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub24_U_r_w),
			.i_fld_V_1_addr_0 (w_sub24_V_addr),
			.i_fld_V_1_datain_0 (w_sub24_V_datain),
			.o_fld_V_1_dataout_0 (w_sub24_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub24_V_r_w),
			.i_fld_result_3_addr_0 (w_sub24_result_addr),
			.i_fld_result_3_datain_0 (w_sub24_result_datain),
			.o_fld_result_3_dataout_0 (w_sub24_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub24_result_r_w),
			.o_run_busy (w_sub24_run_busy),
			.i_run_req (r_sub24_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub22
		sub22_inst(
			.i_fld_T_0_addr_0 (w_sub22_T_addr),
			.i_fld_T_0_datain_0 (w_sub22_T_datain),
			.o_fld_T_0_dataout_0 (w_sub22_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub22_T_r_w),
			.i_fld_U_2_addr_0 (w_sub22_U_addr),
			.i_fld_U_2_datain_0 (w_sub22_U_datain),
			.o_fld_U_2_dataout_0 (w_sub22_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub22_U_r_w),
			.i_fld_V_1_addr_0 (w_sub22_V_addr),
			.i_fld_V_1_datain_0 (w_sub22_V_datain),
			.o_fld_V_1_dataout_0 (w_sub22_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub22_V_r_w),
			.i_fld_result_3_addr_0 (w_sub22_result_addr),
			.i_fld_result_3_datain_0 (w_sub22_result_datain),
			.o_fld_result_3_dataout_0 (w_sub22_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub22_result_r_w),
			.o_run_busy (w_sub22_run_busy),
			.i_run_req (r_sub22_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub23
		sub23_inst(
			.i_fld_T_0_addr_0 (w_sub23_T_addr),
			.i_fld_T_0_datain_0 (w_sub23_T_datain),
			.o_fld_T_0_dataout_0 (w_sub23_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub23_T_r_w),
			.i_fld_U_2_addr_0 (w_sub23_U_addr),
			.i_fld_U_2_datain_0 (w_sub23_U_datain),
			.o_fld_U_2_dataout_0 (w_sub23_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub23_U_r_w),
			.i_fld_V_1_addr_0 (w_sub23_V_addr),
			.i_fld_V_1_datain_0 (w_sub23_V_datain),
			.o_fld_V_1_dataout_0 (w_sub23_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub23_V_r_w),
			.i_fld_result_3_addr_0 (w_sub23_result_addr),
			.i_fld_result_3_datain_0 (w_sub23_result_datain),
			.o_fld_result_3_dataout_0 (w_sub23_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub23_result_r_w),
			.o_run_busy (w_sub23_run_busy),
			.i_run_req (r_sub23_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub12
		sub12_inst(
			.i_fld_T_0_addr_0 (w_sub12_T_addr),
			.i_fld_T_0_datain_0 (w_sub12_T_datain),
			.o_fld_T_0_dataout_0 (w_sub12_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub12_T_r_w),
			.i_fld_U_2_addr_0 (w_sub12_U_addr),
			.i_fld_U_2_datain_0 (w_sub12_U_datain),
			.o_fld_U_2_dataout_0 (w_sub12_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub12_U_r_w),
			.i_fld_V_1_addr_0 (w_sub12_V_addr),
			.i_fld_V_1_datain_0 (w_sub12_V_datain),
			.o_fld_V_1_dataout_0 (w_sub12_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub12_V_r_w),
			.i_fld_result_3_addr_0 (w_sub12_result_addr),
			.i_fld_result_3_datain_0 (w_sub12_result_datain),
			.o_fld_result_3_dataout_0 (w_sub12_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub12_result_r_w),
			.o_run_busy (w_sub12_run_busy),
			.i_run_req (r_sub12_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub03
		sub03_inst(
			.i_fld_T_0_addr_0 (w_sub03_T_addr),
			.i_fld_T_0_datain_0 (w_sub03_T_datain),
			.o_fld_T_0_dataout_0 (w_sub03_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub03_T_r_w),
			.i_fld_U_2_addr_0 (w_sub03_U_addr),
			.i_fld_U_2_datain_0 (w_sub03_U_datain),
			.o_fld_U_2_dataout_0 (w_sub03_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub03_U_r_w),
			.i_fld_V_1_addr_0 (w_sub03_V_addr),
			.i_fld_V_1_datain_0 (w_sub03_V_datain),
			.o_fld_V_1_dataout_0 (w_sub03_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub03_V_r_w),
			.i_fld_result_3_addr_0 (w_sub03_result_addr),
			.i_fld_result_3_datain_0 (w_sub03_result_datain),
			.o_fld_result_3_dataout_0 (w_sub03_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub03_result_r_w),
			.o_run_busy (w_sub03_run_busy),
			.i_run_req (r_sub03_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub02
		sub02_inst(
			.i_fld_T_0_addr_0 (w_sub02_T_addr),
			.i_fld_T_0_datain_0 (w_sub02_T_datain),
			.o_fld_T_0_dataout_0 (w_sub02_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub02_T_r_w),
			.i_fld_U_2_addr_0 (w_sub02_U_addr),
			.i_fld_U_2_datain_0 (w_sub02_U_datain),
			.o_fld_U_2_dataout_0 (w_sub02_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub02_U_r_w),
			.i_fld_V_1_addr_0 (w_sub02_V_addr),
			.i_fld_V_1_datain_0 (w_sub02_V_datain),
			.o_fld_V_1_dataout_0 (w_sub02_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub02_V_r_w),
			.i_fld_result_3_addr_0 (w_sub02_result_addr),
			.i_fld_result_3_datain_0 (w_sub02_result_datain),
			.o_fld_result_3_dataout_0 (w_sub02_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub02_result_r_w),
			.o_run_busy (w_sub02_run_busy),
			.i_run_req (r_sub02_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub11
		sub11_inst(
			.i_fld_T_0_addr_0 (w_sub11_T_addr),
			.i_fld_T_0_datain_0 (w_sub11_T_datain),
			.o_fld_T_0_dataout_0 (w_sub11_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub11_T_r_w),
			.i_fld_U_2_addr_0 (w_sub11_U_addr),
			.i_fld_U_2_datain_0 (w_sub11_U_datain),
			.o_fld_U_2_dataout_0 (w_sub11_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub11_U_r_w),
			.i_fld_V_1_addr_0 (w_sub11_V_addr),
			.i_fld_V_1_datain_0 (w_sub11_V_datain),
			.o_fld_V_1_dataout_0 (w_sub11_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub11_V_r_w),
			.i_fld_result_3_addr_0 (w_sub11_result_addr),
			.i_fld_result_3_datain_0 (w_sub11_result_datain),
			.o_fld_result_3_dataout_0 (w_sub11_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub11_result_r_w),
			.o_run_busy (w_sub11_run_busy),
			.i_run_req (r_sub11_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub14
		sub14_inst(
			.i_fld_T_0_addr_0 (w_sub14_T_addr),
			.i_fld_T_0_datain_0 (w_sub14_T_datain),
			.o_fld_T_0_dataout_0 (w_sub14_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub14_T_r_w),
			.i_fld_U_2_addr_0 (w_sub14_U_addr),
			.i_fld_U_2_datain_0 (w_sub14_U_datain),
			.o_fld_U_2_dataout_0 (w_sub14_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub14_U_r_w),
			.i_fld_V_1_addr_0 (w_sub14_V_addr),
			.i_fld_V_1_datain_0 (w_sub14_V_datain),
			.o_fld_V_1_dataout_0 (w_sub14_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub14_V_r_w),
			.i_fld_result_3_addr_0 (w_sub14_result_addr),
			.i_fld_result_3_datain_0 (w_sub14_result_datain),
			.o_fld_result_3_dataout_0 (w_sub14_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub14_result_r_w),
			.o_run_busy (w_sub14_run_busy),
			.i_run_req (r_sub14_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub01
		sub01_inst(
			.i_fld_T_0_addr_0 (w_sub01_T_addr),
			.i_fld_T_0_datain_0 (w_sub01_T_datain),
			.o_fld_T_0_dataout_0 (w_sub01_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub01_T_r_w),
			.i_fld_U_2_addr_0 (w_sub01_U_addr),
			.i_fld_U_2_datain_0 (w_sub01_U_datain),
			.o_fld_U_2_dataout_0 (w_sub01_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub01_U_r_w),
			.i_fld_V_1_addr_0 (w_sub01_V_addr),
			.i_fld_V_1_datain_0 (w_sub01_V_datain),
			.o_fld_V_1_dataout_0 (w_sub01_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub01_V_r_w),
			.i_fld_result_3_addr_0 (w_sub01_result_addr),
			.i_fld_result_3_datain_0 (w_sub01_result_datain),
			.o_fld_result_3_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub01_result_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub00
		sub00_inst(
			.i_fld_T_0_addr_0 (w_sub00_T_addr),
			.i_fld_T_0_datain_0 (w_sub00_T_datain),
			.o_fld_T_0_dataout_0 (w_sub00_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub00_T_r_w),
			.i_fld_U_2_addr_0 (w_sub00_U_addr),
			.i_fld_U_2_datain_0 (w_sub00_U_datain),
			.o_fld_U_2_dataout_0 (w_sub00_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub00_U_r_w),
			.i_fld_V_1_addr_0 (w_sub00_V_addr),
			.i_fld_V_1_datain_0 (w_sub00_V_datain),
			.o_fld_V_1_dataout_0 (w_sub00_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub00_V_r_w),
			.i_fld_result_3_addr_0 (w_sub00_result_addr),
			.i_fld_result_3_datain_0 (w_sub00_result_datain),
			.o_fld_result_3_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub00_result_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub13
		sub13_inst(
			.i_fld_T_0_addr_0 (w_sub13_T_addr),
			.i_fld_T_0_datain_0 (w_sub13_T_datain),
			.o_fld_T_0_dataout_0 (w_sub13_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub13_T_r_w),
			.i_fld_U_2_addr_0 (w_sub13_U_addr),
			.i_fld_U_2_datain_0 (w_sub13_U_datain),
			.o_fld_U_2_dataout_0 (w_sub13_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub13_U_r_w),
			.i_fld_V_1_addr_0 (w_sub13_V_addr),
			.i_fld_V_1_datain_0 (w_sub13_V_datain),
			.o_fld_V_1_dataout_0 (w_sub13_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub13_V_r_w),
			.i_fld_result_3_addr_0 (w_sub13_result_addr),
			.i_fld_result_3_datain_0 (w_sub13_result_datain),
			.o_fld_result_3_dataout_0 (w_sub13_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub13_result_r_w),
			.o_run_busy (w_sub13_run_busy),
			.i_run_req (r_sub13_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub07
		sub07_inst(
			.i_fld_T_0_addr_0 (w_sub07_T_addr),
			.i_fld_T_0_datain_0 (w_sub07_T_datain),
			.o_fld_T_0_dataout_0 (w_sub07_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub07_T_r_w),
			.i_fld_U_2_addr_0 (w_sub07_U_addr),
			.i_fld_U_2_datain_0 (w_sub07_U_datain),
			.o_fld_U_2_dataout_0 (w_sub07_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub07_U_r_w),
			.i_fld_V_1_addr_0 (w_sub07_V_addr),
			.i_fld_V_1_datain_0 (w_sub07_V_datain),
			.o_fld_V_1_dataout_0 (w_sub07_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub07_V_r_w),
			.i_fld_result_3_addr_0 (w_sub07_result_addr),
			.i_fld_result_3_datain_0 (w_sub07_result_datain),
			.o_fld_result_3_dataout_0 (w_sub07_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub07_result_r_w),
			.o_run_busy (w_sub07_run_busy),
			.i_run_req (r_sub07_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub16
		sub16_inst(
			.i_fld_T_0_addr_0 (w_sub16_T_addr),
			.i_fld_T_0_datain_0 (w_sub16_T_datain),
			.o_fld_T_0_dataout_0 (w_sub16_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub16_T_r_w),
			.i_fld_U_2_addr_0 (w_sub16_U_addr),
			.i_fld_U_2_datain_0 (w_sub16_U_datain),
			.o_fld_U_2_dataout_0 (w_sub16_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub16_U_r_w),
			.i_fld_V_1_addr_0 (w_sub16_V_addr),
			.i_fld_V_1_datain_0 (w_sub16_V_datain),
			.o_fld_V_1_dataout_0 (w_sub16_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub16_V_r_w),
			.i_fld_result_3_addr_0 (w_sub16_result_addr),
			.i_fld_result_3_datain_0 (w_sub16_result_datain),
			.o_fld_result_3_dataout_0 (w_sub16_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub16_result_r_w),
			.o_run_busy (w_sub16_run_busy),
			.i_run_req (r_sub16_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub06
		sub06_inst(
			.i_fld_T_0_addr_0 (w_sub06_T_addr),
			.i_fld_T_0_datain_0 (w_sub06_T_datain),
			.o_fld_T_0_dataout_0 (w_sub06_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub06_T_r_w),
			.i_fld_U_2_addr_0 (w_sub06_U_addr),
			.i_fld_U_2_datain_0 (w_sub06_U_datain),
			.o_fld_U_2_dataout_0 (w_sub06_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub06_U_r_w),
			.i_fld_V_1_addr_0 (w_sub06_V_addr),
			.i_fld_V_1_datain_0 (w_sub06_V_datain),
			.o_fld_V_1_dataout_0 (w_sub06_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub06_V_r_w),
			.i_fld_result_3_addr_0 (w_sub06_result_addr),
			.i_fld_result_3_datain_0 (w_sub06_result_datain),
			.o_fld_result_3_dataout_0 (w_sub06_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub06_result_r_w),
			.o_run_busy (w_sub06_run_busy),
			.i_run_req (r_sub06_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub15
		sub15_inst(
			.i_fld_T_0_addr_0 (w_sub15_T_addr),
			.i_fld_T_0_datain_0 (w_sub15_T_datain),
			.o_fld_T_0_dataout_0 (w_sub15_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub15_T_r_w),
			.i_fld_U_2_addr_0 (w_sub15_U_addr),
			.i_fld_U_2_datain_0 (w_sub15_U_datain),
			.o_fld_U_2_dataout_0 (w_sub15_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub15_U_r_w),
			.i_fld_V_1_addr_0 (w_sub15_V_addr),
			.i_fld_V_1_datain_0 (w_sub15_V_datain),
			.o_fld_V_1_dataout_0 (w_sub15_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub15_V_r_w),
			.i_fld_result_3_addr_0 (w_sub15_result_addr),
			.i_fld_result_3_datain_0 (w_sub15_result_datain),
			.o_fld_result_3_dataout_0 (w_sub15_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub15_result_r_w),
			.o_run_busy (w_sub15_run_busy),
			.i_run_req (r_sub15_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub05
		sub05_inst(
			.i_fld_T_0_addr_0 (w_sub05_T_addr),
			.i_fld_T_0_datain_0 (w_sub05_T_datain),
			.o_fld_T_0_dataout_0 (w_sub05_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub05_T_r_w),
			.i_fld_U_2_addr_0 (w_sub05_U_addr),
			.i_fld_U_2_datain_0 (w_sub05_U_datain),
			.o_fld_U_2_dataout_0 (w_sub05_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub05_U_r_w),
			.i_fld_V_1_addr_0 (w_sub05_V_addr),
			.i_fld_V_1_datain_0 (w_sub05_V_datain),
			.o_fld_V_1_dataout_0 (w_sub05_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub05_V_r_w),
			.i_fld_result_3_addr_0 (w_sub05_result_addr),
			.i_fld_result_3_datain_0 (w_sub05_result_datain),
			.o_fld_result_3_dataout_0 (w_sub05_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub05_result_r_w),
			.o_run_busy (w_sub05_run_busy),
			.i_run_req (r_sub05_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub18
		sub18_inst(
			.i_fld_T_0_addr_0 (w_sub18_T_addr),
			.i_fld_T_0_datain_0 (w_sub18_T_datain),
			.o_fld_T_0_dataout_0 (w_sub18_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub18_T_r_w),
			.i_fld_U_2_addr_0 (w_sub18_U_addr),
			.i_fld_U_2_datain_0 (w_sub18_U_datain),
			.o_fld_U_2_dataout_0 (w_sub18_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub18_U_r_w),
			.i_fld_V_1_addr_0 (w_sub18_V_addr),
			.i_fld_V_1_datain_0 (w_sub18_V_datain),
			.o_fld_V_1_dataout_0 (w_sub18_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub18_V_r_w),
			.i_fld_result_3_addr_0 (w_sub18_result_addr),
			.i_fld_result_3_datain_0 (w_sub18_result_datain),
			.o_fld_result_3_dataout_0 (w_sub18_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub18_result_r_w),
			.o_run_busy (w_sub18_run_busy),
			.i_run_req (r_sub18_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub04
		sub04_inst(
			.i_fld_T_0_addr_0 (w_sub04_T_addr),
			.i_fld_T_0_datain_0 (w_sub04_T_datain),
			.o_fld_T_0_dataout_0 (w_sub04_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub04_T_r_w),
			.i_fld_U_2_addr_0 (w_sub04_U_addr),
			.i_fld_U_2_datain_0 (w_sub04_U_datain),
			.o_fld_U_2_dataout_0 (w_sub04_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub04_U_r_w),
			.i_fld_V_1_addr_0 (w_sub04_V_addr),
			.i_fld_V_1_datain_0 (w_sub04_V_datain),
			.o_fld_V_1_dataout_0 (w_sub04_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub04_V_r_w),
			.i_fld_result_3_addr_0 (w_sub04_result_addr),
			.i_fld_result_3_datain_0 (w_sub04_result_datain),
			.o_fld_result_3_dataout_0 (w_sub04_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub04_result_r_w),
			.o_run_busy (w_sub04_run_busy),
			.i_run_req (r_sub04_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub17
		sub17_inst(
			.i_fld_T_0_addr_0 (w_sub17_T_addr),
			.i_fld_T_0_datain_0 (w_sub17_T_datain),
			.o_fld_T_0_dataout_0 (w_sub17_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub17_T_r_w),
			.i_fld_U_2_addr_0 (w_sub17_U_addr),
			.i_fld_U_2_datain_0 (w_sub17_U_datain),
			.o_fld_U_2_dataout_0 (w_sub17_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub17_U_r_w),
			.i_fld_V_1_addr_0 (w_sub17_V_addr),
			.i_fld_V_1_datain_0 (w_sub17_V_datain),
			.o_fld_V_1_dataout_0 (w_sub17_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub17_V_r_w),
			.i_fld_result_3_addr_0 (w_sub17_result_addr),
			.i_fld_result_3_datain_0 (w_sub17_result_datain),
			.o_fld_result_3_dataout_0 (w_sub17_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub17_result_r_w),
			.o_run_busy (w_sub17_run_busy),
			.i_run_req (r_sub17_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub10
		sub10_inst(
			.i_fld_T_0_addr_0 (w_sub10_T_addr),
			.i_fld_T_0_datain_0 (w_sub10_T_datain),
			.o_fld_T_0_dataout_0 (w_sub10_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub10_T_r_w),
			.i_fld_U_2_addr_0 (w_sub10_U_addr),
			.i_fld_U_2_datain_0 (w_sub10_U_datain),
			.o_fld_U_2_dataout_0 (w_sub10_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub10_U_r_w),
			.i_fld_V_1_addr_0 (w_sub10_V_addr),
			.i_fld_V_1_datain_0 (w_sub10_V_datain),
			.o_fld_V_1_dataout_0 (w_sub10_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub10_V_r_w),
			.i_fld_result_3_addr_0 (w_sub10_result_addr),
			.i_fld_result_3_datain_0 (w_sub10_result_datain),
			.o_fld_result_3_dataout_0 (w_sub10_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub10_result_r_w),
			.o_run_busy (w_sub10_run_busy),
			.i_run_req (r_sub10_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub20
		sub20_inst(
			.i_fld_T_0_addr_0 (w_sub20_T_addr),
			.i_fld_T_0_datain_0 (w_sub20_T_datain),
			.o_fld_T_0_dataout_0 (w_sub20_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub20_T_r_w),
			.i_fld_U_2_addr_0 (w_sub20_U_addr),
			.i_fld_U_2_datain_0 (w_sub20_U_datain),
			.o_fld_U_2_dataout_0 (w_sub20_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub20_U_r_w),
			.i_fld_V_1_addr_0 (w_sub20_V_addr),
			.i_fld_V_1_datain_0 (w_sub20_V_datain),
			.o_fld_V_1_dataout_0 (w_sub20_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub20_V_r_w),
			.i_fld_result_3_addr_0 (w_sub20_result_addr),
			.i_fld_result_3_datain_0 (w_sub20_result_datain),
			.o_fld_result_3_dataout_0 (w_sub20_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub20_result_r_w),
			.o_run_busy (w_sub20_run_busy),
			.i_run_req (r_sub20_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub21
		sub21_inst(
			.i_fld_T_0_addr_0 (w_sub21_T_addr),
			.i_fld_T_0_datain_0 (w_sub21_T_datain),
			.o_fld_T_0_dataout_0 (w_sub21_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub21_T_r_w),
			.i_fld_U_2_addr_0 (w_sub21_U_addr),
			.i_fld_U_2_datain_0 (w_sub21_U_datain),
			.o_fld_U_2_dataout_0 (w_sub21_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub21_U_r_w),
			.i_fld_V_1_addr_0 (w_sub21_V_addr),
			.i_fld_V_1_datain_0 (w_sub21_V_datain),
			.o_fld_V_1_dataout_0 (w_sub21_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub21_V_r_w),
			.i_fld_result_3_addr_0 (w_sub21_result_addr),
			.i_fld_result_3_datain_0 (w_sub21_result_datain),
			.o_fld_result_3_dataout_0 (w_sub21_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub21_result_r_w),
			.o_run_busy (w_sub21_run_busy),
			.i_run_req (r_sub21_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(10), .WORDS(1024) )
		dpram_T_0(
			.clk (clock),
			.ce_0 (w_fld_T_0_ce_0),
			.addr_0 (w_fld_T_0_addr_0),
			.datain_0 (w_fld_T_0_datain_0),
			.dataout_0 (w_fld_T_0_dataout_0),
			.r_w_0 (w_fld_T_0_r_w_0),
			.ce_1 (w_fld_T_0_ce_1),
			.addr_1 (r_fld_T_0_addr_1),
			.datain_1 (r_fld_T_0_datain_1),
			.dataout_1 (w_fld_T_0_dataout_1),
			.r_w_1 (r_fld_T_0_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(10), .WORDS(1024) )
		dpram_TT_1(
			.clk (clock),
			.ce_0 (w_fld_TT_1_ce_0),
			.addr_0 (w_fld_TT_1_addr_0),
			.datain_0 (w_fld_TT_1_datain_0),
			.dataout_0 (w_fld_TT_1_dataout_0),
			.r_w_0 (w_fld_TT_1_r_w_0),
			.ce_1 (w_fld_TT_1_ce_1),
			.addr_1 (r_fld_TT_1_addr_1),
			.datain_1 (r_fld_TT_1_datain_1),
			.dataout_1 (w_fld_TT_1_dataout_1),
			.r_w_1 (r_fld_TT_1_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(10), .WORDS(1024) )
		dpram_U_2(
			.clk (clock),
			.ce_0 (w_fld_U_2_ce_0),
			.addr_0 (w_fld_U_2_addr_0),
			.datain_0 (w_fld_U_2_datain_0),
			.dataout_0 (w_fld_U_2_dataout_0),
			.r_w_0 (w_fld_U_2_r_w_0),
			.ce_1 (w_fld_U_2_ce_1),
			.addr_1 (r_fld_U_2_addr_1),
			.datain_1 (r_fld_U_2_datain_1),
			.dataout_1 (w_fld_U_2_dataout_1),
			.r_w_1 (r_fld_U_2_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(10), .WORDS(1024) )
		dpram_V_3(
			.clk (clock),
			.ce_0 (w_fld_V_3_ce_0),
			.addr_0 (w_fld_V_3_addr_0),
			.datain_0 (w_fld_V_3_datain_0),
			.dataout_0 (w_fld_V_3_dataout_0),
			.r_w_0 (w_fld_V_3_r_w_0),
			.ce_1 (w_fld_V_3_ce_1),
			.addr_1 (r_fld_V_3_addr_1),
			.datain_1 (r_fld_V_3_datain_1),
			.dataout_1 (w_fld_V_3_dataout_1),
			.r_w_1 (r_fld_V_3_r_w_1)
		);

	DivInt
		DivInt_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.dividend (r_ip_DivInt_dividend_0),
			.divisor (r_ip_DivInt_divisor_0),
			.fractional (w_ip_DivInt_fractional_0),
			.quotient (w_ip_DivInt_quotient_0)
		);

	DivInt
		DivInt_inst_1(
			.clk (clock),
			.ce (w_sys_ce),
			.dividend (r_ip_DivInt_dividend_1),
			.divisor (r_ip_DivInt_divisor_1),
			.fractional (w_ip_DivInt_fractional_1),
			.quotient (w_ip_DivInt_quotient_1)
		);

	AddFloat
		AddFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_AddFloat_portA_0),
			.b (r_ip_AddFloat_portB_0),
			.result (w_ip_AddFloat_result_0)
		);

	MultFloat
		MultFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_MultFloat_multiplicand_0),
			.b (r_ip_MultFloat_multiplier_0),
			.result (w_ip_MultFloat_product_0)
		);

	FixedToFloat
		FixedToFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_FixedToFloat_fixed_0),
			.result (w_ip_FixedToFloat_floating_0)
		);

	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_ip_DivInt_dividend_0 <= r_run_mx_32;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_ip_DivInt_divisor_0 <= w_sys_tmp2686;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_ip_DivInt_dividend_1 <= r_run_mx_32;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_ip_DivInt_divisor_1 <= w_sys_tmp2690;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'hc) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h14)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp39;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'hc)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp38[31], w_sys_tmp38[30:0] };

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp38[31], w_sys_tmp38[30:0] };

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp129[31], w_sys_tmp129[30:0] };

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp129[31], w_sys_tmp129[30:0] };

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp38[31], w_sys_tmp38[30:0] };

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp38[31], w_sys_tmp38[30:0] };

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp38[31], w_sys_tmp38[30:0] };

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'hc) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h16)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp37;

									end
									else
									if((8'h7<=r_sys_run_step && r_sys_run_step<=8'hb) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'hf)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_dy_36;

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==8'h13) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1a)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp19;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h19)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==8'h13) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h1a)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==8'hd) || (r_sys_run_step==8'hf)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp38;

									end
									else
									if((r_sys_run_step==8'he) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h16)) begin
										r_ip_MultFloat_multiplier_0 <= r_run_YY_41;

									end
									else
									if((r_sys_run_step==8'h15) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1b)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp2_float;

									end
									else
									if((8'h7<=r_sys_run_step && r_sys_run_step<=8'hb)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp20;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_ip_FixedToFloat_fixed_0 <= w_sys_tmp21;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						7'h4d: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 7'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h0: begin
							r_sys_run_phase <= 7'h2;
						end

						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'h4;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'h5;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp13) ? 7'h9 : 7'hf);

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'h5;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'ha;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp16) ? 7'hd : 7'h6);

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h20)) begin
										r_sys_run_phase <= 7'ha;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'h10;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp227) ? 7'h13 : 7'h15);

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h9d)) begin
										r_sys_run_phase <= 7'h10;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'h16;

									end
								end

							endcase
						end

						7'h16: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2105) ? 7'h19 : 7'h1b);

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h28)) begin
										r_sys_run_phase <= 7'h16;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'h1c;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2578) ? 7'h20 : 7'h4d);

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'h1c;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'h21;

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2581) ? 7'h24 : 7'h26);

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_run_phase <= 7'h21;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'h27;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2598) ? 7'h2a : 7'h2c);

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'hd)) begin
										r_sys_run_phase <= 7'h27;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'h2d;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h25)) begin
										r_sys_run_phase <= ((w_sys_tmp2687) ? 7'h30 : 7'h32);

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_run_phase <= 7'h2d;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'h33;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2734) ? 7'h36 : 7'h38);

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h9d)) begin
										r_sys_run_phase <= 7'h33;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'h39;

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3676) ? 7'h3c : 7'h3d);

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h28)) begin
										r_sys_run_phase <= 7'h39;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h18: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_phase <= 7'h3f;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h18: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_phase <= 7'h41;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'h42;

									end
								end

							endcase
						end

						7'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3916) ? 7'h45 : 7'h47);

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h75)) begin
										r_sys_run_phase <= 7'h42;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'h48;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4508) ? 7'h4b : 7'h1d);

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1e)) begin
										r_sys_run_phase <= 7'h48;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sys_run_phase <= 7'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 5'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h20)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h9d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h16: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h28)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'hd)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h25)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h25)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h9d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h28)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h75)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1e)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 8'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h20)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h1f)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h9c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==8'h9d)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h16: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h28)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h27)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h1) || (r_sys_run_step==8'h2)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'hd)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'hc)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h25)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h24)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h25)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h24)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h9d)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h9c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h28)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h27)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub00_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub01_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub02_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub03_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub04_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub05_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub06_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub07_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub08_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub09_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub10_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub11_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub12_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub13_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub14_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub15_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub16_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub17_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub18_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub19_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub20_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub21_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub22_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub23_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub24_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h75)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h74)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1e)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h1d)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						7'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						7'h4d: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_T_0_addr_1 <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp23[9:0] );

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2593[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2589[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2585[9:0] );

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1) || (r_sys_run_step==8'h3) || (r_sys_run_step==8'h5) || (r_sys_run_step==8'h7) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'hd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2607[9:0] );

									end
									else
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h2) || (r_sys_run_step==8'h4) || (r_sys_run_step==8'h6) || (r_sys_run_step==8'h8) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'hc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2602[9:0] );

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2693[9:0] );

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h32)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3039[9:0] );

									end
									else
									if((r_sys_run_step==8'h29)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2985[9:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2865[9:0] );

									end
									else
									if((r_sys_run_step==8'h5d) || (r_sys_run_step==8'h5f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3297[9:0] );

									end
									else
									if((r_sys_run_step==8'h49)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3177[9:0] );

									end
									else
									if((r_sys_run_step==8'h64) || (r_sys_run_step==8'h66)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3339[9:0] );

									end
									else
									if((r_sys_run_step==8'h53)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3237[9:0] );

									end
									else
									if((r_sys_run_step==8'h89)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3561[9:0] );

									end
									else
									if((r_sys_run_step==8'h3d) || (r_sys_run_step==8'h3f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3105[9:0] );

									end
									else
									if((r_sys_run_step==8'h94) || (r_sys_run_step==8'h96)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3627[9:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2811[9:0] );

									end
									else
									if((r_sys_run_step==8'h4b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3189[9:0] );

									end
									else
									if((r_sys_run_step==8'h4a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3183[9:0] );

									end
									else
									if((r_sys_run_step==8'h98)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3651[9:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2847[9:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2943[9:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2907[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2769[9:0] );

									end
									else
									if((r_sys_run_step==8'h2c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3003[9:0] );

									end
									else
									if((r_sys_run_step==8'h83) || (r_sys_run_step==8'h85)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3525[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2739[9:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2799[9:0] );

									end
									else
									if((r_sys_run_step==8'h2e) || (r_sys_run_step==8'h30)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3015[9:0] );

									end
									else
									if((r_sys_run_step==8'h4e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3207[9:0] );

									end
									else
									if((r_sys_run_step==8'h59)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3273[9:0] );

									end
									else
									if((r_sys_run_step==8'h65) || (r_sys_run_step==8'h67)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3345[9:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2961[9:0] );

									end
									else
									if((r_sys_run_step==8'h7b) || (r_sys_run_step==8'h7d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3477[9:0] );

									end
									else
									if((r_sys_run_step==8'h16) || (r_sys_run_step==8'h18)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2871[9:0] );

									end
									else
									if((r_sys_run_step==8'h1f) || (r_sys_run_step==8'h21)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2925[9:0] );

									end
									else
									if((r_sys_run_step==8'h58)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3267[9:0] );

									end
									else
									if((r_sys_run_step==8'h63)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3333[9:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2853[9:0] );

									end
									else
									if((r_sys_run_step==8'h81)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3513[9:0] );

									end
									else
									if((r_sys_run_step==8'h75)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3441[9:0] );

									end
									else
									if((r_sys_run_step==8'h88)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3555[9:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2805[9:0] );

									end
									else
									if((r_sys_run_step==8'h69)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3369[9:0] );

									end
									else
									if((r_sys_run_step==8'h8f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3597[9:0] );

									end
									else
									if((r_sys_run_step==8'h31)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3033[9:0] );

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3363[9:0] );

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2955[9:0] );

									end
									else
									if((r_sys_run_step==8'h8a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3567[9:0] );

									end
									else
									if((r_sys_run_step==8'h74)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3435[9:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2859[9:0] );

									end
									else
									if((r_sys_run_step==8'h3a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3087[9:0] );

									end
									else
									if((r_sys_run_step==8'h43)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3141[9:0] );

									end
									else
									if((r_sys_run_step==8'h50)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3219[9:0] );

									end
									else
									if((r_sys_run_step==8'h87)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3549[9:0] );

									end
									else
									if((r_sys_run_step==8'h6d) || (r_sys_run_step==8'h6f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3393[9:0] );

									end
									else
									if((r_sys_run_step==8'h9a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3663[9:0] );

									end
									else
									if((r_sys_run_step==8'h82)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3519[9:0] );

									end
									else
									if((r_sys_run_step==8'hf) || (r_sys_run_step==8'h11)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2829[9:0] );

									end
									else
									if((r_sys_run_step==8'h55) || (r_sys_run_step==8'h57)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3249[9:0] );

									end
									else
									if((r_sys_run_step==8'h5a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3279[9:0] );

									end
									else
									if((r_sys_run_step==8'h84) || (r_sys_run_step==8'h86)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3531[9:0] );

									end
									else
									if((r_sys_run_step==8'he) || (r_sys_run_step==8'h10)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2823[9:0] );

									end
									else
									if((r_sys_run_step==8'h41)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3129[9:0] );

									end
									else
									if((r_sys_run_step==8'h6) || (r_sys_run_step==8'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2775[9:0] );

									end
									else
									if((r_sys_run_step==8'h72)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3423[9:0] );

									end
									else
									if((r_sys_run_step==8'h35) || (r_sys_run_step==8'h37)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3057[9:0] );

									end
									else
									if((r_sys_run_step==8'h4c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3195[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2745[9:0] );

									end
									else
									if((r_sys_run_step==8'h3b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3093[9:0] );

									end
									else
									if((r_sys_run_step==8'h3e) || (r_sys_run_step==8'h40)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3111[9:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2967[9:0] );

									end
									else
									if((r_sys_run_step==8'h62)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3327[9:0] );

									end
									else
									if((r_sys_run_step==8'h73)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3429[9:0] );

									end
									else
									if((r_sys_run_step==8'h45) || (r_sys_run_step==8'h47)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3153[9:0] );

									end
									else
									if((r_sys_run_step==8'h4d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3201[9:0] );

									end
									else
									if((r_sys_run_step==8'h54) || (r_sys_run_step==8'h56)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3243[9:0] );

									end
									else
									if((r_sys_run_step==8'h91)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3609[9:0] );

									end
									else
									if((r_sys_run_step==8'h8c) || (r_sys_run_step==8'h8e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3579[9:0] );

									end
									else
									if((r_sys_run_step==8'h71)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3417[9:0] );

									end
									else
									if((r_sys_run_step==8'h9b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3669[9:0] );

									end
									else
									if((r_sys_run_step==8'h79)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3465[9:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2949[9:0] );

									end
									else
									if((r_sys_run_step==8'h7c) || (r_sys_run_step==8'h7e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3483[9:0] );

									end
									else
									if((r_sys_run_step==8'h36) || (r_sys_run_step==8'h38)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3063[9:0] );

									end
									else
									if((r_sys_run_step==8'h2b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2997[9:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2901[9:0] );

									end
									else
									if((r_sys_run_step==8'h92)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3615[9:0] );

									end
									else
									if((r_sys_run_step==8'h42)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3135[9:0] );

									end
									else
									if((r_sys_run_step==8'h7f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3501[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2763[9:0] );

									end
									else
									if((r_sys_run_step==8'h52)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3231[9:0] );

									end
									else
									if((r_sys_run_step==8'h6a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3375[9:0] );

									end
									else
									if((r_sys_run_step==8'h61)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3321[9:0] );

									end
									else
									if((r_sys_run_step==8'h7a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3471[9:0] );

									end
									else
									if((r_sys_run_step==8'h5b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3285[9:0] );

									end
									else
									if((r_sys_run_step==8'h97)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3645[9:0] );

									end
									else
									if((r_sys_run_step==8'h1e) || (r_sys_run_step==8'h20)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2919[9:0] );

									end
									else
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'h9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2781[9:0] );

									end
									else
									if((r_sys_run_step==8'h80)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3507[9:0] );

									end
									else
									if((r_sys_run_step==8'h51)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3225[9:0] );

									end
									else
									if((r_sys_run_step==8'h5c) || (r_sys_run_step==8'h5e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3291[9:0] );

									end
									else
									if((r_sys_run_step==8'h93) || (r_sys_run_step==8'h95)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3621[9:0] );

									end
									else
									if((r_sys_run_step==8'h76)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3447[9:0] );

									end
									else
									if((r_sys_run_step==8'h4f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3213[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2757[9:0] );

									end
									else
									if((r_sys_run_step==8'h6c) || (r_sys_run_step==8'h6e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3387[9:0] );

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2979[9:0] );

									end
									else
									if((r_sys_run_step==8'h60)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3315[9:0] );

									end
									else
									if((r_sys_run_step==8'h77)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3453[9:0] );

									end
									else
									if((r_sys_run_step==8'h17) || (r_sys_run_step==8'h19)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2877[9:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2817[9:0] );

									end
									else
									if((r_sys_run_step==8'h8b) || (r_sys_run_step==8'h8d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3573[9:0] );

									end
									else
									if((r_sys_run_step==8'h2d) || (r_sys_run_step==8'h2f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3009[9:0] );

									end
									else
									if((r_sys_run_step==8'h33)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3045[9:0] );

									end
									else
									if((r_sys_run_step==8'h3c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3099[9:0] );

									end
									else
									if((r_sys_run_step==8'h70)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3411[9:0] );

									end
									else
									if((r_sys_run_step==8'h39)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3081[9:0] );

									end
									else
									if((r_sys_run_step==8'h46) || (r_sys_run_step==8'h48)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3159[9:0] );

									end
									else
									if((r_sys_run_step==8'h2a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2991[9:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2913[9:0] );

									end
									else
									if((r_sys_run_step==8'h99)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3657[9:0] );

									end
									else
									if((r_sys_run_step==8'h90)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3603[9:0] );

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2973[9:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2895[9:0] );

									end
									else
									if((r_sys_run_step==8'h44)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3147[9:0] );

									end
									else
									if((r_sys_run_step==8'h34)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3051[9:0] );

									end
									else
									if((r_sys_run_step==8'h78)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3459[9:0] );

									end
									else
									if((r_sys_run_step==8'h6b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3381[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2751[9:0] );

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h25)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3903[9:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3789[9:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3759[9:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3801[9:0] );

									end
									else
									if((r_sys_run_step==8'h1f) || (r_sys_run_step==8'h21)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3867[9:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3795[9:0] );

									end
									else
									if((r_sys_run_step==8'h6) || (r_sys_run_step==8'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3717[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3687[9:0] );

									end
									else
									if((r_sys_run_step==8'h17) || (r_sys_run_step==8'h19)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3819[9:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3849[9:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3885[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3711[9:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3891[9:0] );

									end
									else
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'h9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3723[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3693[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3681[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3699[9:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3741[9:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3843[9:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3753[9:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3747[9:0] );

									end
									else
									if((r_sys_run_step==8'h16) || (r_sys_run_step==8'h18)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3813[9:0] );

									end
									else
									if((r_sys_run_step==8'h1e) || (r_sys_run_step==8'h20)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3861[9:0] );

									end
									else
									if((r_sys_run_step==8'hf) || (r_sys_run_step==8'h11)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3771[9:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3909[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3705[9:0] );

									end
									else
									if((r_sys_run_step==8'he) || (r_sys_run_step==8'h10)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3765[9:0] );

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3897[9:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3807[9:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3855[9:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3837[9:0] );

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4377[9:0] );

									end
									else
									if((r_sys_run_step==8'h2f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4152[9:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4047[9:0] );

									end
									else
									if((r_sys_run_step==8'h4f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4312[9:0] );

									end
									else
									if((r_sys_run_step==8'h3d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4222[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3921[9:0] );

									end
									else
									if((r_sys_run_step==8'h50)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4317[9:0] );

									end
									else
									if((r_sys_run_step==8'h58)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4357[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3933[9:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3992[9:0] );

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4037[9:0] );

									end
									else
									if((r_sys_run_step==8'h62)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4407[9:0] );

									end
									else
									if((r_sys_run_step==8'h6a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4447[9:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3951[9:0] );

									end
									else
									if((r_sys_run_step==8'h31)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4162[9:0] );

									end
									else
									if((r_sys_run_step==8'h40)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4237[9:0] );

									end
									else
									if((r_sys_run_step==8'h4e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4307[9:0] );

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3987[9:0] );

									end
									else
									if((r_sys_run_step==8'h3a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4207[9:0] );

									end
									else
									if((r_sys_run_step==8'h49)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4282[9:0] );

									end
									else
									if((r_sys_run_step==8'h1f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4072[9:0] );

									end
									else
									if((r_sys_run_step==8'h3c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4217[9:0] );

									end
									else
									if((r_sys_run_step==8'h42)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4247[9:0] );

									end
									else
									if((r_sys_run_step==8'h65)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4422[9:0] );

									end
									else
									if((r_sys_run_step==8'h54)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4337[9:0] );

									end
									else
									if((r_sys_run_step==8'h61)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4402[9:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3962[9:0] );

									end
									else
									if((r_sys_run_step==8'h3e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4227[9:0] );

									end
									else
									if((r_sys_run_step==8'h6e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4467[9:0] );

									end
									else
									if((r_sys_run_step==8'h30)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4157[9:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4102[9:0] );

									end
									else
									if((r_sys_run_step==8'h53)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4332[9:0] );

									end
									else
									if((r_sys_run_step==8'h64)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4417[9:0] );

									end
									else
									if((r_sys_run_step==8'h5e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4387[9:0] );

									end
									else
									if((r_sys_run_step==8'h29)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4122[9:0] );

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4027[9:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3967[9:0] );

									end
									else
									if((r_sys_run_step==8'h48)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4277[9:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4002[9:0] );

									end
									else
									if((r_sys_run_step==8'h33)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4172[9:0] );

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4117[9:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4062[9:0] );

									end
									else
									if((r_sys_run_step==8'h60)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4397[9:0] );

									end
									else
									if((r_sys_run_step==8'h39)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4202[9:0] );

									end
									else
									if((r_sys_run_step==8'h45)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4262[9:0] );

									end
									else
									if((r_sys_run_step==8'h72)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4487[9:0] );

									end
									else
									if((r_sys_run_step==8'h2c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4137[9:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4057[9:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4052[9:0] );

									end
									else
									if((r_sys_run_step==8'h75)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4502[9:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3982[9:0] );

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4042[9:0] );

									end
									else
									if((r_sys_run_step==8'h35)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4182[9:0] );

									end
									else
									if((r_sys_run_step==8'h6d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4462[9:0] );

									end
									else
									if((r_sys_run_step==8'h2a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4127[9:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4012[9:0] );

									end
									else
									if((r_sys_run_step==8'h2e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4147[9:0] );

									end
									else
									if((r_sys_run_step==8'h47)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4272[9:0] );

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4437[9:0] );

									end
									else
									if((r_sys_run_step==8'h70)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4477[9:0] );

									end
									else
									if((r_sys_run_step==8'h74)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4497[9:0] );

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4097[9:0] );

									end
									else
									if((r_sys_run_step==8'h63)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4412[9:0] );

									end
									else
									if((r_sys_run_step==8'h36)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4187[9:0] );

									end
									else
									if((r_sys_run_step==8'h5f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4392[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3927[9:0] );

									end
									else
									if((r_sys_run_step==8'h34)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4177[9:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4092[9:0] );

									end
									else
									if((r_sys_run_step==8'h69)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4442[9:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4022[9:0] );

									end
									else
									if((r_sys_run_step==8'h4d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4302[9:0] );

									end
									else
									if((r_sys_run_step==8'h38)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4197[9:0] );

									end
									else
									if((r_sys_run_step==8'h5a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4367[9:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4087[9:0] );

									end
									else
									if((r_sys_run_step==8'h44)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4257[9:0] );

									end
									else
									if((r_sys_run_step==8'h46)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4267[9:0] );

									end
									else
									if((r_sys_run_step==8'h41)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4242[9:0] );

									end
									else
									if((r_sys_run_step==8'h5d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4382[9:0] );

									end
									else
									if((r_sys_run_step==8'h4a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4287[9:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4017[9:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4032[9:0] );

									end
									else
									if((r_sys_run_step==8'h52)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4327[9:0] );

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4112[9:0] );

									end
									else
									if((r_sys_run_step==8'h73)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4492[9:0] );

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3957[9:0] );

									end
									else
									if((r_sys_run_step==8'h32)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4167[9:0] );

									end
									else
									if((r_sys_run_step==8'h56)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4347[9:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3977[9:0] );

									end
									else
									if((r_sys_run_step==8'h2b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4132[9:0] );

									end
									else
									if((r_sys_run_step==8'h6f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4472[9:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3972[9:0] );

									end
									else
									if((r_sys_run_step==8'h4b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4292[9:0] );

									end
									else
									if((r_sys_run_step==8'h20)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4077[9:0] );

									end
									else
									if((r_sys_run_step==8'h71)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4482[9:0] );

									end
									else
									if((r_sys_run_step==8'h37)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4192[9:0] );

									end
									else
									if((r_sys_run_step==8'h4c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4297[9:0] );

									end
									else
									if((r_sys_run_step==8'h67)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4432[9:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4007[9:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4107[9:0] );

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4067[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3939[9:0] );

									end
									else
									if((r_sys_run_step==8'h66)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4427[9:0] );

									end
									else
									if((r_sys_run_step==8'h6b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4452[9:0] );

									end
									else
									if((r_sys_run_step==8'h2d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4142[9:0] );

									end
									else
									if((r_sys_run_step==8'h6c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4457[9:0] );

									end
									else
									if((r_sys_run_step==8'h55)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4342[9:0] );

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3997[9:0] );

									end
									else
									if((r_sys_run_step==8'h3f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4232[9:0] );

									end
									else
									if((r_sys_run_step==8'h59)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4362[9:0] );

									end
									else
									if((r_sys_run_step==8'h21)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4082[9:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3945[9:0] );

									end
									else
									if((r_sys_run_step==8'h43)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4252[9:0] );

									end
									else
									if((r_sys_run_step==8'h51)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4322[9:0] );

									end
									else
									if((r_sys_run_step==8'h5b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4372[9:0] );

									end
									else
									if((r_sys_run_step==8'h57)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4352[9:0] );

									end
									else
									if((r_sys_run_step==8'h3b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4212[9:0] );

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'hb)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4564[9:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4614[9:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4584[9:0] );

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4549[9:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4554[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4531[9:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4639[9:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4649[9:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4624[9:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4644[9:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4537[9:0] );

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4589[9:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4594[9:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4604[9:0] );

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4619[9:0] );

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4659[9:0] );

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4629[9:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4569[9:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4654[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4525[9:0] );

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4579[9:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4559[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4519[9:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4543[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4513[9:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4574[9:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4609[9:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4599[9:0] );

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4634[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp26;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp2592;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp2587;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'hd)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp2605;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp2696;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h15)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp73_float;

									end
									else
									if((r_sys_run_step==8'h5f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp96_float;

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp70_float;

									end
									else
									if((r_sys_run_step==8'h5b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp60_float;

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp90_float;

									end
									else
									if((r_sys_run_step==8'h54)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp101_float;

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp53_float;

									end
									else
									if((r_sys_run_step==8'h30)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp109_float;

									end
									else
									if((r_sys_run_step==8'h5d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp30_float;

									end
									else
									if((r_sys_run_step==8'h59)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp100_float;

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==8'h65)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp99_float;

									end
									else
									if((r_sys_run_step==8'h2a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==8'h5a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp86_float;

									end
									else
									if((r_sys_run_step==8'h2b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp106_float;

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp52_float;

									end
									else
									if((r_sys_run_step==8'h5e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==8'h73)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp56_float;

									end
									else
									if((r_sys_run_step==8'h45)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp48_float;

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp18_float;

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp54_float;

									end
									else
									if((r_sys_run_step==8'h48)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp95_float;

									end
									else
									if((r_sys_run_step==8'h4d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==8'h39)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp55_float;

									end
									else
									if((r_sys_run_step==8'h50)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp62_float;

									end
									else
									if((r_sys_run_step==8'h6f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp27_float;

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp75_float;

									end
									else
									if((r_sys_run_step==8'h44)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp64_float;

									end
									else
									if((r_sys_run_step==8'h66)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp85_float;

									end
									else
									if((r_sys_run_step==8'h4a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp63_float;

									end
									else
									if((r_sys_run_step==8'h55)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp81_float;

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp107_float;

									end
									else
									if((r_sys_run_step==8'h32)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp89_float;

									end
									else
									if((r_sys_run_step==8'h1f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp93_float;

									end
									else
									if((r_sys_run_step==8'h53)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==8'h6e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp42_float;

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==8'h34)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp50_float;

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp72_float;

									end
									else
									if((r_sys_run_step==8'h4b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp47_float;

									end
									else
									if((r_sys_run_step==8'h29)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp33_float;

									end
									else
									if((r_sys_run_step==8'h52)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp24_float;

									end
									else
									if((r_sys_run_step==8'h38)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp78_float;

									end
									else
									if((r_sys_run_step==8'h62)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp45_float;

									end
									else
									if((r_sys_run_step==8'h4c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp31_float;

									end
									else
									if((r_sys_run_step==8'h61)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp59_float;

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp35_float;

									end
									else
									if((r_sys_run_step==8'h6d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp57_float;

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp91_float;

									end
									else
									if((r_sys_run_step==8'h43)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp79_float;

									end
									else
									if((r_sys_run_step==8'h49)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp87_float;

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp37_float;

									end
									else
									if((r_sys_run_step==8'h35)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp22_float;

									end
									else
									if((r_sys_run_step==8'h75)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp28_float;

									end
									else
									if((r_sys_run_step==8'h4f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp80_float;

									end
									else
									if((r_sys_run_step==8'h46)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp23_float;

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp92_float;

									end
									else
									if((r_sys_run_step==8'h74)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp43_float;

									end
									else
									if((r_sys_run_step==8'h4e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp102_float;

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp71_float;

									end
									else
									if((r_sys_run_step==8'h20)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp76_float;

									end
									else
									if((r_sys_run_step==8'h2f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp20_float;

									end
									else
									if((r_sys_run_step==8'h5c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp46_float;

									end
									else
									if((r_sys_run_step==8'h67)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp58_float;

									end
									else
									if((r_sys_run_step==8'h3d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp88_float;

									end
									else
									if((r_sys_run_step==8'h69)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp29_float;

									end
									else
									if((r_sys_run_step==8'h33)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp66_float;

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp74_float;

									end
									else
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h7)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp3923;

									end
									else
									if((r_sys_run_step==8'h2d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp67_float;

									end
									else
									if((r_sys_run_step==8'h71)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp97_float;

									end
									else
									if((r_sys_run_step==8'h42)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp103_float;

									end
									else
									if((r_sys_run_step==8'h58)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp25_float;

									end
									else
									if((r_sys_run_step==8'h6b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp98_float;

									end
									else
									if((r_sys_run_step==8'h57)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp40_float;

									end
									else
									if((r_sys_run_step==8'h63)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp26_float;

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp36_float;

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==8'h6c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp83_float;

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp19_float;

									end
									else
									if((r_sys_run_step==8'h3e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp65_float;

									end
									else
									if((r_sys_run_step==8'h70)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp14_float;

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp68_float;

									end
									else
									if((r_sys_run_step==8'h6a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp51_float;

									end
									else
									if((r_sys_run_step==8'h64)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==8'h3c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp104_float;

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp34_float;

									end
									else
									if((r_sys_run_step==8'h72)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp84_float;

									end
									else
									if((r_sys_run_step==8'h51)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp41_float;

									end
									else
									if((r_sys_run_step==8'h56)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp61_float;

									end
									else
									if((r_sys_run_step==8'h31)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp105_float;

									end
									else
									if((r_sys_run_step==8'h2c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp77_float;

									end
									else
									if((r_sys_run_step==8'h47)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==8'h3a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp49_float;

									end
									else
									if((r_sys_run_step==8'h3b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp21_float;

									end
									else
									if((r_sys_run_step==8'h40)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp32_float;

									end
									else
									if((r_sys_run_step==8'h36)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp44_float;

									end
									else
									if((r_sys_run_step==8'h37)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp94_float;

									end
									else
									if((r_sys_run_step==8'h3f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp39_float;

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp108_float;

									end
									else
									if((r_sys_run_step==8'h21)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp69_float;

									end
									else
									if((r_sys_run_step==8'h41)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==8'h2e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp38_float;

									end
									else
									if((r_sys_run_step==8'h60)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp82_float;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp23_float;

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp21_float;

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp18_float;

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp25_float;

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp24_float;

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp26_float;

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp19_float;

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp20_float;

									end
									else
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h7)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp4515;

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp14_float;

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp27_float;

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp22_float;

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp5_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_T_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h3)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'hd)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h9b)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h26)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h75)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h1e)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin
							r_fld_T_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_TT_1_addr_1 <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_fld_TT_1_addr_1 <= $signed( w_sys_tmp28[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_fld_TT_1_datain_1 <= w_sys_tmp26;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_TT_1_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_fld_TT_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin
							r_fld_TT_1_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_U_2_addr_1 <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h18) || (r_sys_run_step==8'h1a) || (8'h1c<=r_sys_run_step && r_sys_run_step<=8'h20)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp33[9:0] );

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h8c) || (r_sys_run_step==8'h8e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1912[9:0] );

									end
									else
									if((r_sys_run_step==8'h44)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1048[9:0] );

									end
									else
									if((r_sys_run_step==8'h76)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1648[9:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp472[9:0] );

									end
									else
									if((r_sys_run_step==8'h5b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1324[9:0] );

									end
									else
									if((r_sys_run_step==8'h2a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp736[9:0] );

									end
									else
									if((r_sys_run_step==8'h91)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1972[9:0] );

									end
									else
									if((r_sys_run_step==8'h81)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1780[9:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp544[9:0] );

									end
									else
									if((r_sys_run_step==8'h72)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1600[9:0] );

									end
									else
									if((r_sys_run_step==8'h7b) || (r_sys_run_step==8'h7d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1708[9:0] );

									end
									else
									if((r_sys_run_step==8'h35) || (r_sys_run_step==8'h37)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp868[9:0] );

									end
									else
									if((r_sys_run_step==8'h69)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1492[9:0] );

									end
									else
									if((r_sys_run_step==8'h61)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1396[9:0] );

									end
									else
									if((r_sys_run_step==8'h3e) || (r_sys_run_step==8'h40)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp976[9:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp448[9:0] );

									end
									else
									if((r_sys_run_step==8'he) || (r_sys_run_step==8'h10)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp400[9:0] );

									end
									else
									if((r_sys_run_step==8'h39)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp916[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp268[9:0] );

									end
									else
									if((r_sys_run_step==8'h8f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1948[9:0] );

									end
									else
									if((r_sys_run_step==8'h46) || (r_sys_run_step==8'h48)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1072[9:0] );

									end
									else
									if((r_sys_run_step==8'h71)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1588[9:0] );

									end
									else
									if((r_sys_run_step==8'h79)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1684[9:0] );

									end
									else
									if((r_sys_run_step==8'h2b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp748[9:0] );

									end
									else
									if((r_sys_run_step==8'h55) || (r_sys_run_step==8'h57)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1252[9:0] );

									end
									else
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'h9)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp316[9:0] );

									end
									else
									if((r_sys_run_step==8'h75)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1636[9:0] );

									end
									else
									if((r_sys_run_step==8'h16) || (r_sys_run_step==8'h18)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp496[9:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp352[9:0] );

									end
									else
									if((r_sys_run_step==8'h87)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1852[9:0] );

									end
									else
									if((r_sys_run_step==8'h88)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1864[9:0] );

									end
									else
									if((r_sys_run_step==8'h6) || (r_sys_run_step==8'h8)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp304[9:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp580[9:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp376[9:0] );

									end
									else
									if((r_sys_run_step==8'h6a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1504[9:0] );

									end
									else
									if((r_sys_run_step==8'h41)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1012[9:0] );

									end
									else
									if((r_sys_run_step==8'h50)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1192[9:0] );

									end
									else
									if((r_sys_run_step==8'h7c) || (r_sys_run_step==8'h7e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1720[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp232[9:0] );

									end
									else
									if((r_sys_run_step==8'h77)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1660[9:0] );

									end
									else
									if((r_sys_run_step==8'h45) || (r_sys_run_step==8'h47)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1060[9:0] );

									end
									else
									if((r_sys_run_step==8'h93) || (r_sys_run_step==8'h95)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1996[9:0] );

									end
									else
									if((r_sys_run_step==8'h84) || (r_sys_run_step==8'h86)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1816[9:0] );

									end
									else
									if((r_sys_run_step==8'h51)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1204[9:0] );

									end
									else
									if((r_sys_run_step==8'h90)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1960[9:0] );

									end
									else
									if((r_sys_run_step==8'h3b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp940[9:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp568[9:0] );

									end
									else
									if((r_sys_run_step==8'h52)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1216[9:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp460[9:0] );

									end
									else
									if((r_sys_run_step==8'h53)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1228[9:0] );

									end
									else
									if((r_sys_run_step==8'h31)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp820[9:0] );

									end
									else
									if((r_sys_run_step==8'hf) || (r_sys_run_step==8'h11)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp412[9:0] );

									end
									else
									if((r_sys_run_step==8'h2d) || (r_sys_run_step==8'h2f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp772[9:0] );

									end
									else
									if((r_sys_run_step==8'h80)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1768[9:0] );

									end
									else
									if((r_sys_run_step==8'h4d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1156[9:0] );

									end
									else
									if((r_sys_run_step==8'h74)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1624[9:0] );

									end
									else
									if((r_sys_run_step==8'h97)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2044[9:0] );

									end
									else
									if((r_sys_run_step==8'h92)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1984[9:0] );

									end
									else
									if((r_sys_run_step==8'h82)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1792[9:0] );

									end
									else
									if((r_sys_run_step==8'h7a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1696[9:0] );

									end
									else
									if((r_sys_run_step==8'h6b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1516[9:0] );

									end
									else
									if((r_sys_run_step==8'h36) || (r_sys_run_step==8'h38)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp880[9:0] );

									end
									else
									if((r_sys_run_step==8'h1e) || (r_sys_run_step==8'h20)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp592[9:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp688[9:0] );

									end
									else
									if((r_sys_run_step==8'h1f) || (r_sys_run_step==8'h21)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp604[9:0] );

									end
									else
									if((r_sys_run_step==8'h78)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1672[9:0] );

									end
									else
									if((r_sys_run_step==8'h33)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp844[9:0] );

									end
									else
									if((r_sys_run_step==8'h29)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp724[9:0] );

									end
									else
									if((r_sys_run_step==8'h2e) || (r_sys_run_step==8'h30)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp784[9:0] );

									end
									else
									if((r_sys_run_step==8'h5c) || (r_sys_run_step==8'h5e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1336[9:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp640[9:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp484[9:0] );

									end
									else
									if((r_sys_run_step==8'h5a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1312[9:0] );

									end
									else
									if((r_sys_run_step==8'h42)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1024[9:0] );

									end
									else
									if((r_sys_run_step==8'h49)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1108[9:0] );

									end
									else
									if((r_sys_run_step==8'h7f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1756[9:0] );

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp712[9:0] );

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp664[9:0] );

									end
									else
									if((r_sys_run_step==8'h89)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1876[9:0] );

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1480[9:0] );

									end
									else
									if((r_sys_run_step==8'h98)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2056[9:0] );

									end
									else
									if((r_sys_run_step==8'h2c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp760[9:0] );

									end
									else
									if((r_sys_run_step==8'h3d) || (r_sys_run_step==8'h3f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp964[9:0] );

									end
									else
									if((r_sys_run_step==8'h5d) || (r_sys_run_step==8'h5f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1348[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp256[9:0] );

									end
									else
									if((r_sys_run_step==8'h70)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1576[9:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp652[9:0] );

									end
									else
									if((r_sys_run_step==8'h4e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1168[9:0] );

									end
									else
									if((r_sys_run_step==8'h60)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1384[9:0] );

									end
									else
									if((r_sys_run_step==8'h94) || (r_sys_run_step==8'h96)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2008[9:0] );

									end
									else
									if((r_sys_run_step==8'h9a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2080[9:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp364[9:0] );

									end
									else
									if((r_sys_run_step==8'h99)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2068[9:0] );

									end
									else
									if((r_sys_run_step==8'h58)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1288[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp292[9:0] );

									end
									else
									if((r_sys_run_step==8'h17) || (r_sys_run_step==8'h19)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp508[9:0] );

									end
									else
									if((r_sys_run_step==8'h3a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp928[9:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp676[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp280[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp244[9:0] );

									end
									else
									if((r_sys_run_step==8'h3c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp952[9:0] );

									end
									else
									if((r_sys_run_step==8'h4b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1132[9:0] );

									end
									else
									if((r_sys_run_step==8'h4c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1144[9:0] );

									end
									else
									if((r_sys_run_step==8'h8a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1888[9:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp556[9:0] );

									end
									else
									if((r_sys_run_step==8'h6d) || (r_sys_run_step==8'h6f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1540[9:0] );

									end
									else
									if((r_sys_run_step==8'h9b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2092[9:0] );

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp700[9:0] );

									end
									else
									if((r_sys_run_step==8'h54) || (r_sys_run_step==8'h56)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1240[9:0] );

									end
									else
									if((r_sys_run_step==8'h83) || (r_sys_run_step==8'h85)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1804[9:0] );

									end
									else
									if((r_sys_run_step==8'h64) || (r_sys_run_step==8'h66)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1432[9:0] );

									end
									else
									if((r_sys_run_step==8'h4f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1180[9:0] );

									end
									else
									if((r_sys_run_step==8'h73)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1612[9:0] );

									end
									else
									if((r_sys_run_step==8'h32)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp832[9:0] );

									end
									else
									if((r_sys_run_step==8'h59)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1300[9:0] );

									end
									else
									if((r_sys_run_step==8'h62)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1408[9:0] );

									end
									else
									if((r_sys_run_step==8'h34)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp856[9:0] );

									end
									else
									if((r_sys_run_step==8'h43)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1036[9:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp388[9:0] );

									end
									else
									if((r_sys_run_step==8'h4a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1120[9:0] );

									end
									else
									if((r_sys_run_step==8'h6c) || (r_sys_run_step==8'h6e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1528[9:0] );

									end
									else
									if((r_sys_run_step==8'h8b) || (r_sys_run_step==8'h8d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1900[9:0] );

									end
									else
									if((r_sys_run_step==8'h65) || (r_sys_run_step==8'h67)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1444[9:0] );

									end
									else
									if((r_sys_run_step==8'h63)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1420[9:0] );

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2146[9:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2422[9:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2254[9:0] );

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2542[9:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2434[9:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2230[9:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2458[9:0] );

									end
									else
									if((r_sys_run_step==8'h16) || (r_sys_run_step==8'h18)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2374[9:0] );

									end
									else
									if((r_sys_run_step==8'hf) || (r_sys_run_step==8'h11)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2290[9:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2326[9:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2338[9:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2554[9:0] );

									end
									else
									if((r_sys_run_step==8'h1f) || (r_sys_run_step==8'h21)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2482[9:0] );

									end
									else
									if((r_sys_run_step==8'h1e) || (r_sys_run_step==8'h20)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2470[9:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2566[9:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2242[9:0] );

									end
									else
									if((r_sys_run_step==8'h6) || (r_sys_run_step==8'h8)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2182[9:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2266[9:0] );

									end
									else
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'h9)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2194[9:0] );

									end
									else
									if((r_sys_run_step==8'he) || (r_sys_run_step==8'h10)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2278[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2122[9:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2362[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2158[9:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2530[9:0] );

									end
									else
									if((r_sys_run_step==8'h17) || (r_sys_run_step==8'h19)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2386[9:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2518[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2170[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2110[9:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2350[9:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2446[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2134[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h18) || (r_sys_run_step==8'h1a) || (8'h1c<=r_sys_run_step && r_sys_run_step<=8'h20)) begin
										r_fld_U_2_datain_1 <= w_sys_tmp19;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_U_2_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h18) || (r_sys_run_step==8'h1a) || (8'h1c<=r_sys_run_step && r_sys_run_step<=8'h20)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h9b)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h26)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_fld_U_2_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_V_3_addr_1 <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp42[9:0] );

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h8c) || (r_sys_run_step==8'h8e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1912[9:0] );

									end
									else
									if((r_sys_run_step==8'h44)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1048[9:0] );

									end
									else
									if((r_sys_run_step==8'h76)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1648[9:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp472[9:0] );

									end
									else
									if((r_sys_run_step==8'h5b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1324[9:0] );

									end
									else
									if((r_sys_run_step==8'h2a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp736[9:0] );

									end
									else
									if((r_sys_run_step==8'h91)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1972[9:0] );

									end
									else
									if((r_sys_run_step==8'h81)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1780[9:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp544[9:0] );

									end
									else
									if((r_sys_run_step==8'h72)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1600[9:0] );

									end
									else
									if((r_sys_run_step==8'h7b) || (r_sys_run_step==8'h7d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1708[9:0] );

									end
									else
									if((r_sys_run_step==8'h35) || (r_sys_run_step==8'h37)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp868[9:0] );

									end
									else
									if((r_sys_run_step==8'h69)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1492[9:0] );

									end
									else
									if((r_sys_run_step==8'h61)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1396[9:0] );

									end
									else
									if((r_sys_run_step==8'h3e) || (r_sys_run_step==8'h40)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp976[9:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp448[9:0] );

									end
									else
									if((r_sys_run_step==8'he) || (r_sys_run_step==8'h10)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp400[9:0] );

									end
									else
									if((r_sys_run_step==8'h39)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp916[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp268[9:0] );

									end
									else
									if((r_sys_run_step==8'h8f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1948[9:0] );

									end
									else
									if((r_sys_run_step==8'h46) || (r_sys_run_step==8'h48)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1072[9:0] );

									end
									else
									if((r_sys_run_step==8'h71)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1588[9:0] );

									end
									else
									if((r_sys_run_step==8'h79)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1684[9:0] );

									end
									else
									if((r_sys_run_step==8'h2b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp748[9:0] );

									end
									else
									if((r_sys_run_step==8'h55) || (r_sys_run_step==8'h57)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1252[9:0] );

									end
									else
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'h9)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp316[9:0] );

									end
									else
									if((r_sys_run_step==8'h75)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1636[9:0] );

									end
									else
									if((r_sys_run_step==8'h16) || (r_sys_run_step==8'h18)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp496[9:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp352[9:0] );

									end
									else
									if((r_sys_run_step==8'h87)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1852[9:0] );

									end
									else
									if((r_sys_run_step==8'h88)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1864[9:0] );

									end
									else
									if((r_sys_run_step==8'h6) || (r_sys_run_step==8'h8)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp304[9:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp580[9:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp376[9:0] );

									end
									else
									if((r_sys_run_step==8'h6a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1504[9:0] );

									end
									else
									if((r_sys_run_step==8'h41)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1012[9:0] );

									end
									else
									if((r_sys_run_step==8'h50)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1192[9:0] );

									end
									else
									if((r_sys_run_step==8'h7c) || (r_sys_run_step==8'h7e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1720[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp232[9:0] );

									end
									else
									if((r_sys_run_step==8'h77)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1660[9:0] );

									end
									else
									if((r_sys_run_step==8'h45) || (r_sys_run_step==8'h47)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1060[9:0] );

									end
									else
									if((r_sys_run_step==8'h93) || (r_sys_run_step==8'h95)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1996[9:0] );

									end
									else
									if((r_sys_run_step==8'h84) || (r_sys_run_step==8'h86)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1816[9:0] );

									end
									else
									if((r_sys_run_step==8'h51)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1204[9:0] );

									end
									else
									if((r_sys_run_step==8'h90)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1960[9:0] );

									end
									else
									if((r_sys_run_step==8'h3b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp940[9:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp568[9:0] );

									end
									else
									if((r_sys_run_step==8'h52)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1216[9:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp460[9:0] );

									end
									else
									if((r_sys_run_step==8'h53)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1228[9:0] );

									end
									else
									if((r_sys_run_step==8'h31)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp820[9:0] );

									end
									else
									if((r_sys_run_step==8'hf) || (r_sys_run_step==8'h11)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp412[9:0] );

									end
									else
									if((r_sys_run_step==8'h2d) || (r_sys_run_step==8'h2f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp772[9:0] );

									end
									else
									if((r_sys_run_step==8'h80)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1768[9:0] );

									end
									else
									if((r_sys_run_step==8'h4d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1156[9:0] );

									end
									else
									if((r_sys_run_step==8'h74)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1624[9:0] );

									end
									else
									if((r_sys_run_step==8'h97)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2044[9:0] );

									end
									else
									if((r_sys_run_step==8'h92)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1984[9:0] );

									end
									else
									if((r_sys_run_step==8'h82)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1792[9:0] );

									end
									else
									if((r_sys_run_step==8'h7a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1696[9:0] );

									end
									else
									if((r_sys_run_step==8'h6b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1516[9:0] );

									end
									else
									if((r_sys_run_step==8'h36) || (r_sys_run_step==8'h38)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp880[9:0] );

									end
									else
									if((r_sys_run_step==8'h1e) || (r_sys_run_step==8'h20)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp592[9:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp688[9:0] );

									end
									else
									if((r_sys_run_step==8'h1f) || (r_sys_run_step==8'h21)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp604[9:0] );

									end
									else
									if((r_sys_run_step==8'h78)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1672[9:0] );

									end
									else
									if((r_sys_run_step==8'h33)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp844[9:0] );

									end
									else
									if((r_sys_run_step==8'h29)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp724[9:0] );

									end
									else
									if((r_sys_run_step==8'h2e) || (r_sys_run_step==8'h30)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp784[9:0] );

									end
									else
									if((r_sys_run_step==8'h5c) || (r_sys_run_step==8'h5e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1336[9:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp640[9:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp484[9:0] );

									end
									else
									if((r_sys_run_step==8'h5a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1312[9:0] );

									end
									else
									if((r_sys_run_step==8'h42)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1024[9:0] );

									end
									else
									if((r_sys_run_step==8'h49)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1108[9:0] );

									end
									else
									if((r_sys_run_step==8'h7f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1756[9:0] );

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp712[9:0] );

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp664[9:0] );

									end
									else
									if((r_sys_run_step==8'h89)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1876[9:0] );

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1480[9:0] );

									end
									else
									if((r_sys_run_step==8'h98)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2056[9:0] );

									end
									else
									if((r_sys_run_step==8'h2c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp760[9:0] );

									end
									else
									if((r_sys_run_step==8'h3d) || (r_sys_run_step==8'h3f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp964[9:0] );

									end
									else
									if((r_sys_run_step==8'h5d) || (r_sys_run_step==8'h5f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1348[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp256[9:0] );

									end
									else
									if((r_sys_run_step==8'h70)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1576[9:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp652[9:0] );

									end
									else
									if((r_sys_run_step==8'h4e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1168[9:0] );

									end
									else
									if((r_sys_run_step==8'h60)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1384[9:0] );

									end
									else
									if((r_sys_run_step==8'h94) || (r_sys_run_step==8'h96)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2008[9:0] );

									end
									else
									if((r_sys_run_step==8'h9a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2080[9:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp364[9:0] );

									end
									else
									if((r_sys_run_step==8'h99)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2068[9:0] );

									end
									else
									if((r_sys_run_step==8'h58)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1288[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp292[9:0] );

									end
									else
									if((r_sys_run_step==8'h17) || (r_sys_run_step==8'h19)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp508[9:0] );

									end
									else
									if((r_sys_run_step==8'h3a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp928[9:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp676[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp280[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp244[9:0] );

									end
									else
									if((r_sys_run_step==8'h3c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp952[9:0] );

									end
									else
									if((r_sys_run_step==8'h4b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1132[9:0] );

									end
									else
									if((r_sys_run_step==8'h4c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1144[9:0] );

									end
									else
									if((r_sys_run_step==8'h8a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1888[9:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp556[9:0] );

									end
									else
									if((r_sys_run_step==8'h6d) || (r_sys_run_step==8'h6f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1540[9:0] );

									end
									else
									if((r_sys_run_step==8'h9b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2092[9:0] );

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp700[9:0] );

									end
									else
									if((r_sys_run_step==8'h54) || (r_sys_run_step==8'h56)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1240[9:0] );

									end
									else
									if((r_sys_run_step==8'h83) || (r_sys_run_step==8'h85)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1804[9:0] );

									end
									else
									if((r_sys_run_step==8'h64) || (r_sys_run_step==8'h66)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1432[9:0] );

									end
									else
									if((r_sys_run_step==8'h4f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1180[9:0] );

									end
									else
									if((r_sys_run_step==8'h73)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1612[9:0] );

									end
									else
									if((r_sys_run_step==8'h32)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp832[9:0] );

									end
									else
									if((r_sys_run_step==8'h59)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1300[9:0] );

									end
									else
									if((r_sys_run_step==8'h62)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1408[9:0] );

									end
									else
									if((r_sys_run_step==8'h34)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp856[9:0] );

									end
									else
									if((r_sys_run_step==8'h43)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1036[9:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp388[9:0] );

									end
									else
									if((r_sys_run_step==8'h4a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1120[9:0] );

									end
									else
									if((r_sys_run_step==8'h6c) || (r_sys_run_step==8'h6e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1528[9:0] );

									end
									else
									if((r_sys_run_step==8'h8b) || (r_sys_run_step==8'h8d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1900[9:0] );

									end
									else
									if((r_sys_run_step==8'h65) || (r_sys_run_step==8'h67)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1444[9:0] );

									end
									else
									if((r_sys_run_step==8'h63)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1420[9:0] );

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2146[9:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2422[9:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2254[9:0] );

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2542[9:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2434[9:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2230[9:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2458[9:0] );

									end
									else
									if((r_sys_run_step==8'h16) || (r_sys_run_step==8'h18)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2374[9:0] );

									end
									else
									if((r_sys_run_step==8'hf) || (r_sys_run_step==8'h11)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2290[9:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2326[9:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2338[9:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2554[9:0] );

									end
									else
									if((r_sys_run_step==8'h1f) || (r_sys_run_step==8'h21)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2482[9:0] );

									end
									else
									if((r_sys_run_step==8'h1e) || (r_sys_run_step==8'h20)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2470[9:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2566[9:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2242[9:0] );

									end
									else
									if((r_sys_run_step==8'h6) || (r_sys_run_step==8'h8)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2182[9:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2266[9:0] );

									end
									else
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'h9)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2194[9:0] );

									end
									else
									if((r_sys_run_step==8'he) || (r_sys_run_step==8'h10)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2278[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2122[9:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2362[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2158[9:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2530[9:0] );

									end
									else
									if((r_sys_run_step==8'h17) || (r_sys_run_step==8'h19)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2386[9:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2518[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2170[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2110[9:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2350[9:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2446[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2134[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_fld_V_3_datain_1 <= w_sys_tmp26;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_V_3_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h9b)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h26)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_fld_V_3_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_29 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_29 <= w_sys_tmp15;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_29 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h9d)) begin
										r_run_k_29 <= w_sys_tmp2103;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_29 <= w_sys_tmp2104;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h28)) begin
										r_run_k_29 <= w_sys_tmp2577;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_29 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_run_k_29 <= w_sys_tmp2597;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_29 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h9d)) begin
										r_run_k_29 <= w_sys_tmp3674;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_29 <= w_sys_tmp3675;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h28)) begin
										r_run_k_29 <= w_sys_tmp3914;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_29 <= w_sys_tmp3915;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h75)) begin
										r_run_k_29 <= w_sys_tmp4506;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_29 <= w_sys_tmp4507;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1e)) begin
										r_run_k_29 <= w_sys_tmp4663;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_j_30 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_run_j_30 <= w_sys_tmp49;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_j_30 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h2) || (r_sys_run_step==8'h4) || (r_sys_run_step==8'h6) || (r_sys_run_step==8'h8) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'hc)) begin
										r_run_j_30 <= w_sys_tmp2612;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h25)) begin
										r_run_j_30 <= w_sys_tmp2685;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_run_j_30 <= w_sys_tmp2697;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_n_31 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_n_31 <= w_sys_tmp2580;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_mx_32 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_my_33 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_dt_34 <= w_sys_tmp5;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_dx_35 <= w_sys_tmp7;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_dy_36 <= w_sys_tmp8;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_r1_37 <= w_sys_tmp9;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_r2_38 <= w_sys_tmp10;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_r3_39 <= w_sys_tmp11;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_r4_40 <= w_sys_tmp12;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h10) || (r_sys_run_step==8'h11)) begin
										r_run_YY_41 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==8'hc) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h14)) begin
										r_run_YY_41 <= w_sys_tmp19;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_kx_42 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_ky_43 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_nlast_44 <= w_sys_tmp6;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy0_j_45 <= r_run_j_30;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_run_copy0_j_45 <= w_sys_tmp46;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy1_j_46 <= r_run_j_30;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h18) || (r_sys_run_step==8'h1a) || (8'h1c<=r_sys_run_step && r_sys_run_step<=8'h20)) begin
										r_run_copy1_j_46 <= w_sys_tmp47;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy2_j_47 <= r_run_j_30;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_run_copy2_j_47 <= w_sys_tmp48;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy0_j_48 <= r_run_j_30;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1) || (r_sys_run_step==8'h3) || (r_sys_run_step==8'h5) || (r_sys_run_step==8'h7) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'hd)) begin
										r_run_copy0_j_48 <= w_sys_tmp2611;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h13: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub19_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub19_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h9c)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp3663[9:0] );

									end
									else
									if((r_sys_run_step==8'h9d)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp3669[9:0] );

									end
									else
									if((r_sys_run_step==8'h98)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp3627[9:0] );

									end
									else
									if((r_sys_run_step==8'h9b)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp3657[9:0] );

									end
									else
									if((r_sys_run_step==8'h99)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp3645[9:0] );

									end
									else
									if((r_sys_run_step==8'h9a)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp3651[9:0] );

									end
									else
									if((r_sys_run_step==8'h97)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp3621[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h97<=r_sys_run_step && r_sys_run_step<=8'h9d)) begin
										r_sub19_T_datain <= w_sys_tmp2741;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h97<=r_sys_run_step && r_sys_run_step<=8'h9d)) begin
										r_sub19_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub19_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h98)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp2008[9:0] );

									end
									else
									if((r_sys_run_step==8'h9c)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp2080[9:0] );

									end
									else
									if((r_sys_run_step==8'h9b)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp2068[9:0] );

									end
									else
									if((r_sys_run_step==8'h97)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp1996[9:0] );

									end
									else
									if((r_sys_run_step==8'h9a)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp2056[9:0] );

									end
									else
									if((r_sys_run_step==8'h99)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp2044[9:0] );

									end
									else
									if((r_sys_run_step==8'h9d)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp2092[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h97<=r_sys_run_step && r_sys_run_step<=8'h9d)) begin
										r_sub19_V_datain <= w_sys_tmp240;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h97<=r_sys_run_step && r_sys_run_step<=8'h9d)) begin
										r_sub19_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub19_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h98)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp2008[9:0] );

									end
									else
									if((r_sys_run_step==8'h9c)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp2080[9:0] );

									end
									else
									if((r_sys_run_step==8'h9b)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp2068[9:0] );

									end
									else
									if((r_sys_run_step==8'h97)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp1996[9:0] );

									end
									else
									if((r_sys_run_step==8'h9a)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp2056[9:0] );

									end
									else
									if((r_sys_run_step==8'h99)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp2044[9:0] );

									end
									else
									if((r_sys_run_step==8'h9d)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp2092[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h97<=r_sys_run_step && r_sys_run_step<=8'h9d)) begin
										r_sub19_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h97<=r_sys_run_step && r_sys_run_step<=8'h9d)) begin
										r_sub19_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub19_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp4502[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp4497[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp4482[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp4492[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp4487[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h4)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub19_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h9: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub09_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub09_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4b)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp3177[9:0] );

									end
									else
									if((r_sys_run_step==8'h4e)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp3195[9:0] );

									end
									else
									if((r_sys_run_step==8'h4d)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp3189[9:0] );

									end
									else
									if((r_sys_run_step==8'h4c)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp3183[9:0] );

									end
									else
									if((r_sys_run_step==8'h4a)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp3159[9:0] );

									end
									else
									if((r_sys_run_step==8'h49)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp3153[9:0] );

									end
									else
									if((r_sys_run_step==8'h4f)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp3201[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h49<=r_sys_run_step && r_sys_run_step<=8'h4f)) begin
										r_sub09_T_datain <= w_sys_tmp2741;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h49<=r_sys_run_step && r_sys_run_step<=8'h4f)) begin
										r_sub09_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub09_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4e)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp1144[9:0] );

									end
									else
									if((r_sys_run_step==8'h4c)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp1120[9:0] );

									end
									else
									if((r_sys_run_step==8'h4f)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp1156[9:0] );

									end
									else
									if((r_sys_run_step==8'h49)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp1060[9:0] );

									end
									else
									if((r_sys_run_step==8'h4a)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp1072[9:0] );

									end
									else
									if((r_sys_run_step==8'h4d)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp1132[9:0] );

									end
									else
									if((r_sys_run_step==8'h4b)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp1108[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h49<=r_sys_run_step && r_sys_run_step<=8'h4f)) begin
										r_sub09_V_datain <= w_sys_tmp240;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h49<=r_sys_run_step && r_sys_run_step<=8'h4f)) begin
										r_sub09_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub09_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4e)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp1144[9:0] );

									end
									else
									if((r_sys_run_step==8'h4c)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp1120[9:0] );

									end
									else
									if((r_sys_run_step==8'h4f)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp1156[9:0] );

									end
									else
									if((r_sys_run_step==8'h49)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp1060[9:0] );

									end
									else
									if((r_sys_run_step==8'h4a)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp1072[9:0] );

									end
									else
									if((r_sys_run_step==8'h4d)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp1132[9:0] );

									end
									else
									if((r_sys_run_step==8'h4b)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp1108[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h49<=r_sys_run_step && r_sys_run_step<=8'h4f)) begin
										r_sub09_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h49<=r_sys_run_step && r_sys_run_step<=8'h4f)) begin
										r_sub09_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub09_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4207[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4202[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4192[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4197[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4212[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h4)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub09_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h8: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub08_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub08_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h43)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp3129[9:0] );

									end
									else
									if((r_sys_run_step==8'h44)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp3135[9:0] );

									end
									else
									if((r_sys_run_step==8'h42)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp3111[9:0] );

									end
									else
									if((r_sys_run_step==8'h41)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp3105[9:0] );

									end
									else
									if((r_sys_run_step==8'h48)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp3159[9:0] );

									end
									else
									if((r_sys_run_step==8'h47)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp3153[9:0] );

									end
									else
									if((r_sys_run_step==8'h46)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp3147[9:0] );

									end
									else
									if((r_sys_run_step==8'h45)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp3141[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h41<=r_sys_run_step && r_sys_run_step<=8'h48)) begin
										r_sub08_T_datain <= w_sys_tmp2741;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h41<=r_sys_run_step && r_sys_run_step<=8'h48)) begin
										r_sub08_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub08_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h41)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp964[9:0] );

									end
									else
									if((r_sys_run_step==8'h46)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp1048[9:0] );

									end
									else
									if((r_sys_run_step==8'h43)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp1012[9:0] );

									end
									else
									if((r_sys_run_step==8'h45)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp1036[9:0] );

									end
									else
									if((r_sys_run_step==8'h47)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp1060[9:0] );

									end
									else
									if((r_sys_run_step==8'h48)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp1072[9:0] );

									end
									else
									if((r_sys_run_step==8'h44)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp1024[9:0] );

									end
									else
									if((r_sys_run_step==8'h42)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp976[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h41<=r_sys_run_step && r_sys_run_step<=8'h48)) begin
										r_sub08_V_datain <= w_sys_tmp240;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h41<=r_sys_run_step && r_sys_run_step<=8'h48)) begin
										r_sub08_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub08_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h41)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp964[9:0] );

									end
									else
									if((r_sys_run_step==8'h46)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp1048[9:0] );

									end
									else
									if((r_sys_run_step==8'h43)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp1012[9:0] );

									end
									else
									if((r_sys_run_step==8'h45)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp1036[9:0] );

									end
									else
									if((r_sys_run_step==8'h47)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp1060[9:0] );

									end
									else
									if((r_sys_run_step==8'h48)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp1072[9:0] );

									end
									else
									if((r_sys_run_step==8'h44)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp1024[9:0] );

									end
									else
									if((r_sys_run_step==8'h42)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp976[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h41<=r_sys_run_step && r_sys_run_step<=8'h48)) begin
										r_sub08_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h41<=r_sys_run_step && r_sys_run_step<=8'h48)) begin
										r_sub08_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub08_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4162[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4177[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4182[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4187[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4172[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4167[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub08_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h18: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub24_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub24_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h23)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp3867[9:0] );

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp3909[9:0] );

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp3903[9:0] );

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp3885[9:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp3897[9:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp3861[9:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp3891[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h22<=r_sys_run_step && r_sys_run_step<=8'h28)) begin
										r_sub24_T_datain <= w_sys_tmp3683;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h22<=r_sys_run_step && r_sys_run_step<=8'h28)) begin
										r_sub24_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub24_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h28)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp2566[9:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp2530[9:0] );

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp2518[9:0] );

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp2554[9:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp2542[9:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp2482[9:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp2470[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h22<=r_sys_run_step && r_sys_run_step<=8'h28)) begin
										r_sub24_V_datain <= w_sys_tmp2118;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h22<=r_sys_run_step && r_sys_run_step<=8'h28)) begin
										r_sub24_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub24_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h28)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp2566[9:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp2530[9:0] );

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp2518[9:0] );

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp2554[9:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp2542[9:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp2482[9:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp2470[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h22<=r_sys_run_step && r_sys_run_step<=8'h28)) begin
										r_sub24_U_datain <= w_sys_tmp2112;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h22<=r_sys_run_step && r_sys_run_step<=8'h28)) begin
										r_sub24_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub24_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp4659[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp4649[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp4644[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp4654[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp4639[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h4)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub24_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h16: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub22_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub22_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h12)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp3765[9:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp3795[9:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp3789[9:0] );

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp3819[9:0] );

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp3813[9:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp3807[9:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp3771[9:0] );

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp3801[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h12<=r_sys_run_step && r_sys_run_step<=8'h19)) begin
										r_sub22_T_datain <= w_sys_tmp3683;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h12<=r_sys_run_step && r_sys_run_step<=8'h19)) begin
										r_sub22_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub22_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h19)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp2386[9:0] );

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp2374[9:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp2290[9:0] );

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp2350[9:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp2338[9:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp2326[9:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp2278[9:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp2362[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h12<=r_sys_run_step && r_sys_run_step<=8'h19)) begin
										r_sub22_V_datain <= w_sys_tmp2118;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h12<=r_sys_run_step && r_sys_run_step<=8'h19)) begin
										r_sub22_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub22_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h19)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp2386[9:0] );

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp2374[9:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp2290[9:0] );

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp2350[9:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp2338[9:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp2326[9:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp2278[9:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp2362[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h12<=r_sys_run_step && r_sys_run_step<=8'h19)) begin
										r_sub22_U_datain <= w_sys_tmp2112;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h12<=r_sys_run_step && r_sys_run_step<=8'h19)) begin
										r_sub22_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub22_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp4584[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp4589[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp4579[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp4599[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp4594[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp4604[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub22_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h17: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub23_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub23_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h21)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp3867[9:0] );

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp3849[9:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp3819[9:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp3843[9:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp3813[9:0] );

									end
									else
									if((r_sys_run_step==8'h20)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp3861[9:0] );

									end
									else
									if((r_sys_run_step==8'h1f)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp3855[9:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp3837[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h1a<=r_sys_run_step && r_sys_run_step<=8'h21)) begin
										r_sub23_T_datain <= w_sys_tmp3683;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h1a<=r_sys_run_step && r_sys_run_step<=8'h21)) begin
										r_sub23_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub23_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1b)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp2386[9:0] );

									end
									else
									if((r_sys_run_step==8'h1f)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp2458[9:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp2374[9:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp2422[9:0] );

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp2446[9:0] );

									end
									else
									if((r_sys_run_step==8'h21)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp2482[9:0] );

									end
									else
									if((r_sys_run_step==8'h20)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp2470[9:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp2434[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h1a<=r_sys_run_step && r_sys_run_step<=8'h21)) begin
										r_sub23_V_datain <= w_sys_tmp2118;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h1a<=r_sys_run_step && r_sys_run_step<=8'h21)) begin
										r_sub23_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub23_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1b)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp2386[9:0] );

									end
									else
									if((r_sys_run_step==8'h1f)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp2458[9:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp2374[9:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp2422[9:0] );

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp2446[9:0] );

									end
									else
									if((r_sys_run_step==8'h21)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp2482[9:0] );

									end
									else
									if((r_sys_run_step==8'h20)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp2470[9:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp2434[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h1a<=r_sys_run_step && r_sys_run_step<=8'h21)) begin
										r_sub23_U_datain <= w_sys_tmp2112;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h1a<=r_sys_run_step && r_sys_run_step<=8'h21)) begin
										r_sub23_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub23_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp4624[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp4614[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp4629[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp4609[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp4634[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp4619[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub23_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'hc: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub12_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub12_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h61)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp3297[9:0] );

									end
									else
									if((r_sys_run_step==8'h66)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp3339[9:0] );

									end
									else
									if((r_sys_run_step==8'h65)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp3333[9:0] );

									end
									else
									if((r_sys_run_step==8'h67)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp3345[9:0] );

									end
									else
									if((r_sys_run_step==8'h63)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp3321[9:0] );

									end
									else
									if((r_sys_run_step==8'h62)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp3315[9:0] );

									end
									else
									if((r_sys_run_step==8'h64)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp3327[9:0] );

									end
									else
									if((r_sys_run_step==8'h60)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp3291[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h60<=r_sys_run_step && r_sys_run_step<=8'h67)) begin
										r_sub12_T_datain <= w_sys_tmp2741;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h60<=r_sys_run_step && r_sys_run_step<=8'h67)) begin
										r_sub12_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub12_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h61)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp1348[9:0] );

									end
									else
									if((r_sys_run_step==8'h64)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp1408[9:0] );

									end
									else
									if((r_sys_run_step==8'h66)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp1432[9:0] );

									end
									else
									if((r_sys_run_step==8'h60)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp1336[9:0] );

									end
									else
									if((r_sys_run_step==8'h63)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp1396[9:0] );

									end
									else
									if((r_sys_run_step==8'h67)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp1444[9:0] );

									end
									else
									if((r_sys_run_step==8'h65)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp1420[9:0] );

									end
									else
									if((r_sys_run_step==8'h62)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp1384[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h60<=r_sys_run_step && r_sys_run_step<=8'h67)) begin
										r_sub12_V_datain <= w_sys_tmp240;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h60<=r_sys_run_step && r_sys_run_step<=8'h67)) begin
										r_sub12_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub12_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h61)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp1348[9:0] );

									end
									else
									if((r_sys_run_step==8'h64)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp1408[9:0] );

									end
									else
									if((r_sys_run_step==8'h66)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp1432[9:0] );

									end
									else
									if((r_sys_run_step==8'h60)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp1336[9:0] );

									end
									else
									if((r_sys_run_step==8'h63)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp1396[9:0] );

									end
									else
									if((r_sys_run_step==8'h67)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp1444[9:0] );

									end
									else
									if((r_sys_run_step==8'h65)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp1420[9:0] );

									end
									else
									if((r_sys_run_step==8'h62)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp1384[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h60<=r_sys_run_step && r_sys_run_step<=8'h67)) begin
										r_sub12_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h60<=r_sys_run_step && r_sys_run_step<=8'h67)) begin
										r_sub12_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub12_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp4282[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp4292[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp4297[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp4277[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp4287[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp4302[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub12_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h3: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h20)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp2919[9:0] );

									end
									else
									if((r_sys_run_step==8'h1f)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp2913[9:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp2871[9:0] );

									end
									else
									if((r_sys_run_step==8'h21)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp2925[9:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp2895[9:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp2877[9:0] );

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp2907[9:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp2901[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h1a<=r_sys_run_step && r_sys_run_step<=8'h21)) begin
										r_sub03_T_datain <= w_sys_tmp2741;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h1a<=r_sys_run_step && r_sys_run_step<=8'h21)) begin
										r_sub03_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub03_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1c)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp544[9:0] );

									end
									else
									if((r_sys_run_step==8'h1f)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp580[9:0] );

									end
									else
									if((r_sys_run_step==8'h20)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp592[9:0] );

									end
									else
									if((r_sys_run_step==8'h21)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp604[9:0] );

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp568[9:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp496[9:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp508[9:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp556[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h1a<=r_sys_run_step && r_sys_run_step<=8'h21)) begin
										r_sub03_V_datain <= w_sys_tmp240;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h1a<=r_sys_run_step && r_sys_run_step<=8'h21)) begin
										r_sub03_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub03_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1c)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp544[9:0] );

									end
									else
									if((r_sys_run_step==8'h1f)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp580[9:0] );

									end
									else
									if((r_sys_run_step==8'h20)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp592[9:0] );

									end
									else
									if((r_sys_run_step==8'h21)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp604[9:0] );

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp568[9:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp496[9:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp508[9:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp556[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h1a<=r_sys_run_step && r_sys_run_step<=8'h21)) begin
										r_sub03_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h1a<=r_sys_run_step && r_sys_run_step<=8'h21)) begin
										r_sub03_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub03_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4037[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4042[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4027[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4022[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4017[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4032[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub03_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h2: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h17)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp2865[9:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp2829[9:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp2853[9:0] );

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp2871[9:0] );

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp2859[9:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp2847[9:0] );

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp2877[9:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp2823[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h12<=r_sys_run_step && r_sys_run_step<=8'h19)) begin
										r_sub02_T_datain <= w_sys_tmp2741;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h12<=r_sys_run_step && r_sys_run_step<=8'h19)) begin
										r_sub02_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub02_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h14)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp448[9:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp400[9:0] );

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp472[9:0] );

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp496[9:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp460[9:0] );

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp508[9:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp484[9:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp412[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h12<=r_sys_run_step && r_sys_run_step<=8'h19)) begin
										r_sub02_V_datain <= w_sys_tmp240;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h12<=r_sys_run_step && r_sys_run_step<=8'h19)) begin
										r_sub02_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub02_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h14)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp448[9:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp400[9:0] );

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp472[9:0] );

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp496[9:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp460[9:0] );

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp508[9:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp484[9:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp412[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h12<=r_sys_run_step && r_sys_run_step<=8'h19)) begin
										r_sub02_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h12<=r_sys_run_step && r_sys_run_step<=8'h19)) begin
										r_sub02_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub02_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3987[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3997[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp4012[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3992[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp4002[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp4007[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub02_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'hb: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub11_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub11_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5f)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp3297[9:0] );

									end
									else
									if((r_sys_run_step==8'h5b)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp3273[9:0] );

									end
									else
									if((r_sys_run_step==8'h59)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp3249[9:0] );

									end
									else
									if((r_sys_run_step==8'h5c)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp3279[9:0] );

									end
									else
									if((r_sys_run_step==8'h5d)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp3285[9:0] );

									end
									else
									if((r_sys_run_step==8'h5e)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp3291[9:0] );

									end
									else
									if((r_sys_run_step==8'h5a)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp3267[9:0] );

									end
									else
									if((r_sys_run_step==8'h58)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp3243[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h58<=r_sys_run_step && r_sys_run_step<=8'h5f)) begin
										r_sub11_T_datain <= w_sys_tmp2741;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h58<=r_sys_run_step && r_sys_run_step<=8'h5f)) begin
										r_sub11_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub11_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5f)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp1348[9:0] );

									end
									else
									if((r_sys_run_step==8'h5b)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp1300[9:0] );

									end
									else
									if((r_sys_run_step==8'h59)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp1252[9:0] );

									end
									else
									if((r_sys_run_step==8'h5e)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp1336[9:0] );

									end
									else
									if((r_sys_run_step==8'h5d)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp1324[9:0] );

									end
									else
									if((r_sys_run_step==8'h5a)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp1288[9:0] );

									end
									else
									if((r_sys_run_step==8'h5c)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp1312[9:0] );

									end
									else
									if((r_sys_run_step==8'h58)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp1240[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h58<=r_sys_run_step && r_sys_run_step<=8'h5f)) begin
										r_sub11_V_datain <= w_sys_tmp240;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h58<=r_sys_run_step && r_sys_run_step<=8'h5f)) begin
										r_sub11_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub11_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5f)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp1348[9:0] );

									end
									else
									if((r_sys_run_step==8'h5b)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp1300[9:0] );

									end
									else
									if((r_sys_run_step==8'h59)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp1252[9:0] );

									end
									else
									if((r_sys_run_step==8'h5e)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp1336[9:0] );

									end
									else
									if((r_sys_run_step==8'h5d)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp1324[9:0] );

									end
									else
									if((r_sys_run_step==8'h5a)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp1288[9:0] );

									end
									else
									if((r_sys_run_step==8'h5c)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp1312[9:0] );

									end
									else
									if((r_sys_run_step==8'h58)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp1240[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h58<=r_sys_run_step && r_sys_run_step<=8'h5f)) begin
										r_sub11_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h58<=r_sys_run_step && r_sys_run_step<=8'h5f)) begin
										r_sub11_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub11_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp4267[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp4257[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp4252[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp4247[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp4272[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp4262[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub11_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'he: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub14_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub14_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h74)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp3423[9:0] );

									end
									else
									if((r_sys_run_step==8'h71)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp3393[9:0] );

									end
									else
									if((r_sys_run_step==8'h73)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp3417[9:0] );

									end
									else
									if((r_sys_run_step==8'h72)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp3411[9:0] );

									end
									else
									if((r_sys_run_step==8'h70)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp3387[9:0] );

									end
									else
									if((r_sys_run_step==8'h76)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp3435[9:0] );

									end
									else
									if((r_sys_run_step==8'h75)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp3429[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h70<=r_sys_run_step && r_sys_run_step<=8'h76)) begin
										r_sub14_T_datain <= w_sys_tmp2741;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h70<=r_sys_run_step && r_sys_run_step<=8'h76)) begin
										r_sub14_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub14_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h74)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp1600[9:0] );

									end
									else
									if((r_sys_run_step==8'h70)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp1528[9:0] );

									end
									else
									if((r_sys_run_step==8'h72)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp1576[9:0] );

									end
									else
									if((r_sys_run_step==8'h75)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp1612[9:0] );

									end
									else
									if((r_sys_run_step==8'h76)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp1624[9:0] );

									end
									else
									if((r_sys_run_step==8'h73)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp1588[9:0] );

									end
									else
									if((r_sys_run_step==8'h71)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp1540[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h70<=r_sys_run_step && r_sys_run_step<=8'h76)) begin
										r_sub14_V_datain <= w_sys_tmp240;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h70<=r_sys_run_step && r_sys_run_step<=8'h76)) begin
										r_sub14_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub14_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h74)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp1600[9:0] );

									end
									else
									if((r_sys_run_step==8'h70)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp1528[9:0] );

									end
									else
									if((r_sys_run_step==8'h72)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp1576[9:0] );

									end
									else
									if((r_sys_run_step==8'h75)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp1612[9:0] );

									end
									else
									if((r_sys_run_step==8'h76)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp1624[9:0] );

									end
									else
									if((r_sys_run_step==8'h73)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp1588[9:0] );

									end
									else
									if((r_sys_run_step==8'h71)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp1540[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h70<=r_sys_run_step && r_sys_run_step<=8'h76)) begin
										r_sub14_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h70<=r_sys_run_step && r_sys_run_step<=8'h76)) begin
										r_sub14_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub14_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp4347[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp4342[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp4337[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp4357[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp4352[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h4)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub14_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'ha)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp2775[9:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp2781[9:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp2829[9:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp2805[9:0] );

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp2811[9:0] );

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp2823[9:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp2817[9:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp2799[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'ha<=r_sys_run_step && r_sys_run_step<=8'h11)) begin
										r_sub01_T_datain <= w_sys_tmp2741;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'ha<=r_sys_run_step && r_sys_run_step<=8'h11)) begin
										r_sub01_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub01_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'ha)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp304[9:0] );

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp400[9:0] );

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp376[9:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp388[9:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp316[9:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp364[9:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp352[9:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp412[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'ha<=r_sys_run_step && r_sys_run_step<=8'h11)) begin
										r_sub01_V_datain <= w_sys_tmp240;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'ha<=r_sys_run_step && r_sys_run_step<=8'h11)) begin
										r_sub01_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub01_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'ha)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp304[9:0] );

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp400[9:0] );

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp376[9:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp388[9:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp316[9:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp364[9:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp352[9:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp412[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'ha<=r_sys_run_step && r_sys_run_step<=8'h11)) begin
										r_sub01_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'ha<=r_sys_run_step && r_sys_run_step<=8'h11)) begin
										r_sub01_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub01_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3982[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3977[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3972[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3962[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3967[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3957[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h8)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp2775[9:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp2781[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp2757[9:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp2763[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp2739[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp2745[9:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp2769[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp2751[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h9)) begin
										r_sub00_T_datain <= w_sys_tmp2741;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h9)) begin
										r_sub00_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub00_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h8)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp304[9:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp280[9:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp316[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp256[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp244[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp232[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp268[9:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp292[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h9)) begin
										r_sub00_V_datain <= w_sys_tmp240;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h9)) begin
										r_sub00_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub00_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h8)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp304[9:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp280[9:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp316[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp256[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp244[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp232[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp268[9:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp292[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h9)) begin
										r_sub00_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h9)) begin
										r_sub00_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub00_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3939[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3921[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3951[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3945[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3933[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3927[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'hd: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub13_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub13_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6f)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp3393[9:0] );

									end
									else
									if((r_sys_run_step==8'h6c)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp3375[9:0] );

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp3339[9:0] );

									end
									else
									if((r_sys_run_step==8'h69)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp3345[9:0] );

									end
									else
									if((r_sys_run_step==8'h6b)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp3369[9:0] );

									end
									else
									if((r_sys_run_step==8'h6e)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp3387[9:0] );

									end
									else
									if((r_sys_run_step==8'h6a)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp3363[9:0] );

									end
									else
									if((r_sys_run_step==8'h6d)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp3381[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h68<=r_sys_run_step && r_sys_run_step<=8'h6f)) begin
										r_sub13_T_datain <= w_sys_tmp2741;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h68<=r_sys_run_step && r_sys_run_step<=8'h6f)) begin
										r_sub13_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub13_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6d)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp1516[9:0] );

									end
									else
									if((r_sys_run_step==8'h6c)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp1504[9:0] );

									end
									else
									if((r_sys_run_step==8'h6b)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp1492[9:0] );

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp1432[9:0] );

									end
									else
									if((r_sys_run_step==8'h6e)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp1528[9:0] );

									end
									else
									if((r_sys_run_step==8'h69)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp1444[9:0] );

									end
									else
									if((r_sys_run_step==8'h6a)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp1480[9:0] );

									end
									else
									if((r_sys_run_step==8'h6f)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp1540[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h68<=r_sys_run_step && r_sys_run_step<=8'h6f)) begin
										r_sub13_V_datain <= w_sys_tmp240;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h68<=r_sys_run_step && r_sys_run_step<=8'h6f)) begin
										r_sub13_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub13_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6d)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp1516[9:0] );

									end
									else
									if((r_sys_run_step==8'h6c)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp1504[9:0] );

									end
									else
									if((r_sys_run_step==8'h6b)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp1492[9:0] );

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp1432[9:0] );

									end
									else
									if((r_sys_run_step==8'h6e)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp1528[9:0] );

									end
									else
									if((r_sys_run_step==8'h69)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp1444[9:0] );

									end
									else
									if((r_sys_run_step==8'h6a)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp1480[9:0] );

									end
									else
									if((r_sys_run_step==8'h6f)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp1540[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h68<=r_sys_run_step && r_sys_run_step<=8'h6f)) begin
										r_sub13_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h68<=r_sys_run_step && r_sys_run_step<=8'h6f)) begin
										r_sub13_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub13_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp4332[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp4307[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp4312[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp4317[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp4322[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp4327[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub13_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h7: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub07_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub07_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3d)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp3093[9:0] );

									end
									else
									if((r_sys_run_step==8'h3e)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp3099[9:0] );

									end
									else
									if((r_sys_run_step==8'h40)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp3111[9:0] );

									end
									else
									if((r_sys_run_step==8'h3f)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp3105[9:0] );

									end
									else
									if((r_sys_run_step==8'h39)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp3057[9:0] );

									end
									else
									if((r_sys_run_step==8'h3b)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp3081[9:0] );

									end
									else
									if((r_sys_run_step==8'h3a)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp3063[9:0] );

									end
									else
									if((r_sys_run_step==8'h3c)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp3087[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h39<=r_sys_run_step && r_sys_run_step<=8'h40)) begin
										r_sub07_T_datain <= w_sys_tmp2741;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h39<=r_sys_run_step && r_sys_run_step<=8'h40)) begin
										r_sub07_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub07_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3f)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp964[9:0] );

									end
									else
									if((r_sys_run_step==8'h3c)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp928[9:0] );

									end
									else
									if((r_sys_run_step==8'h3a)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp880[9:0] );

									end
									else
									if((r_sys_run_step==8'h39)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp868[9:0] );

									end
									else
									if((r_sys_run_step==8'h3d)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp940[9:0] );

									end
									else
									if((r_sys_run_step==8'h3b)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp916[9:0] );

									end
									else
									if((r_sys_run_step==8'h3e)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp952[9:0] );

									end
									else
									if((r_sys_run_step==8'h40)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp976[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h39<=r_sys_run_step && r_sys_run_step<=8'h40)) begin
										r_sub07_V_datain <= w_sys_tmp240;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h39<=r_sys_run_step && r_sys_run_step<=8'h40)) begin
										r_sub07_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub07_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3f)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp964[9:0] );

									end
									else
									if((r_sys_run_step==8'h3c)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp928[9:0] );

									end
									else
									if((r_sys_run_step==8'h3a)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp880[9:0] );

									end
									else
									if((r_sys_run_step==8'h39)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp868[9:0] );

									end
									else
									if((r_sys_run_step==8'h3d)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp940[9:0] );

									end
									else
									if((r_sys_run_step==8'h3b)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp916[9:0] );

									end
									else
									if((r_sys_run_step==8'h3e)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp952[9:0] );

									end
									else
									if((r_sys_run_step==8'h40)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp976[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h39<=r_sys_run_step && r_sys_run_step<=8'h40)) begin
										r_sub07_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h39<=r_sys_run_step && r_sys_run_step<=8'h40)) begin
										r_sub07_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub07_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4137[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4132[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4147[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4152[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4157[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4142[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub07_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h10: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub16_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub16_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h84)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp3519[9:0] );

									end
									else
									if((r_sys_run_step==8'h82)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp3507[9:0] );

									end
									else
									if((r_sys_run_step==8'h81)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp3501[9:0] );

									end
									else
									if((r_sys_run_step==8'h85)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp3525[9:0] );

									end
									else
									if((r_sys_run_step==8'h7f)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp3477[9:0] );

									end
									else
									if((r_sys_run_step==8'h80)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp3483[9:0] );

									end
									else
									if((r_sys_run_step==8'h86)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp3531[9:0] );

									end
									else
									if((r_sys_run_step==8'h83)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp3513[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h7f<=r_sys_run_step && r_sys_run_step<=8'h86)) begin
										r_sub16_T_datain <= w_sys_tmp2741;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h7f<=r_sys_run_step && r_sys_run_step<=8'h86)) begin
										r_sub16_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub16_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h81)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp1756[9:0] );

									end
									else
									if((r_sys_run_step==8'h7f)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp1708[9:0] );

									end
									else
									if((r_sys_run_step==8'h85)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp1804[9:0] );

									end
									else
									if((r_sys_run_step==8'h80)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp1720[9:0] );

									end
									else
									if((r_sys_run_step==8'h82)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp1768[9:0] );

									end
									else
									if((r_sys_run_step==8'h86)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp1816[9:0] );

									end
									else
									if((r_sys_run_step==8'h84)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp1792[9:0] );

									end
									else
									if((r_sys_run_step==8'h83)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp1780[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h7f<=r_sys_run_step && r_sys_run_step<=8'h86)) begin
										r_sub16_V_datain <= w_sys_tmp240;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h7f<=r_sys_run_step && r_sys_run_step<=8'h86)) begin
										r_sub16_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub16_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h81)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp1756[9:0] );

									end
									else
									if((r_sys_run_step==8'h7f)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp1708[9:0] );

									end
									else
									if((r_sys_run_step==8'h85)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp1804[9:0] );

									end
									else
									if((r_sys_run_step==8'h80)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp1720[9:0] );

									end
									else
									if((r_sys_run_step==8'h82)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp1768[9:0] );

									end
									else
									if((r_sys_run_step==8'h86)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp1816[9:0] );

									end
									else
									if((r_sys_run_step==8'h84)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp1792[9:0] );

									end
									else
									if((r_sys_run_step==8'h83)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp1780[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h7f<=r_sys_run_step && r_sys_run_step<=8'h86)) begin
										r_sub16_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h7f<=r_sys_run_step && r_sys_run_step<=8'h86)) begin
										r_sub16_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub16_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp4407[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp4417[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp4412[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp4402[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp4397[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp4392[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub16_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h6: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub06_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub06_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h34)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp3039[9:0] );

									end
									else
									if((r_sys_run_step==8'h32)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp3015[9:0] );

									end
									else
									if((r_sys_run_step==8'h31)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp3009[9:0] );

									end
									else
									if((r_sys_run_step==8'h35)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp3045[9:0] );

									end
									else
									if((r_sys_run_step==8'h36)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp3051[9:0] );

									end
									else
									if((r_sys_run_step==8'h37)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp3057[9:0] );

									end
									else
									if((r_sys_run_step==8'h33)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp3033[9:0] );

									end
									else
									if((r_sys_run_step==8'h38)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp3063[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h31<=r_sys_run_step && r_sys_run_step<=8'h38)) begin
										r_sub06_T_datain <= w_sys_tmp2741;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h31<=r_sys_run_step && r_sys_run_step<=8'h38)) begin
										r_sub06_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub06_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h34)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp832[9:0] );

									end
									else
									if((r_sys_run_step==8'h38)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp880[9:0] );

									end
									else
									if((r_sys_run_step==8'h35)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp844[9:0] );

									end
									else
									if((r_sys_run_step==8'h37)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp868[9:0] );

									end
									else
									if((r_sys_run_step==8'h31)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp772[9:0] );

									end
									else
									if((r_sys_run_step==8'h36)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp856[9:0] );

									end
									else
									if((r_sys_run_step==8'h32)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp784[9:0] );

									end
									else
									if((r_sys_run_step==8'h33)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp820[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h31<=r_sys_run_step && r_sys_run_step<=8'h38)) begin
										r_sub06_V_datain <= w_sys_tmp240;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h31<=r_sys_run_step && r_sys_run_step<=8'h38)) begin
										r_sub06_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub06_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h34)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp832[9:0] );

									end
									else
									if((r_sys_run_step==8'h38)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp880[9:0] );

									end
									else
									if((r_sys_run_step==8'h35)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp844[9:0] );

									end
									else
									if((r_sys_run_step==8'h37)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp868[9:0] );

									end
									else
									if((r_sys_run_step==8'h31)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp772[9:0] );

									end
									else
									if((r_sys_run_step==8'h36)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp856[9:0] );

									end
									else
									if((r_sys_run_step==8'h32)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp784[9:0] );

									end
									else
									if((r_sys_run_step==8'h33)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp820[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h31<=r_sys_run_step && r_sys_run_step<=8'h38)) begin
										r_sub06_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h31<=r_sys_run_step && r_sys_run_step<=8'h38)) begin
										r_sub06_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub06_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4102[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4117[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4127[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4122[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4107[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4112[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub06_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub15_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub15_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h77)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp3441[9:0] );

									end
									else
									if((r_sys_run_step==8'h78)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp3447[9:0] );

									end
									else
									if((r_sys_run_step==8'h7a)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp3459[9:0] );

									end
									else
									if((r_sys_run_step==8'h7d)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp3477[9:0] );

									end
									else
									if((r_sys_run_step==8'h7c)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp3471[9:0] );

									end
									else
									if((r_sys_run_step==8'h7b)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp3465[9:0] );

									end
									else
									if((r_sys_run_step==8'h7e)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp3483[9:0] );

									end
									else
									if((r_sys_run_step==8'h79)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp3453[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h77<=r_sys_run_step && r_sys_run_step<=8'h7e)) begin
										r_sub15_T_datain <= w_sys_tmp2741;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h77<=r_sys_run_step && r_sys_run_step<=8'h7e)) begin
										r_sub15_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub15_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7c)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp1696[9:0] );

									end
									else
									if((r_sys_run_step==8'h7b)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp1684[9:0] );

									end
									else
									if((r_sys_run_step==8'h7d)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp1708[9:0] );

									end
									else
									if((r_sys_run_step==8'h7e)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp1720[9:0] );

									end
									else
									if((r_sys_run_step==8'h78)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp1648[9:0] );

									end
									else
									if((r_sys_run_step==8'h77)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp1636[9:0] );

									end
									else
									if((r_sys_run_step==8'h79)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp1660[9:0] );

									end
									else
									if((r_sys_run_step==8'h7a)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp1672[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h77<=r_sys_run_step && r_sys_run_step<=8'h7e)) begin
										r_sub15_V_datain <= w_sys_tmp240;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h77<=r_sys_run_step && r_sys_run_step<=8'h7e)) begin
										r_sub15_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub15_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7c)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp1696[9:0] );

									end
									else
									if((r_sys_run_step==8'h7b)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp1684[9:0] );

									end
									else
									if((r_sys_run_step==8'h7d)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp1708[9:0] );

									end
									else
									if((r_sys_run_step==8'h7e)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp1720[9:0] );

									end
									else
									if((r_sys_run_step==8'h78)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp1648[9:0] );

									end
									else
									if((r_sys_run_step==8'h77)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp1636[9:0] );

									end
									else
									if((r_sys_run_step==8'h79)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp1660[9:0] );

									end
									else
									if((r_sys_run_step==8'h7a)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp1672[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h77<=r_sys_run_step && r_sys_run_step<=8'h7e)) begin
										r_sub15_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h77<=r_sys_run_step && r_sys_run_step<=8'h7e)) begin
										r_sub15_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub15_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp4367[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp4387[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp4362[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp4382[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp4377[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp4372[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub15_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h5: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub05_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub05_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2b)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp2985[9:0] );

									end
									else
									if((r_sys_run_step==8'h30)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp3015[9:0] );

									end
									else
									if((r_sys_run_step==8'h2f)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp3009[9:0] );

									end
									else
									if((r_sys_run_step==8'h2c)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp2991[9:0] );

									end
									else
									if((r_sys_run_step==8'h2e)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp3003[9:0] );

									end
									else
									if((r_sys_run_step==8'h2a)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp2979[9:0] );

									end
									else
									if((r_sys_run_step==8'h29)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp2973[9:0] );

									end
									else
									if((r_sys_run_step==8'h2d)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp2997[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h29<=r_sys_run_step && r_sys_run_step<=8'h30)) begin
										r_sub05_T_datain <= w_sys_tmp2741;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h29<=r_sys_run_step && r_sys_run_step<=8'h30)) begin
										r_sub05_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub05_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2d)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp748[9:0] );

									end
									else
									if((r_sys_run_step==8'h2f)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp772[9:0] );

									end
									else
									if((r_sys_run_step==8'h2b)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp724[9:0] );

									end
									else
									if((r_sys_run_step==8'h30)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp784[9:0] );

									end
									else
									if((r_sys_run_step==8'h2a)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp712[9:0] );

									end
									else
									if((r_sys_run_step==8'h2c)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp736[9:0] );

									end
									else
									if((r_sys_run_step==8'h2e)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp760[9:0] );

									end
									else
									if((r_sys_run_step==8'h29)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp700[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h29<=r_sys_run_step && r_sys_run_step<=8'h30)) begin
										r_sub05_V_datain <= w_sys_tmp240;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h29<=r_sys_run_step && r_sys_run_step<=8'h30)) begin
										r_sub05_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub05_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2d)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp748[9:0] );

									end
									else
									if((r_sys_run_step==8'h2f)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp772[9:0] );

									end
									else
									if((r_sys_run_step==8'h2b)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp724[9:0] );

									end
									else
									if((r_sys_run_step==8'h30)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp784[9:0] );

									end
									else
									if((r_sys_run_step==8'h2a)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp712[9:0] );

									end
									else
									if((r_sys_run_step==8'h2c)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp736[9:0] );

									end
									else
									if((r_sys_run_step==8'h2e)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp760[9:0] );

									end
									else
									if((r_sys_run_step==8'h29)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp700[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h29<=r_sys_run_step && r_sys_run_step<=8'h30)) begin
										r_sub05_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h29<=r_sys_run_step && r_sys_run_step<=8'h30)) begin
										r_sub05_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub05_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4087[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4097[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4092[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4082[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4072[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4077[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub05_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h12: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub18_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub18_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h94)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp3615[9:0] );

									end
									else
									if((r_sys_run_step==8'h8f)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp3573[9:0] );

									end
									else
									if((r_sys_run_step==8'h93)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp3609[9:0] );

									end
									else
									if((r_sys_run_step==8'h90)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp3579[9:0] );

									end
									else
									if((r_sys_run_step==8'h91)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp3597[9:0] );

									end
									else
									if((r_sys_run_step==8'h96)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp3627[9:0] );

									end
									else
									if((r_sys_run_step==8'h95)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp3621[9:0] );

									end
									else
									if((r_sys_run_step==8'h92)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp3603[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h8f<=r_sys_run_step && r_sys_run_step<=8'h96)) begin
										r_sub18_T_datain <= w_sys_tmp2741;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h8f<=r_sys_run_step && r_sys_run_step<=8'h96)) begin
										r_sub18_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub18_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h96)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp2008[9:0] );

									end
									else
									if((r_sys_run_step==8'h90)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp1912[9:0] );

									end
									else
									if((r_sys_run_step==8'h92)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp1960[9:0] );

									end
									else
									if((r_sys_run_step==8'h8f)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp1900[9:0] );

									end
									else
									if((r_sys_run_step==8'h93)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp1972[9:0] );

									end
									else
									if((r_sys_run_step==8'h91)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp1948[9:0] );

									end
									else
									if((r_sys_run_step==8'h95)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp1996[9:0] );

									end
									else
									if((r_sys_run_step==8'h94)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp1984[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h8f<=r_sys_run_step && r_sys_run_step<=8'h96)) begin
										r_sub18_V_datain <= w_sys_tmp240;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h8f<=r_sys_run_step && r_sys_run_step<=8'h96)) begin
										r_sub18_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub18_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h96)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp2008[9:0] );

									end
									else
									if((r_sys_run_step==8'h90)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp1912[9:0] );

									end
									else
									if((r_sys_run_step==8'h92)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp1960[9:0] );

									end
									else
									if((r_sys_run_step==8'h8f)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp1900[9:0] );

									end
									else
									if((r_sys_run_step==8'h93)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp1972[9:0] );

									end
									else
									if((r_sys_run_step==8'h91)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp1948[9:0] );

									end
									else
									if((r_sys_run_step==8'h95)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp1996[9:0] );

									end
									else
									if((r_sys_run_step==8'h94)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp1984[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h8f<=r_sys_run_step && r_sys_run_step<=8'h96)) begin
										r_sub18_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h8f<=r_sys_run_step && r_sys_run_step<=8'h96)) begin
										r_sub18_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub18_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp4477[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp4457[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp4462[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp4472[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp4467[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp4452[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub18_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h4: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub04_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub04_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h22)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp2919[9:0] );

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp2961[9:0] );

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp2967[9:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp2949[9:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp2955[9:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp2925[9:0] );

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp2943[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h22<=r_sys_run_step && r_sys_run_step<=8'h28)) begin
										r_sub04_T_datain <= w_sys_tmp2741;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h22<=r_sys_run_step && r_sys_run_step<=8'h28)) begin
										r_sub04_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub04_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h27)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp676[9:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp592[9:0] );

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp688[9:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp604[9:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp664[9:0] );

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp640[9:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp652[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h22<=r_sys_run_step && r_sys_run_step<=8'h28)) begin
										r_sub04_V_datain <= w_sys_tmp240;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h22<=r_sys_run_step && r_sys_run_step<=8'h28)) begin
										r_sub04_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub04_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h27)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp676[9:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp592[9:0] );

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp688[9:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp604[9:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp664[9:0] );

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp640[9:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp652[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h22<=r_sys_run_step && r_sys_run_step<=8'h28)) begin
										r_sub04_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h22<=r_sys_run_step && r_sys_run_step<=8'h28)) begin
										r_sub04_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub04_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4052[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4067[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4062[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4057[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4047[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h4)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub04_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h11: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub17_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub17_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h8d)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp3573[9:0] );

									end
									else
									if((r_sys_run_step==8'h89)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp3549[9:0] );

									end
									else
									if((r_sys_run_step==8'h8a)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp3555[9:0] );

									end
									else
									if((r_sys_run_step==8'h8b)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp3561[9:0] );

									end
									else
									if((r_sys_run_step==8'h8e)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp3579[9:0] );

									end
									else
									if((r_sys_run_step==8'h87)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp3525[9:0] );

									end
									else
									if((r_sys_run_step==8'h8c)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp3567[9:0] );

									end
									else
									if((r_sys_run_step==8'h88)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp3531[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h87<=r_sys_run_step && r_sys_run_step<=8'h8e)) begin
										r_sub17_T_datain <= w_sys_tmp2741;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h87<=r_sys_run_step && r_sys_run_step<=8'h8e)) begin
										r_sub17_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub17_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h8a)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp1864[9:0] );

									end
									else
									if((r_sys_run_step==8'h8e)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp1912[9:0] );

									end
									else
									if((r_sys_run_step==8'h87)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp1804[9:0] );

									end
									else
									if((r_sys_run_step==8'h8d)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp1900[9:0] );

									end
									else
									if((r_sys_run_step==8'h8c)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp1888[9:0] );

									end
									else
									if((r_sys_run_step==8'h8b)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp1876[9:0] );

									end
									else
									if((r_sys_run_step==8'h89)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp1852[9:0] );

									end
									else
									if((r_sys_run_step==8'h88)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp1816[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h87<=r_sys_run_step && r_sys_run_step<=8'h8e)) begin
										r_sub17_V_datain <= w_sys_tmp240;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h87<=r_sys_run_step && r_sys_run_step<=8'h8e)) begin
										r_sub17_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub17_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h8a)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp1864[9:0] );

									end
									else
									if((r_sys_run_step==8'h8e)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp1912[9:0] );

									end
									else
									if((r_sys_run_step==8'h87)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp1804[9:0] );

									end
									else
									if((r_sys_run_step==8'h8d)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp1900[9:0] );

									end
									else
									if((r_sys_run_step==8'h8c)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp1888[9:0] );

									end
									else
									if((r_sys_run_step==8'h8b)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp1876[9:0] );

									end
									else
									if((r_sys_run_step==8'h89)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp1852[9:0] );

									end
									else
									if((r_sys_run_step==8'h88)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp1816[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h87<=r_sys_run_step && r_sys_run_step<=8'h8e)) begin
										r_sub17_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h87<=r_sys_run_step && r_sys_run_step<=8'h8e)) begin
										r_sub17_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub17_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp4447[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp4442[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp4427[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp4432[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp4437[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp4422[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub17_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'ha: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub10_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub10_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h52)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp3219[9:0] );

									end
									else
									if((r_sys_run_step==8'h55)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp3237[9:0] );

									end
									else
									if((r_sys_run_step==8'h53)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp3225[9:0] );

									end
									else
									if((r_sys_run_step==8'h50)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp3207[9:0] );

									end
									else
									if((r_sys_run_step==8'h57)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp3249[9:0] );

									end
									else
									if((r_sys_run_step==8'h51)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp3213[9:0] );

									end
									else
									if((r_sys_run_step==8'h56)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp3243[9:0] );

									end
									else
									if((r_sys_run_step==8'h54)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp3231[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h50<=r_sys_run_step && r_sys_run_step<=8'h57)) begin
										r_sub10_T_datain <= w_sys_tmp2741;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h50<=r_sys_run_step && r_sys_run_step<=8'h57)) begin
										r_sub10_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub10_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h52)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp1192[9:0] );

									end
									else
									if((r_sys_run_step==8'h57)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp1252[9:0] );

									end
									else
									if((r_sys_run_step==8'h51)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp1180[9:0] );

									end
									else
									if((r_sys_run_step==8'h54)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp1216[9:0] );

									end
									else
									if((r_sys_run_step==8'h55)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp1228[9:0] );

									end
									else
									if((r_sys_run_step==8'h53)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp1204[9:0] );

									end
									else
									if((r_sys_run_step==8'h50)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp1168[9:0] );

									end
									else
									if((r_sys_run_step==8'h56)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp1240[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h50<=r_sys_run_step && r_sys_run_step<=8'h57)) begin
										r_sub10_V_datain <= w_sys_tmp240;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h50<=r_sys_run_step && r_sys_run_step<=8'h57)) begin
										r_sub10_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub10_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h52)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp1192[9:0] );

									end
									else
									if((r_sys_run_step==8'h57)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp1252[9:0] );

									end
									else
									if((r_sys_run_step==8'h51)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp1180[9:0] );

									end
									else
									if((r_sys_run_step==8'h54)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp1216[9:0] );

									end
									else
									if((r_sys_run_step==8'h55)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp1228[9:0] );

									end
									else
									if((r_sys_run_step==8'h53)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp1204[9:0] );

									end
									else
									if((r_sys_run_step==8'h50)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp1168[9:0] );

									end
									else
									if((r_sys_run_step==8'h56)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp1240[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h50<=r_sys_run_step && r_sys_run_step<=8'h57)) begin
										r_sub10_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h50<=r_sys_run_step && r_sys_run_step<=8'h57)) begin
										r_sub10_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub10_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp4237[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp4232[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp4242[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp4222[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp4227[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp4217[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub10_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h14: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub20_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub20_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp3693[9:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp3705[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp3681[9:0] );

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp3717[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp3699[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp3687[9:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp3711[9:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp3723[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h9)) begin
										r_sub20_T_datain <= w_sys_tmp3683;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h9)) begin
										r_sub20_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub20_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp2146[9:0] );

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp2182[9:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp2158[9:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp2170[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp2110[9:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp2194[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp2122[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp2134[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h9)) begin
										r_sub20_V_datain <= w_sys_tmp2118;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h9)) begin
										r_sub20_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub20_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp2146[9:0] );

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp2182[9:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp2158[9:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp2170[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp2110[9:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp2194[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp2122[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp2134[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h9)) begin
										r_sub20_U_datain <= w_sys_tmp2112;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h9)) begin
										r_sub20_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub20_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp4543[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp4513[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp4537[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp4531[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp4525[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp4519[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub20_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h15: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub21_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub21_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h10)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp3765[9:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp3759[9:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp3717[9:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp3741[9:0] );

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp3753[9:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp3747[9:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp3771[9:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp3723[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'ha<=r_sys_run_step && r_sys_run_step<=8'h11)) begin
										r_sub21_T_datain <= w_sys_tmp3683;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'ha<=r_sys_run_step && r_sys_run_step<=8'h11)) begin
										r_sub21_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub21_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'hd)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp2242[9:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp2230[9:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp2182[9:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp2266[9:0] );

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp2254[9:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp2290[9:0] );

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp2278[9:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp2194[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'ha<=r_sys_run_step && r_sys_run_step<=8'h11)) begin
										r_sub21_V_datain <= w_sys_tmp2118;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'ha<=r_sys_run_step && r_sys_run_step<=8'h11)) begin
										r_sub21_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub21_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'hd)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp2242[9:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp2230[9:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp2182[9:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp2266[9:0] );

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp2254[9:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp2290[9:0] );

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp2278[9:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp2194[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'ha<=r_sys_run_step && r_sys_run_step<=8'h11)) begin
										r_sub21_U_datain <= w_sys_tmp2112;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'ha<=r_sys_run_step && r_sys_run_step<=8'h11)) begin
										r_sub21_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub21_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp4564[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp4574[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp4569[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp4549[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp4554[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp4559[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub21_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h16)) begin
										r_sys_tmp0_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp0_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h16)) begin
										r_sys_tmp1_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp1_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h12) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h19)) begin
										r_sys_tmp2_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp2_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h11) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h17)) begin
										r_sys_tmp3_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp3_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'hf) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h19)) begin
										r_sys_tmp4_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==8'hc) || (r_sys_run_step==8'hd)) begin
										r_sys_tmp4_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp4_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp5_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp5_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp6_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp6_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp7_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp7_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp8_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp8_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp9_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp9_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp10_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp10_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp11_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp11_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp12_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp12_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp13_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp13_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp14_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp14_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp15_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp15_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp16_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp16_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp17_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp17_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp18_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp18_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp19_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp19_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp20_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp20_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp21_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp21_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp22_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp22_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp23_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp23_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp24_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp24_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp25_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp25_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp26_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp26_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp27_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp27_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp28_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp29_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp30_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp31_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp32_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp33_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp34_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp35_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp36_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp37_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp38_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp39_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp40_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp41_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp42_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp43_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp44_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp45_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp46_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp47_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp48_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp49_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp50_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp51_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp52_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp53_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp54_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp55_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp56_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp57_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp58_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp59_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp60_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp61_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp62_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp63_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp64_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp65_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp66_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp67_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp68_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp69_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp70_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp71_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp72_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp73_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp74_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp75_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp76_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp77_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp78_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp79_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp80_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp81_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp82_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp83_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp84_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp85_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp86_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp87_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp88_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp89_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp90_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp91_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp92_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp93_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp94_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp95_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp96_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp97_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp98_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp99_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp100_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp101_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp102_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp103_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp104_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp105_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp106_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp107_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp108_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp109_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
