/*
TimeStamp:	2016/6/27		14:41
*/


module c1(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy	
);

	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 5:0] r_sys_run_phase;
	reg         [ 3:0] r_sys_run_stage;
	reg         [ 6:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 3:0] w_sys_run_stage_p1;
	wire        [ 6:0] w_sys_run_step_p1;
	wire signed [ 8:0] w_fld_u_0_addr_0;
	wire        [31:0] w_fld_u_0_datain_0;
	wire        [31:0] w_fld_u_0_dataout_0;
	wire               w_fld_u_0_r_w_0;
	wire               w_fld_u_0_ce_0;
	reg  signed [ 8:0] r_fld_u_0_addr_1;
	reg         [31:0] r_fld_u_0_datain_1;
	wire        [31:0] w_fld_u_0_dataout_1;
	reg                r_fld_u_0_r_w_1;
	wire               w_fld_u_0_ce_1;
	wire signed [ 8:0] w_fld_uu_1_addr_0;
	wire        [31:0] w_fld_uu_1_datain_0;
	wire        [31:0] w_fld_uu_1_dataout_0;
	wire               w_fld_uu_1_r_w_0;
	wire               w_fld_uu_1_ce_0;
	reg  signed [ 8:0] r_fld_uu_1_addr_1;
	reg         [31:0] r_fld_uu_1_datain_1;
	wire        [31:0] w_fld_uu_1_dataout_1;
	reg                r_fld_uu_1_r_w_1;
	wire               w_fld_uu_1_ce_1;
	reg  signed [31:0] r_run_k_11;
	reg  signed [31:0] r_run_j_12;
	reg  signed [31:0] r_run_n_13;
	reg  signed [31:0] r_run_mx_14;
	reg  signed [31:0] r_run_my_15;
	reg  signed [31:0] r_run_nlast_16;
	reg  signed [31:0] r_run_copy0_j_17;
	reg  signed [31:0] r_run_copy0_j_18;
	reg  signed [31:0] r_run_copy1_j_19;
	reg  signed [31:0] r_run_copy2_j_20;
	reg                r_sub08_run_req;
	wire               w_sub08_run_busy;
	wire signed [ 9:0] w_sub08_u_addr;
	reg  signed [ 9:0] r_sub08_u_addr;
	wire        [31:0] w_sub08_u_datain;
	reg         [31:0] r_sub08_u_datain;
	wire        [31:0] w_sub08_u_dataout;
	wire               w_sub08_u_r_w;
	reg                r_sub08_u_r_w;
	wire signed [ 9:0] w_sub08_result_addr;
	reg  signed [ 9:0] r_sub08_result_addr;
	wire        [31:0] w_sub08_result_datain;
	reg         [31:0] r_sub08_result_datain;
	wire        [31:0] w_sub08_result_dataout;
	wire               w_sub08_result_r_w;
	reg                r_sub08_result_r_w;
	reg                r_sub03_run_req;
	wire               w_sub03_run_busy;
	wire signed [ 9:0] w_sub03_u_addr;
	reg  signed [ 9:0] r_sub03_u_addr;
	wire        [31:0] w_sub03_u_datain;
	reg         [31:0] r_sub03_u_datain;
	wire        [31:0] w_sub03_u_dataout;
	wire               w_sub03_u_r_w;
	reg                r_sub03_u_r_w;
	wire signed [ 9:0] w_sub03_result_addr;
	reg  signed [ 9:0] r_sub03_result_addr;
	wire        [31:0] w_sub03_result_datain;
	reg         [31:0] r_sub03_result_datain;
	wire        [31:0] w_sub03_result_dataout;
	wire               w_sub03_result_r_w;
	reg                r_sub03_result_r_w;
	reg                r_sub02_run_req;
	wire               w_sub02_run_busy;
	wire signed [ 9:0] w_sub02_u_addr;
	reg  signed [ 9:0] r_sub02_u_addr;
	wire        [31:0] w_sub02_u_datain;
	reg         [31:0] r_sub02_u_datain;
	wire        [31:0] w_sub02_u_dataout;
	wire               w_sub02_u_r_w;
	reg                r_sub02_u_r_w;
	wire signed [ 9:0] w_sub02_result_addr;
	reg  signed [ 9:0] r_sub02_result_addr;
	wire        [31:0] w_sub02_result_datain;
	reg         [31:0] r_sub02_result_datain;
	wire        [31:0] w_sub02_result_dataout;
	wire               w_sub02_result_r_w;
	reg                r_sub02_result_r_w;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [ 9:0] w_sub01_u_addr;
	reg  signed [ 9:0] r_sub01_u_addr;
	wire        [31:0] w_sub01_u_datain;
	reg         [31:0] r_sub01_u_datain;
	wire        [31:0] w_sub01_u_dataout;
	wire               w_sub01_u_r_w;
	reg                r_sub01_u_r_w;
	wire signed [ 9:0] w_sub01_result_addr;
	reg  signed [ 9:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [ 9:0] w_sub00_u_addr;
	reg  signed [ 9:0] r_sub00_u_addr;
	wire        [31:0] w_sub00_u_datain;
	reg         [31:0] r_sub00_u_datain;
	wire        [31:0] w_sub00_u_dataout;
	wire               w_sub00_u_r_w;
	reg                r_sub00_u_r_w;
	wire signed [ 9:0] w_sub00_result_addr;
	reg  signed [ 9:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	reg                r_sub07_run_req;
	wire               w_sub07_run_busy;
	wire signed [ 9:0] w_sub07_u_addr;
	reg  signed [ 9:0] r_sub07_u_addr;
	wire        [31:0] w_sub07_u_datain;
	reg         [31:0] r_sub07_u_datain;
	wire        [31:0] w_sub07_u_dataout;
	wire               w_sub07_u_r_w;
	reg                r_sub07_u_r_w;
	wire signed [ 9:0] w_sub07_result_addr;
	reg  signed [ 9:0] r_sub07_result_addr;
	wire        [31:0] w_sub07_result_datain;
	reg         [31:0] r_sub07_result_datain;
	wire        [31:0] w_sub07_result_dataout;
	wire               w_sub07_result_r_w;
	reg                r_sub07_result_r_w;
	reg                r_sub06_run_req;
	wire               w_sub06_run_busy;
	wire signed [ 9:0] w_sub06_u_addr;
	reg  signed [ 9:0] r_sub06_u_addr;
	wire        [31:0] w_sub06_u_datain;
	reg         [31:0] r_sub06_u_datain;
	wire        [31:0] w_sub06_u_dataout;
	wire               w_sub06_u_r_w;
	reg                r_sub06_u_r_w;
	wire signed [ 9:0] w_sub06_result_addr;
	reg  signed [ 9:0] r_sub06_result_addr;
	wire        [31:0] w_sub06_result_datain;
	reg         [31:0] r_sub06_result_datain;
	wire        [31:0] w_sub06_result_dataout;
	wire               w_sub06_result_r_w;
	reg                r_sub06_result_r_w;
	reg                r_sub05_run_req;
	wire               w_sub05_run_busy;
	wire signed [ 9:0] w_sub05_u_addr;
	reg  signed [ 9:0] r_sub05_u_addr;
	wire        [31:0] w_sub05_u_datain;
	reg         [31:0] r_sub05_u_datain;
	wire        [31:0] w_sub05_u_dataout;
	wire               w_sub05_u_r_w;
	reg                r_sub05_u_r_w;
	wire signed [ 9:0] w_sub05_result_addr;
	reg  signed [ 9:0] r_sub05_result_addr;
	wire        [31:0] w_sub05_result_datain;
	reg         [31:0] r_sub05_result_datain;
	wire        [31:0] w_sub05_result_dataout;
	wire               w_sub05_result_r_w;
	reg                r_sub05_result_r_w;
	reg                r_sub04_run_req;
	wire               w_sub04_run_busy;
	wire signed [ 9:0] w_sub04_u_addr;
	reg  signed [ 9:0] r_sub04_u_addr;
	wire        [31:0] w_sub04_u_datain;
	reg         [31:0] r_sub04_u_datain;
	wire        [31:0] w_sub04_u_dataout;
	wire               w_sub04_u_r_w;
	reg                r_sub04_u_r_w;
	wire signed [ 9:0] w_sub04_result_addr;
	reg  signed [ 9:0] r_sub04_result_addr;
	wire        [31:0] w_sub04_result_datain;
	reg         [31:0] r_sub04_result_datain;
	wire        [31:0] w_sub04_result_dataout;
	wire               w_sub04_result_r_w;
	reg                r_sub04_result_r_w;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg         [31:0] r_sys_tmp4_float;
	reg         [31:0] r_sys_tmp5_float;
	reg         [31:0] r_sys_tmp6_float;
	reg         [31:0] r_sys_tmp7_float;
	reg         [31:0] r_sys_tmp8_float;
	reg         [31:0] r_sys_tmp9_float;
	reg         [31:0] r_sys_tmp10_float;
	reg         [31:0] r_sys_tmp11_float;
	reg         [31:0] r_sys_tmp12_float;
	reg         [31:0] r_sys_tmp13_float;
	reg         [31:0] r_sys_tmp14_float;
	reg         [31:0] r_sys_tmp15_float;
	reg         [31:0] r_sys_tmp16_float;
	reg         [31:0] r_sys_tmp17_float;
	reg         [31:0] r_sys_tmp18_float;
	reg         [31:0] r_sys_tmp19_float;
	reg         [31:0] r_sys_tmp20_float;
	reg         [31:0] r_sys_tmp21_float;
	reg         [31:0] r_sys_tmp22_float;
	reg         [31:0] r_sys_tmp23_float;
	reg         [31:0] r_sys_tmp24_float;
	reg         [31:0] r_sys_tmp25_float;
	reg         [31:0] r_sys_tmp26_float;
	reg         [31:0] r_sys_tmp27_float;
	reg         [31:0] r_sys_tmp28_float;
	reg         [31:0] r_sys_tmp29_float;
	reg         [31:0] r_sys_tmp30_float;
	reg         [31:0] r_sys_tmp31_float;
	reg         [31:0] r_sys_tmp32_float;
	reg         [31:0] r_sys_tmp33_float;
	reg         [31:0] r_sys_tmp34_float;
	reg         [31:0] r_sys_tmp35_float;
	reg         [31:0] r_sys_tmp36_float;
	reg         [31:0] r_sys_tmp37_float;
	reg         [31:0] r_sys_tmp38_float;
	reg         [31:0] r_sys_tmp39_float;
	reg         [31:0] r_sys_tmp40_float;
	reg         [31:0] r_sys_tmp41_float;
	reg         [31:0] r_sys_tmp42_float;
	reg         [31:0] r_sys_tmp43_float;
	reg         [31:0] r_sys_tmp44_float;
	reg         [31:0] r_sys_tmp45_float;
	reg         [31:0] r_sys_tmp46_float;
	reg         [31:0] r_sys_tmp47_float;
	wire signed [31:0] w_sys_tmp1;
	wire signed [31:0] w_sys_tmp3;
	wire               w_sys_tmp4;
	wire               w_sys_tmp5;
	wire signed [31:0] w_sys_tmp6;
	wire               w_sys_tmp7;
	wire               w_sys_tmp8;
	wire signed [31:0] w_sys_tmp11;
	wire signed [31:0] w_sys_tmp12;
	wire signed [31:0] w_sys_tmp13;
	wire        [31:0] w_sys_tmp14;
	wire signed [31:0] w_sys_tmp16;
	wire signed [31:0] w_sys_tmp17;
	wire signed [31:0] w_sys_tmp20;
	wire signed [31:0] w_sys_tmp21;
	wire               w_sys_tmp250;
	wire               w_sys_tmp251;
	wire signed [31:0] w_sys_tmp252;
	wire               w_sys_tmp253;
	wire               w_sys_tmp254;
	wire signed [31:0] w_sys_tmp257;
	wire signed [31:0] w_sys_tmp258;
	wire        [31:0] w_sys_tmp259;
	wire signed [31:0] w_sys_tmp261;
	wire signed [31:0] w_sys_tmp262;
	wire        [31:0] w_sys_tmp263;
	wire signed [31:0] w_sys_tmp265;
	wire signed [31:0] w_sys_tmp266;
	wire        [31:0] w_sys_tmp268;
	wire signed [31:0] w_sys_tmp270;
	wire signed [31:0] w_sys_tmp271;
	wire signed [31:0] w_sys_tmp274;
	wire signed [31:0] w_sys_tmp275;
	wire signed [31:0] w_sys_tmp276;
	wire signed [31:0] w_sys_tmp277;
	wire               w_sys_tmp696;
	wire               w_sys_tmp697;
	wire signed [31:0] w_sys_tmp698;
	wire signed [31:0] w_sys_tmp701;
	wire signed [31:0] w_sys_tmp702;
	wire        [31:0] w_sys_tmp703;
	wire signed [31:0] w_sys_tmp707;
	wire signed [31:0] w_sys_tmp708;
	wire signed [31:0] w_sys_tmp713;
	wire signed [31:0] w_sys_tmp714;
	wire signed [31:0] w_sys_tmp719;
	wire signed [31:0] w_sys_tmp720;
	wire signed [31:0] w_sys_tmp725;
	wire signed [31:0] w_sys_tmp726;
	wire signed [31:0] w_sys_tmp731;
	wire signed [31:0] w_sys_tmp732;
	wire signed [31:0] w_sys_tmp737;
	wire signed [31:0] w_sys_tmp738;
	wire signed [31:0] w_sys_tmp743;
	wire signed [31:0] w_sys_tmp744;
	wire signed [31:0] w_sys_tmp749;
	wire signed [31:0] w_sys_tmp750;
	wire signed [31:0] w_sys_tmp755;
	wire signed [31:0] w_sys_tmp756;
	wire signed [31:0] w_sys_tmp761;
	wire signed [31:0] w_sys_tmp762;
	wire signed [31:0] w_sys_tmp767;
	wire signed [31:0] w_sys_tmp768;
	wire signed [31:0] w_sys_tmp785;
	wire signed [31:0] w_sys_tmp786;
	wire signed [31:0] w_sys_tmp791;
	wire signed [31:0] w_sys_tmp792;
	wire signed [31:0] w_sys_tmp797;
	wire signed [31:0] w_sys_tmp798;
	wire signed [31:0] w_sys_tmp803;
	wire signed [31:0] w_sys_tmp804;
	wire signed [31:0] w_sys_tmp809;
	wire signed [31:0] w_sys_tmp810;
	wire signed [31:0] w_sys_tmp815;
	wire signed [31:0] w_sys_tmp816;
	wire signed [31:0] w_sys_tmp821;
	wire signed [31:0] w_sys_tmp822;
	wire signed [31:0] w_sys_tmp827;
	wire signed [31:0] w_sys_tmp828;
	wire signed [31:0] w_sys_tmp833;
	wire signed [31:0] w_sys_tmp834;
	wire signed [31:0] w_sys_tmp839;
	wire signed [31:0] w_sys_tmp840;
	wire signed [31:0] w_sys_tmp857;
	wire signed [31:0] w_sys_tmp858;
	wire signed [31:0] w_sys_tmp863;
	wire signed [31:0] w_sys_tmp864;
	wire signed [31:0] w_sys_tmp869;
	wire signed [31:0] w_sys_tmp870;
	wire signed [31:0] w_sys_tmp875;
	wire signed [31:0] w_sys_tmp876;
	wire signed [31:0] w_sys_tmp881;
	wire signed [31:0] w_sys_tmp882;
	wire signed [31:0] w_sys_tmp887;
	wire signed [31:0] w_sys_tmp888;
	wire signed [31:0] w_sys_tmp893;
	wire signed [31:0] w_sys_tmp894;
	wire signed [31:0] w_sys_tmp899;
	wire signed [31:0] w_sys_tmp900;
	wire signed [31:0] w_sys_tmp905;
	wire signed [31:0] w_sys_tmp906;
	wire signed [31:0] w_sys_tmp911;
	wire signed [31:0] w_sys_tmp912;
	wire signed [31:0] w_sys_tmp917;
	wire signed [31:0] w_sys_tmp918;
	wire signed [31:0] w_sys_tmp923;
	wire signed [31:0] w_sys_tmp924;
	wire signed [31:0] w_sys_tmp929;
	wire signed [31:0] w_sys_tmp930;
	wire signed [31:0] w_sys_tmp935;
	wire signed [31:0] w_sys_tmp936;
	wire signed [31:0] w_sys_tmp941;
	wire signed [31:0] w_sys_tmp942;
	wire signed [31:0] w_sys_tmp947;
	wire signed [31:0] w_sys_tmp948;
	wire signed [31:0] w_sys_tmp953;
	wire signed [31:0] w_sys_tmp954;
	wire signed [31:0] w_sys_tmp959;
	wire signed [31:0] w_sys_tmp960;
	wire signed [31:0] w_sys_tmp965;
	wire signed [31:0] w_sys_tmp966;
	wire signed [31:0] w_sys_tmp971;
	wire signed [31:0] w_sys_tmp972;
	wire signed [31:0] w_sys_tmp977;
	wire signed [31:0] w_sys_tmp978;
	wire signed [31:0] w_sys_tmp995;
	wire signed [31:0] w_sys_tmp996;
	wire signed [31:0] w_sys_tmp1001;
	wire signed [31:0] w_sys_tmp1002;
	wire signed [31:0] w_sys_tmp1007;
	wire signed [31:0] w_sys_tmp1008;
	wire signed [31:0] w_sys_tmp1013;
	wire signed [31:0] w_sys_tmp1014;
	wire signed [31:0] w_sys_tmp1019;
	wire signed [31:0] w_sys_tmp1020;
	wire signed [31:0] w_sys_tmp1025;
	wire signed [31:0] w_sys_tmp1026;
	wire signed [31:0] w_sys_tmp1031;
	wire signed [31:0] w_sys_tmp1032;
	wire signed [31:0] w_sys_tmp1037;
	wire signed [31:0] w_sys_tmp1038;
	wire signed [31:0] w_sys_tmp1043;
	wire signed [31:0] w_sys_tmp1044;
	wire signed [31:0] w_sys_tmp1049;
	wire signed [31:0] w_sys_tmp1050;
	wire signed [31:0] w_sys_tmp1067;
	wire signed [31:0] w_sys_tmp1068;
	wire signed [31:0] w_sys_tmp1073;
	wire signed [31:0] w_sys_tmp1074;
	wire signed [31:0] w_sys_tmp1079;
	wire signed [31:0] w_sys_tmp1080;
	wire signed [31:0] w_sys_tmp1085;
	wire signed [31:0] w_sys_tmp1086;
	wire signed [31:0] w_sys_tmp1091;
	wire signed [31:0] w_sys_tmp1092;
	wire signed [31:0] w_sys_tmp1097;
	wire signed [31:0] w_sys_tmp1098;
	wire signed [31:0] w_sys_tmp1103;
	wire signed [31:0] w_sys_tmp1104;
	wire signed [31:0] w_sys_tmp1109;
	wire signed [31:0] w_sys_tmp1110;
	wire signed [31:0] w_sys_tmp1115;
	wire signed [31:0] w_sys_tmp1116;
	wire signed [31:0] w_sys_tmp1120;
	wire signed [31:0] w_sys_tmp1121;
	wire               w_sys_tmp1122;
	wire               w_sys_tmp1123;
	wire signed [31:0] w_sys_tmp1124;
	wire signed [31:0] w_sys_tmp1127;
	wire signed [31:0] w_sys_tmp1128;
	wire        [31:0] w_sys_tmp1129;
	wire signed [31:0] w_sys_tmp1133;
	wire signed [31:0] w_sys_tmp1134;
	wire signed [31:0] w_sys_tmp1139;
	wire signed [31:0] w_sys_tmp1140;
	wire signed [31:0] w_sys_tmp1145;
	wire signed [31:0] w_sys_tmp1146;
	wire signed [31:0] w_sys_tmp1151;
	wire signed [31:0] w_sys_tmp1152;
	wire signed [31:0] w_sys_tmp1157;
	wire signed [31:0] w_sys_tmp1158;
	wire signed [31:0] w_sys_tmp1163;
	wire signed [31:0] w_sys_tmp1164;
	wire signed [31:0] w_sys_tmp1169;
	wire signed [31:0] w_sys_tmp1170;
	wire signed [31:0] w_sys_tmp1175;
	wire signed [31:0] w_sys_tmp1176;
	wire signed [31:0] w_sys_tmp1181;
	wire signed [31:0] w_sys_tmp1182;
	wire signed [31:0] w_sys_tmp1187;
	wire signed [31:0] w_sys_tmp1188;
	wire signed [31:0] w_sys_tmp1193;
	wire signed [31:0] w_sys_tmp1194;
	wire signed [31:0] w_sys_tmp1211;
	wire signed [31:0] w_sys_tmp1212;
	wire signed [31:0] w_sys_tmp1217;
	wire signed [31:0] w_sys_tmp1218;
	wire signed [31:0] w_sys_tmp1223;
	wire signed [31:0] w_sys_tmp1224;
	wire signed [31:0] w_sys_tmp1229;
	wire signed [31:0] w_sys_tmp1230;
	wire signed [31:0] w_sys_tmp1235;
	wire signed [31:0] w_sys_tmp1236;
	wire signed [31:0] w_sys_tmp1241;
	wire signed [31:0] w_sys_tmp1242;
	wire signed [31:0] w_sys_tmp1247;
	wire signed [31:0] w_sys_tmp1248;
	wire signed [31:0] w_sys_tmp1253;
	wire signed [31:0] w_sys_tmp1254;
	wire signed [31:0] w_sys_tmp1259;
	wire signed [31:0] w_sys_tmp1260;
	wire signed [31:0] w_sys_tmp1271;
	wire signed [31:0] w_sys_tmp1272;
	wire signed [31:0] w_sys_tmp1277;
	wire signed [31:0] w_sys_tmp1278;
	wire signed [31:0] w_sys_tmp1283;
	wire signed [31:0] w_sys_tmp1284;
	wire signed [31:0] w_sys_tmp1289;
	wire signed [31:0] w_sys_tmp1290;
	wire signed [31:0] w_sys_tmp1295;
	wire signed [31:0] w_sys_tmp1296;
	wire signed [31:0] w_sys_tmp1301;
	wire signed [31:0] w_sys_tmp1302;
	wire signed [31:0] w_sys_tmp1307;
	wire signed [31:0] w_sys_tmp1308;
	wire signed [31:0] w_sys_tmp1313;
	wire signed [31:0] w_sys_tmp1314;
	wire signed [31:0] w_sys_tmp1319;
	wire signed [31:0] w_sys_tmp1320;
	wire signed [31:0] w_sys_tmp1324;
	wire signed [31:0] w_sys_tmp1325;
	wire               w_sys_tmp1326;
	wire               w_sys_tmp1327;
	wire signed [31:0] w_sys_tmp1328;
	wire signed [31:0] w_sys_tmp1331;
	wire signed [31:0] w_sys_tmp1332;
	wire        [31:0] w_sys_tmp1333;
	wire signed [31:0] w_sys_tmp1337;
	wire signed [31:0] w_sys_tmp1338;
	wire signed [31:0] w_sys_tmp1343;
	wire signed [31:0] w_sys_tmp1344;
	wire signed [31:0] w_sys_tmp1349;
	wire signed [31:0] w_sys_tmp1350;
	wire signed [31:0] w_sys_tmp1355;
	wire signed [31:0] w_sys_tmp1356;
	wire signed [31:0] w_sys_tmp1361;
	wire signed [31:0] w_sys_tmp1362;
	wire signed [31:0] w_sys_tmp1367;
	wire signed [31:0] w_sys_tmp1368;
	wire signed [31:0] w_sys_tmp1373;
	wire signed [31:0] w_sys_tmp1374;
	wire signed [31:0] w_sys_tmp1379;
	wire signed [31:0] w_sys_tmp1380;
	wire signed [31:0] w_sys_tmp1385;
	wire signed [31:0] w_sys_tmp1386;
	wire signed [31:0] w_sys_tmp1391;
	wire signed [31:0] w_sys_tmp1392;
	wire signed [31:0] w_sys_tmp1396;
	wire signed [31:0] w_sys_tmp1397;
	wire signed [31:0] w_sys_tmp1401;
	wire signed [31:0] w_sys_tmp1402;
	wire signed [31:0] w_sys_tmp1406;
	wire signed [31:0] w_sys_tmp1407;
	wire signed [31:0] w_sys_tmp1411;
	wire signed [31:0] w_sys_tmp1412;
	wire signed [31:0] w_sys_tmp1416;
	wire signed [31:0] w_sys_tmp1417;
	wire signed [31:0] w_sys_tmp1421;
	wire signed [31:0] w_sys_tmp1422;
	wire signed [31:0] w_sys_tmp1426;
	wire signed [31:0] w_sys_tmp1427;
	wire signed [31:0] w_sys_tmp1431;
	wire signed [31:0] w_sys_tmp1432;
	wire signed [31:0] w_sys_tmp1436;
	wire signed [31:0] w_sys_tmp1437;
	wire signed [31:0] w_sys_tmp1441;
	wire signed [31:0] w_sys_tmp1442;
	wire signed [31:0] w_sys_tmp1446;
	wire signed [31:0] w_sys_tmp1447;
	wire signed [31:0] w_sys_tmp1451;
	wire signed [31:0] w_sys_tmp1452;
	wire signed [31:0] w_sys_tmp1456;
	wire signed [31:0] w_sys_tmp1457;
	wire signed [31:0] w_sys_tmp1461;
	wire signed [31:0] w_sys_tmp1462;
	wire signed [31:0] w_sys_tmp1466;
	wire signed [31:0] w_sys_tmp1467;
	wire signed [31:0] w_sys_tmp1471;
	wire signed [31:0] w_sys_tmp1472;
	wire signed [31:0] w_sys_tmp1476;
	wire signed [31:0] w_sys_tmp1477;
	wire signed [31:0] w_sys_tmp1481;
	wire signed [31:0] w_sys_tmp1482;
	wire signed [31:0] w_sys_tmp1486;
	wire signed [31:0] w_sys_tmp1487;
	wire signed [31:0] w_sys_tmp1491;
	wire signed [31:0] w_sys_tmp1492;
	wire signed [31:0] w_sys_tmp1496;
	wire signed [31:0] w_sys_tmp1497;
	wire signed [31:0] w_sys_tmp1501;
	wire signed [31:0] w_sys_tmp1502;
	wire signed [31:0] w_sys_tmp1506;
	wire signed [31:0] w_sys_tmp1507;
	wire signed [31:0] w_sys_tmp1511;
	wire signed [31:0] w_sys_tmp1512;
	wire signed [31:0] w_sys_tmp1516;
	wire signed [31:0] w_sys_tmp1517;
	wire signed [31:0] w_sys_tmp1521;
	wire signed [31:0] w_sys_tmp1522;
	wire signed [31:0] w_sys_tmp1526;
	wire signed [31:0] w_sys_tmp1527;
	wire signed [31:0] w_sys_tmp1531;
	wire signed [31:0] w_sys_tmp1532;
	wire signed [31:0] w_sys_tmp1536;
	wire signed [31:0] w_sys_tmp1537;
	wire signed [31:0] w_sys_tmp1541;
	wire signed [31:0] w_sys_tmp1542;
	wire signed [31:0] w_sys_tmp1546;
	wire signed [31:0] w_sys_tmp1547;
	wire signed [31:0] w_sys_tmp1551;
	wire signed [31:0] w_sys_tmp1552;
	wire signed [31:0] w_sys_tmp1556;
	wire signed [31:0] w_sys_tmp1557;
	wire signed [31:0] w_sys_tmp1561;
	wire signed [31:0] w_sys_tmp1562;
	wire signed [31:0] w_sys_tmp1566;
	wire signed [31:0] w_sys_tmp1567;
	wire signed [31:0] w_sys_tmp1571;
	wire signed [31:0] w_sys_tmp1572;
	wire signed [31:0] w_sys_tmp1576;
	wire signed [31:0] w_sys_tmp1577;
	wire signed [31:0] w_sys_tmp1581;
	wire signed [31:0] w_sys_tmp1582;
	wire signed [31:0] w_sys_tmp1586;
	wire signed [31:0] w_sys_tmp1587;
	wire signed [31:0] w_sys_tmp1591;
	wire signed [31:0] w_sys_tmp1592;
	wire signed [31:0] w_sys_tmp1596;
	wire signed [31:0] w_sys_tmp1597;
	wire signed [31:0] w_sys_tmp1601;
	wire signed [31:0] w_sys_tmp1602;
	wire signed [31:0] w_sys_tmp1606;
	wire signed [31:0] w_sys_tmp1607;
	wire signed [31:0] w_sys_tmp1611;
	wire signed [31:0] w_sys_tmp1612;
	wire signed [31:0] w_sys_tmp1616;
	wire signed [31:0] w_sys_tmp1617;
	wire signed [31:0] w_sys_tmp1621;
	wire signed [31:0] w_sys_tmp1622;
	wire signed [31:0] w_sys_tmp1626;
	wire signed [31:0] w_sys_tmp1627;
	wire signed [31:0] w_sys_tmp1630;
	wire signed [31:0] w_sys_tmp1631;
	wire               w_sys_tmp1632;
	wire               w_sys_tmp1633;
	wire signed [31:0] w_sys_tmp1634;
	wire signed [31:0] w_sys_tmp1637;
	wire signed [31:0] w_sys_tmp1638;
	wire        [31:0] w_sys_tmp1639;
	wire signed [31:0] w_sys_tmp1643;
	wire signed [31:0] w_sys_tmp1644;
	wire signed [31:0] w_sys_tmp1649;
	wire signed [31:0] w_sys_tmp1650;
	wire signed [31:0] w_sys_tmp1655;
	wire signed [31:0] w_sys_tmp1656;
	wire signed [31:0] w_sys_tmp1661;
	wire signed [31:0] w_sys_tmp1662;
	wire signed [31:0] w_sys_tmp1667;
	wire signed [31:0] w_sys_tmp1668;
	wire signed [31:0] w_sys_tmp1673;
	wire signed [31:0] w_sys_tmp1674;
	wire signed [31:0] w_sys_tmp1679;
	wire signed [31:0] w_sys_tmp1680;
	wire signed [31:0] w_sys_tmp1685;
	wire signed [31:0] w_sys_tmp1686;
	wire signed [31:0] w_sys_tmp1691;
	wire signed [31:0] w_sys_tmp1692;
	wire signed [31:0] w_sys_tmp1697;
	wire signed [31:0] w_sys_tmp1698;
	wire signed [31:0] w_sys_tmp1702;
	wire signed [31:0] w_sys_tmp1703;
	wire signed [31:0] w_sys_tmp1707;
	wire signed [31:0] w_sys_tmp1708;
	wire signed [31:0] w_sys_tmp1712;
	wire signed [31:0] w_sys_tmp1713;
	wire signed [31:0] w_sys_tmp1717;
	wire signed [31:0] w_sys_tmp1718;
	wire signed [31:0] w_sys_tmp1722;
	wire signed [31:0] w_sys_tmp1723;
	wire signed [31:0] w_sys_tmp1727;
	wire signed [31:0] w_sys_tmp1728;
	wire signed [31:0] w_sys_tmp1732;
	wire signed [31:0] w_sys_tmp1733;
	wire signed [31:0] w_sys_tmp1737;
	wire signed [31:0] w_sys_tmp1738;
	wire signed [31:0] w_sys_tmp1742;
	wire signed [31:0] w_sys_tmp1743;
	wire signed [31:0] w_sys_tmp1747;
	wire signed [31:0] w_sys_tmp1748;
	wire signed [31:0] w_sys_tmp1757;
	wire signed [31:0] w_sys_tmp1758;
	wire signed [31:0] w_sys_tmp1762;
	wire signed [31:0] w_sys_tmp1763;
	wire signed [31:0] w_sys_tmp1767;
	wire signed [31:0] w_sys_tmp1768;
	wire signed [31:0] w_sys_tmp1772;
	wire signed [31:0] w_sys_tmp1773;
	wire signed [31:0] w_sys_tmp1777;
	wire signed [31:0] w_sys_tmp1778;
	wire signed [31:0] w_sys_tmp1782;
	wire signed [31:0] w_sys_tmp1783;
	wire signed [31:0] w_sys_tmp1787;
	wire signed [31:0] w_sys_tmp1788;
	wire signed [31:0] w_sys_tmp1792;
	wire signed [31:0] w_sys_tmp1793;
	wire signed [31:0] w_sys_tmp1796;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 4'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 7'h1);
	assign w_fld_u_0_addr_0 = 9'sh0;
	assign w_fld_u_0_datain_0 = 32'h0;
	assign w_fld_u_0_r_w_0 = 1'h0;
	assign w_fld_u_0_ce_0 = w_sys_ce;
	assign w_fld_u_0_ce_1 = w_sys_ce;
	assign w_fld_uu_1_addr_0 = 9'sh0;
	assign w_fld_uu_1_datain_0 = 32'h0;
	assign w_fld_uu_1_r_w_0 = 1'h0;
	assign w_fld_uu_1_ce_0 = w_sys_ce;
	assign w_fld_uu_1_ce_1 = w_sys_ce;
	assign w_sub08_u_addr = ( (|r_sys_processing_methodID) ? r_sub08_u_addr : 10'sh0 ) ;
	assign w_sub08_u_datain = ( (|r_sys_processing_methodID) ? r_sub08_u_datain : 32'h0 ) ;
	assign w_sub08_u_r_w = ( (|r_sys_processing_methodID) ? r_sub08_u_r_w : 1'h0 ) ;
	assign w_sub08_result_addr = ( (|r_sys_processing_methodID) ? r_sub08_result_addr : 10'sh0 ) ;
	assign w_sub08_result_datain = ( (|r_sys_processing_methodID) ? r_sub08_result_datain : 32'h0 ) ;
	assign w_sub08_result_r_w = ( (|r_sys_processing_methodID) ? r_sub08_result_r_w : 1'h0 ) ;
	assign w_sub03_u_addr = ( (|r_sys_processing_methodID) ? r_sub03_u_addr : 10'sh0 ) ;
	assign w_sub03_u_datain = ( (|r_sys_processing_methodID) ? r_sub03_u_datain : 32'h0 ) ;
	assign w_sub03_u_r_w = ( (|r_sys_processing_methodID) ? r_sub03_u_r_w : 1'h0 ) ;
	assign w_sub03_result_addr = ( (|r_sys_processing_methodID) ? r_sub03_result_addr : 10'sh0 ) ;
	assign w_sub03_result_datain = ( (|r_sys_processing_methodID) ? r_sub03_result_datain : 32'h0 ) ;
	assign w_sub03_result_r_w = ( (|r_sys_processing_methodID) ? r_sub03_result_r_w : 1'h0 ) ;
	assign w_sub02_u_addr = ( (|r_sys_processing_methodID) ? r_sub02_u_addr : 10'sh0 ) ;
	assign w_sub02_u_datain = ( (|r_sys_processing_methodID) ? r_sub02_u_datain : 32'h0 ) ;
	assign w_sub02_u_r_w = ( (|r_sys_processing_methodID) ? r_sub02_u_r_w : 1'h0 ) ;
	assign w_sub02_result_addr = ( (|r_sys_processing_methodID) ? r_sub02_result_addr : 10'sh0 ) ;
	assign w_sub02_result_datain = ( (|r_sys_processing_methodID) ? r_sub02_result_datain : 32'h0 ) ;
	assign w_sub02_result_r_w = ( (|r_sys_processing_methodID) ? r_sub02_result_r_w : 1'h0 ) ;
	assign w_sub01_u_addr = ( (|r_sys_processing_methodID) ? r_sub01_u_addr : 10'sh0 ) ;
	assign w_sub01_u_datain = ( (|r_sys_processing_methodID) ? r_sub01_u_datain : 32'h0 ) ;
	assign w_sub01_u_r_w = ( (|r_sys_processing_methodID) ? r_sub01_u_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 10'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub00_u_addr = ( (|r_sys_processing_methodID) ? r_sub00_u_addr : 10'sh0 ) ;
	assign w_sub00_u_datain = ( (|r_sys_processing_methodID) ? r_sub00_u_datain : 32'h0 ) ;
	assign w_sub00_u_r_w = ( (|r_sys_processing_methodID) ? r_sub00_u_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 10'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sub07_u_addr = ( (|r_sys_processing_methodID) ? r_sub07_u_addr : 10'sh0 ) ;
	assign w_sub07_u_datain = ( (|r_sys_processing_methodID) ? r_sub07_u_datain : 32'h0 ) ;
	assign w_sub07_u_r_w = ( (|r_sys_processing_methodID) ? r_sub07_u_r_w : 1'h0 ) ;
	assign w_sub07_result_addr = ( (|r_sys_processing_methodID) ? r_sub07_result_addr : 10'sh0 ) ;
	assign w_sub07_result_datain = ( (|r_sys_processing_methodID) ? r_sub07_result_datain : 32'h0 ) ;
	assign w_sub07_result_r_w = ( (|r_sys_processing_methodID) ? r_sub07_result_r_w : 1'h0 ) ;
	assign w_sub06_u_addr = ( (|r_sys_processing_methodID) ? r_sub06_u_addr : 10'sh0 ) ;
	assign w_sub06_u_datain = ( (|r_sys_processing_methodID) ? r_sub06_u_datain : 32'h0 ) ;
	assign w_sub06_u_r_w = ( (|r_sys_processing_methodID) ? r_sub06_u_r_w : 1'h0 ) ;
	assign w_sub06_result_addr = ( (|r_sys_processing_methodID) ? r_sub06_result_addr : 10'sh0 ) ;
	assign w_sub06_result_datain = ( (|r_sys_processing_methodID) ? r_sub06_result_datain : 32'h0 ) ;
	assign w_sub06_result_r_w = ( (|r_sys_processing_methodID) ? r_sub06_result_r_w : 1'h0 ) ;
	assign w_sub05_u_addr = ( (|r_sys_processing_methodID) ? r_sub05_u_addr : 10'sh0 ) ;
	assign w_sub05_u_datain = ( (|r_sys_processing_methodID) ? r_sub05_u_datain : 32'h0 ) ;
	assign w_sub05_u_r_w = ( (|r_sys_processing_methodID) ? r_sub05_u_r_w : 1'h0 ) ;
	assign w_sub05_result_addr = ( (|r_sys_processing_methodID) ? r_sub05_result_addr : 10'sh0 ) ;
	assign w_sub05_result_datain = ( (|r_sys_processing_methodID) ? r_sub05_result_datain : 32'h0 ) ;
	assign w_sub05_result_r_w = ( (|r_sys_processing_methodID) ? r_sub05_result_r_w : 1'h0 ) ;
	assign w_sub04_u_addr = ( (|r_sys_processing_methodID) ? r_sub04_u_addr : 10'sh0 ) ;
	assign w_sub04_u_datain = ( (|r_sys_processing_methodID) ? r_sub04_u_datain : 32'h0 ) ;
	assign w_sub04_u_r_w = ( (|r_sys_processing_methodID) ? r_sub04_u_r_w : 1'h0 ) ;
	assign w_sub04_result_addr = ( (|r_sys_processing_methodID) ? r_sub04_result_addr : 10'sh0 ) ;
	assign w_sub04_result_datain = ( (|r_sys_processing_methodID) ? r_sub04_result_datain : 32'h0 ) ;
	assign w_sub04_result_r_w = ( (|r_sys_processing_methodID) ? r_sub04_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh0000001f;
	assign w_sys_tmp3 = 32'sh00000002;
	assign w_sys_tmp4 = ( !w_sys_tmp5 );
	assign w_sys_tmp5 = (r_run_my_15 < r_run_k_11);
	assign w_sys_tmp6 = (r_run_k_11 + w_sys_intOne);
	assign w_sys_tmp7 = ( !w_sys_tmp8 );
	assign w_sys_tmp8 = (r_run_mx_14 < r_run_j_12);
	assign w_sys_tmp11 = (w_sys_tmp12 + r_run_k_11);
	assign w_sys_tmp12 = (r_run_j_12 * w_sys_tmp13);
	assign w_sys_tmp13 = 32'sh0000001f;
	assign w_sys_tmp14 = 32'h0;
	assign w_sys_tmp16 = (w_sys_tmp17 + r_run_k_11);
	assign w_sys_tmp17 = (r_run_copy0_j_17 * w_sys_tmp13);
	assign w_sys_tmp20 = (r_run_copy0_j_17 + w_sys_intOne);
	assign w_sys_tmp21 = (r_run_j_12 + w_sys_intOne);
	assign w_sys_tmp250 = ( !w_sys_tmp251 );
	assign w_sys_tmp251 = (r_run_nlast_16 < r_run_n_13);
	assign w_sys_tmp252 = (r_run_n_13 + w_sys_intOne);
	assign w_sys_tmp253 = ( !w_sys_tmp254 );
	assign w_sys_tmp254 = (r_run_my_15 < r_run_j_12);
	assign w_sys_tmp257 = (w_sys_tmp258 + r_run_j_12);
	assign w_sys_tmp258 = 32'sh0000001f;
	assign w_sys_tmp259 = 32'h3f000000;
	assign w_sys_tmp261 = (w_sys_tmp262 + r_run_copy2_j_20);
	assign w_sys_tmp262 = 32'sh000001b9;
	assign w_sys_tmp263 = 32'h0;
	assign w_sys_tmp265 = (w_sys_tmp266 + w_sys_intOne);
	assign w_sys_tmp266 = (r_run_copy1_j_19 * w_sys_tmp258);
	assign w_sys_tmp268 = 32'h3f800000;
	assign w_sys_tmp270 = (w_sys_tmp271 + r_run_my_15);
	assign w_sys_tmp271 = (r_run_copy0_j_18 * w_sys_tmp258);
	assign w_sys_tmp274 = (r_run_copy0_j_18 + w_sys_intOne);
	assign w_sys_tmp275 = (r_run_copy1_j_19 + w_sys_intOne);
	assign w_sys_tmp276 = (r_run_copy2_j_20 + w_sys_intOne);
	assign w_sys_tmp277 = (r_run_j_12 + w_sys_intOne);
	assign w_sys_tmp696 = ( !w_sys_tmp697 );
	assign w_sys_tmp697 = (w_sys_tmp698 < r_run_k_11);
	assign w_sys_tmp698 = 32'sh0000000c;
	assign w_sys_tmp701 = (w_sys_tmp702 + r_run_k_11);
	assign w_sys_tmp702 = 32'sh0000001f;
	assign w_sys_tmp703 = w_fld_u_0_dataout_1;
	assign w_sys_tmp707 = (w_sys_tmp708 + r_run_k_11);
	assign w_sys_tmp708 = 32'sh0000003e;
	assign w_sys_tmp713 = (w_sys_tmp714 + r_run_k_11);
	assign w_sys_tmp714 = 32'sh0000005d;
	assign w_sys_tmp719 = (w_sys_tmp720 + r_run_k_11);
	assign w_sys_tmp720 = 32'sh0000007c;
	assign w_sys_tmp725 = (w_sys_tmp726 + r_run_k_11);
	assign w_sys_tmp726 = 32'sh0000009b;
	assign w_sys_tmp731 = (w_sys_tmp732 + r_run_k_11);
	assign w_sys_tmp732 = 32'sh000000ba;
	assign w_sys_tmp737 = (w_sys_tmp738 + r_run_k_11);
	assign w_sys_tmp738 = 32'sh000000d9;
	assign w_sys_tmp743 = (w_sys_tmp744 + r_run_k_11);
	assign w_sys_tmp744 = 32'sh000000f8;
	assign w_sys_tmp749 = (w_sys_tmp750 + r_run_k_11);
	assign w_sys_tmp750 = 32'sh00000117;
	assign w_sys_tmp755 = (w_sys_tmp756 + r_run_k_11);
	assign w_sys_tmp756 = 32'sh00000136;
	assign w_sys_tmp761 = (w_sys_tmp762 + r_run_k_11);
	assign w_sys_tmp762 = 32'sh00000155;
	assign w_sys_tmp767 = (w_sys_tmp768 + r_run_k_11);
	assign w_sys_tmp768 = 32'sh00000174;
	assign w_sys_tmp785 = (w_sys_tmp786 + r_run_k_11);
	assign w_sys_tmp786 = 32'sh00000193;
	assign w_sys_tmp791 = (w_sys_tmp792 + r_run_k_11);
	assign w_sys_tmp792 = 32'sh000001b2;
	assign w_sys_tmp797 = (w_sys_tmp798 + r_run_k_11);
	assign w_sys_tmp798 = 32'sh000001d1;
	assign w_sys_tmp803 = (w_sys_tmp804 + r_run_k_11);
	assign w_sys_tmp804 = 32'sh000001f0;
	assign w_sys_tmp809 = (w_sys_tmp810 + r_run_k_11);
	assign w_sys_tmp810 = 32'sh0000020f;
	assign w_sys_tmp815 = (w_sys_tmp816 + r_run_k_11);
	assign w_sys_tmp816 = 32'sh0000022e;
	assign w_sys_tmp821 = (w_sys_tmp822 + r_run_k_11);
	assign w_sys_tmp822 = 32'sh0000024d;
	assign w_sys_tmp827 = (w_sys_tmp828 + r_run_k_11);
	assign w_sys_tmp828 = 32'sh0000026c;
	assign w_sys_tmp833 = (w_sys_tmp834 + r_run_k_11);
	assign w_sys_tmp834 = 32'sh0000028b;
	assign w_sys_tmp839 = (w_sys_tmp840 + r_run_k_11);
	assign w_sys_tmp840 = 32'sh000002aa;
	assign w_sys_tmp857 = (w_sys_tmp858 + r_run_k_11);
	assign w_sys_tmp858 = 32'sh000002c9;
	assign w_sys_tmp863 = (w_sys_tmp864 + r_run_k_11);
	assign w_sys_tmp864 = 32'sh000002e8;
	assign w_sys_tmp869 = (w_sys_tmp870 + r_run_k_11);
	assign w_sys_tmp870 = 32'sh00000307;
	assign w_sys_tmp875 = (w_sys_tmp876 + r_run_k_11);
	assign w_sys_tmp876 = 32'sh00000326;
	assign w_sys_tmp881 = (w_sys_tmp882 + r_run_k_11);
	assign w_sys_tmp882 = 32'sh00000345;
	assign w_sys_tmp887 = (w_sys_tmp888 + r_run_k_11);
	assign w_sys_tmp888 = 32'sh00000364;
	assign w_sys_tmp893 = (w_sys_tmp894 + r_run_k_11);
	assign w_sys_tmp894 = 32'sh00000383;
	assign w_sys_tmp899 = (w_sys_tmp900 + r_run_k_11);
	assign w_sys_tmp900 = 32'sh000003a2;
	assign w_sys_tmp905 = (w_sys_tmp906 + r_run_k_11);
	assign w_sys_tmp906 = 32'sh000003c1;
	assign w_sys_tmp911 = (w_sys_tmp912 + r_run_k_11);
	assign w_sys_tmp912 = 32'sh00000029;
	assign w_sys_tmp917 = (w_sys_tmp918 + r_run_k_11);
	assign w_sys_tmp918 = 32'sh00000048;
	assign w_sys_tmp923 = (w_sys_tmp924 + r_run_k_11);
	assign w_sys_tmp924 = 32'sh00000067;
	assign w_sys_tmp929 = (w_sys_tmp930 + r_run_k_11);
	assign w_sys_tmp930 = 32'sh00000086;
	assign w_sys_tmp935 = (w_sys_tmp936 + r_run_k_11);
	assign w_sys_tmp936 = 32'sh000000a5;
	assign w_sys_tmp941 = (w_sys_tmp942 + r_run_k_11);
	assign w_sys_tmp942 = 32'sh000000c4;
	assign w_sys_tmp947 = (w_sys_tmp948 + r_run_k_11);
	assign w_sys_tmp948 = 32'sh000000e3;
	assign w_sys_tmp953 = (w_sys_tmp954 + r_run_k_11);
	assign w_sys_tmp954 = 32'sh00000102;
	assign w_sys_tmp959 = (w_sys_tmp960 + r_run_k_11);
	assign w_sys_tmp960 = 32'sh00000121;
	assign w_sys_tmp965 = (w_sys_tmp966 + r_run_k_11);
	assign w_sys_tmp966 = 32'sh00000140;
	assign w_sys_tmp971 = (w_sys_tmp972 + r_run_k_11);
	assign w_sys_tmp972 = 32'sh0000015f;
	assign w_sys_tmp977 = (w_sys_tmp978 + r_run_k_11);
	assign w_sys_tmp978 = 32'sh0000017e;
	assign w_sys_tmp995 = (w_sys_tmp996 + r_run_k_11);
	assign w_sys_tmp996 = 32'sh0000019d;
	assign w_sys_tmp1001 = (w_sys_tmp1002 + r_run_k_11);
	assign w_sys_tmp1002 = 32'sh000001bc;
	assign w_sys_tmp1007 = (w_sys_tmp1008 + r_run_k_11);
	assign w_sys_tmp1008 = 32'sh000001db;
	assign w_sys_tmp1013 = (w_sys_tmp1014 + r_run_k_11);
	assign w_sys_tmp1014 = 32'sh000001fa;
	assign w_sys_tmp1019 = (w_sys_tmp1020 + r_run_k_11);
	assign w_sys_tmp1020 = 32'sh00000219;
	assign w_sys_tmp1025 = (w_sys_tmp1026 + r_run_k_11);
	assign w_sys_tmp1026 = 32'sh00000238;
	assign w_sys_tmp1031 = (w_sys_tmp1032 + r_run_k_11);
	assign w_sys_tmp1032 = 32'sh00000257;
	assign w_sys_tmp1037 = (w_sys_tmp1038 + r_run_k_11);
	assign w_sys_tmp1038 = 32'sh00000276;
	assign w_sys_tmp1043 = (w_sys_tmp1044 + r_run_k_11);
	assign w_sys_tmp1044 = 32'sh00000295;
	assign w_sys_tmp1049 = (w_sys_tmp1050 + r_run_k_11);
	assign w_sys_tmp1050 = 32'sh000002b4;
	assign w_sys_tmp1067 = (w_sys_tmp1068 + r_run_k_11);
	assign w_sys_tmp1068 = 32'sh000002d3;
	assign w_sys_tmp1073 = (w_sys_tmp1074 + r_run_k_11);
	assign w_sys_tmp1074 = 32'sh000002f2;
	assign w_sys_tmp1079 = (w_sys_tmp1080 + r_run_k_11);
	assign w_sys_tmp1080 = 32'sh00000311;
	assign w_sys_tmp1085 = (w_sys_tmp1086 + r_run_k_11);
	assign w_sys_tmp1086 = 32'sh00000330;
	assign w_sys_tmp1091 = (w_sys_tmp1092 + r_run_k_11);
	assign w_sys_tmp1092 = 32'sh0000034f;
	assign w_sys_tmp1097 = (w_sys_tmp1098 + r_run_k_11);
	assign w_sys_tmp1098 = 32'sh0000036e;
	assign w_sys_tmp1103 = (w_sys_tmp1104 + r_run_k_11);
	assign w_sys_tmp1104 = 32'sh0000038d;
	assign w_sys_tmp1109 = (w_sys_tmp1110 + r_run_k_11);
	assign w_sys_tmp1110 = 32'sh000003ac;
	assign w_sys_tmp1115 = (w_sys_tmp1116 + r_run_k_11);
	assign w_sys_tmp1116 = 32'sh000003cb;
	assign w_sys_tmp1120 = (r_run_k_11 + w_sys_intOne);
	assign w_sys_tmp1121 = 32'sh00000015;
	assign w_sys_tmp1122 = ( !w_sys_tmp1123 );
	assign w_sys_tmp1123 = (w_sys_tmp1124 < r_run_k_11);
	assign w_sys_tmp1124 = 32'sh0000001f;
	assign w_sys_tmp1127 = (w_sys_tmp1128 + r_run_k_11);
	assign w_sys_tmp1128 = 32'sh0000001f;
	assign w_sys_tmp1129 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1133 = (w_sys_tmp1134 + r_run_k_11);
	assign w_sys_tmp1134 = 32'sh0000003e;
	assign w_sys_tmp1139 = (w_sys_tmp1140 + r_run_k_11);
	assign w_sys_tmp1140 = 32'sh0000005d;
	assign w_sys_tmp1145 = (w_sys_tmp1146 + r_run_k_11);
	assign w_sys_tmp1146 = 32'sh0000007c;
	assign w_sys_tmp1151 = (w_sys_tmp1152 + r_run_k_11);
	assign w_sys_tmp1152 = 32'sh0000009b;
	assign w_sys_tmp1157 = (w_sys_tmp1158 + r_run_k_11);
	assign w_sys_tmp1158 = 32'sh000000ba;
	assign w_sys_tmp1163 = (w_sys_tmp1164 + r_run_k_11);
	assign w_sys_tmp1164 = 32'sh000000d9;
	assign w_sys_tmp1169 = (w_sys_tmp1170 + r_run_k_11);
	assign w_sys_tmp1170 = 32'sh000000f8;
	assign w_sys_tmp1175 = (w_sys_tmp1176 + r_run_k_11);
	assign w_sys_tmp1176 = 32'sh00000117;
	assign w_sys_tmp1181 = (w_sys_tmp1182 + r_run_k_11);
	assign w_sys_tmp1182 = 32'sh00000136;
	assign w_sys_tmp1187 = (w_sys_tmp1188 + r_run_k_11);
	assign w_sys_tmp1188 = 32'sh00000155;
	assign w_sys_tmp1193 = (w_sys_tmp1194 + r_run_k_11);
	assign w_sys_tmp1194 = 32'sh00000174;
	assign w_sys_tmp1211 = (w_sys_tmp1212 + r_run_k_11);
	assign w_sys_tmp1212 = 32'sh00000193;
	assign w_sys_tmp1217 = (w_sys_tmp1218 + r_run_k_11);
	assign w_sys_tmp1218 = 32'sh000001b2;
	assign w_sys_tmp1223 = (w_sys_tmp1224 + r_run_k_11);
	assign w_sys_tmp1224 = 32'sh000001d1;
	assign w_sys_tmp1229 = (w_sys_tmp1230 + r_run_k_11);
	assign w_sys_tmp1230 = 32'sh000001f0;
	assign w_sys_tmp1235 = (w_sys_tmp1236 + r_run_k_11);
	assign w_sys_tmp1236 = 32'sh0000020f;
	assign w_sys_tmp1241 = (w_sys_tmp1242 + r_run_k_11);
	assign w_sys_tmp1242 = 32'sh0000022e;
	assign w_sys_tmp1247 = (w_sys_tmp1248 + r_run_k_11);
	assign w_sys_tmp1248 = 32'sh0000024d;
	assign w_sys_tmp1253 = (w_sys_tmp1254 + r_run_k_11);
	assign w_sys_tmp1254 = 32'sh0000026c;
	assign w_sys_tmp1259 = (w_sys_tmp1260 + r_run_k_11);
	assign w_sys_tmp1260 = 32'sh0000028b;
	assign w_sys_tmp1271 = (w_sys_tmp1272 + r_run_k_11);
	assign w_sys_tmp1272 = 32'sh000002aa;
	assign w_sys_tmp1277 = (w_sys_tmp1278 + r_run_k_11);
	assign w_sys_tmp1278 = 32'sh000002c9;
	assign w_sys_tmp1283 = (w_sys_tmp1284 + r_run_k_11);
	assign w_sys_tmp1284 = 32'sh000002e8;
	assign w_sys_tmp1289 = (w_sys_tmp1290 + r_run_k_11);
	assign w_sys_tmp1290 = 32'sh00000307;
	assign w_sys_tmp1295 = (w_sys_tmp1296 + r_run_k_11);
	assign w_sys_tmp1296 = 32'sh00000326;
	assign w_sys_tmp1301 = (w_sys_tmp1302 + r_run_k_11);
	assign w_sys_tmp1302 = 32'sh00000345;
	assign w_sys_tmp1307 = (w_sys_tmp1308 + r_run_k_11);
	assign w_sys_tmp1308 = 32'sh00000364;
	assign w_sys_tmp1313 = (w_sys_tmp1314 + r_run_k_11);
	assign w_sys_tmp1314 = 32'sh00000383;
	assign w_sys_tmp1319 = (w_sys_tmp1320 + r_run_k_11);
	assign w_sys_tmp1320 = 32'sh000003a2;
	assign w_sys_tmp1324 = (r_run_k_11 + w_sys_intOne);
	assign w_sys_tmp1325 = 32'sh00000002;
	assign w_sys_tmp1326 = ( !w_sys_tmp1327 );
	assign w_sys_tmp1327 = (w_sys_tmp1328 < r_run_k_11);
	assign w_sys_tmp1328 = 32'sh0000000b;
	assign w_sys_tmp1331 = (w_sys_tmp1332 + r_run_k_11);
	assign w_sys_tmp1332 = 32'sh0000003e;
	assign w_sys_tmp1333 = w_sub00_result_dataout;
	assign w_sys_tmp1337 = (w_sys_tmp1338 + r_run_k_11);
	assign w_sys_tmp1338 = 32'sh0000005d;
	assign w_sys_tmp1343 = (w_sys_tmp1344 + r_run_k_11);
	assign w_sys_tmp1344 = 32'sh0000007c;
	assign w_sys_tmp1349 = (w_sys_tmp1350 + r_run_k_11);
	assign w_sys_tmp1350 = 32'sh0000009b;
	assign w_sys_tmp1355 = (w_sys_tmp1356 + r_run_k_11);
	assign w_sys_tmp1356 = 32'sh000000ba;
	assign w_sys_tmp1361 = (w_sys_tmp1362 + r_run_k_11);
	assign w_sys_tmp1362 = 32'sh000000d9;
	assign w_sys_tmp1367 = (w_sys_tmp1368 + r_run_k_11);
	assign w_sys_tmp1368 = 32'sh000000f8;
	assign w_sys_tmp1373 = (w_sys_tmp1374 + r_run_k_11);
	assign w_sys_tmp1374 = 32'sh00000117;
	assign w_sys_tmp1379 = (w_sys_tmp1380 + r_run_k_11);
	assign w_sys_tmp1380 = 32'sh00000136;
	assign w_sys_tmp1385 = (w_sys_tmp1386 + r_run_k_11);
	assign w_sys_tmp1386 = 32'sh00000155;
	assign w_sys_tmp1391 = (w_sys_tmp1392 + r_run_k_11);
	assign w_sys_tmp1392 = 32'sh00000174;
	assign w_sys_tmp1396 = (w_sys_tmp1397 + r_run_k_11);
	assign w_sys_tmp1397 = 32'sh00000193;
	assign w_sys_tmp1401 = (w_sys_tmp1402 + r_run_k_11);
	assign w_sys_tmp1402 = 32'sh000001b2;
	assign w_sys_tmp1406 = (w_sys_tmp1407 + r_run_k_11);
	assign w_sys_tmp1407 = 32'sh000001d1;
	assign w_sys_tmp1411 = (w_sys_tmp1412 + r_run_k_11);
	assign w_sys_tmp1412 = 32'sh000001f0;
	assign w_sys_tmp1416 = (w_sys_tmp1417 + r_run_k_11);
	assign w_sys_tmp1417 = 32'sh0000020f;
	assign w_sys_tmp1421 = (w_sys_tmp1422 + r_run_k_11);
	assign w_sys_tmp1422 = 32'sh0000022e;
	assign w_sys_tmp1426 = (w_sys_tmp1427 + r_run_k_11);
	assign w_sys_tmp1427 = 32'sh0000024d;
	assign w_sys_tmp1431 = (w_sys_tmp1432 + r_run_k_11);
	assign w_sys_tmp1432 = 32'sh0000026c;
	assign w_sys_tmp1436 = (w_sys_tmp1437 + r_run_k_11);
	assign w_sys_tmp1437 = 32'sh0000028b;
	assign w_sys_tmp1441 = (w_sys_tmp1442 + r_run_k_11);
	assign w_sys_tmp1442 = 32'sh000002aa;
	assign w_sys_tmp1446 = (w_sys_tmp1447 + r_run_k_11);
	assign w_sys_tmp1447 = 32'sh000002c9;
	assign w_sys_tmp1451 = (w_sys_tmp1452 + r_run_k_11);
	assign w_sys_tmp1452 = 32'sh000002e8;
	assign w_sys_tmp1456 = (w_sys_tmp1457 + r_run_k_11);
	assign w_sys_tmp1457 = 32'sh00000307;
	assign w_sys_tmp1461 = (w_sys_tmp1462 + r_run_k_11);
	assign w_sys_tmp1462 = 32'sh00000326;
	assign w_sys_tmp1466 = (w_sys_tmp1467 + r_run_k_11);
	assign w_sys_tmp1467 = 32'sh00000345;
	assign w_sys_tmp1471 = (w_sys_tmp1472 + r_run_k_11);
	assign w_sys_tmp1472 = 32'sh00000364;
	assign w_sys_tmp1476 = (w_sys_tmp1477 + r_run_k_11);
	assign w_sys_tmp1477 = 32'sh00000383;
	assign w_sys_tmp1481 = (w_sys_tmp1482 + r_run_k_11);
	assign w_sys_tmp1482 = 32'sh000003a2;
	assign w_sys_tmp1486 = (w_sys_tmp1487 + r_run_k_11);
	assign w_sys_tmp1487 = 32'sh00000048;
	assign w_sys_tmp1491 = (w_sys_tmp1492 + r_run_k_11);
	assign w_sys_tmp1492 = 32'sh00000067;
	assign w_sys_tmp1496 = (w_sys_tmp1497 + r_run_k_11);
	assign w_sys_tmp1497 = 32'sh00000086;
	assign w_sys_tmp1501 = (w_sys_tmp1502 + r_run_k_11);
	assign w_sys_tmp1502 = 32'sh000000a5;
	assign w_sys_tmp1506 = (w_sys_tmp1507 + r_run_k_11);
	assign w_sys_tmp1507 = 32'sh000000c4;
	assign w_sys_tmp1511 = (w_sys_tmp1512 + r_run_k_11);
	assign w_sys_tmp1512 = 32'sh000000e3;
	assign w_sys_tmp1516 = (w_sys_tmp1517 + r_run_k_11);
	assign w_sys_tmp1517 = 32'sh00000102;
	assign w_sys_tmp1521 = (w_sys_tmp1522 + r_run_k_11);
	assign w_sys_tmp1522 = 32'sh00000121;
	assign w_sys_tmp1526 = (w_sys_tmp1527 + r_run_k_11);
	assign w_sys_tmp1527 = 32'sh00000140;
	assign w_sys_tmp1531 = (w_sys_tmp1532 + r_run_k_11);
	assign w_sys_tmp1532 = 32'sh0000015f;
	assign w_sys_tmp1536 = (w_sys_tmp1537 + r_run_k_11);
	assign w_sys_tmp1537 = 32'sh0000017e;
	assign w_sys_tmp1541 = (w_sys_tmp1542 + r_run_k_11);
	assign w_sys_tmp1542 = 32'sh0000019d;
	assign w_sys_tmp1546 = (w_sys_tmp1547 + r_run_k_11);
	assign w_sys_tmp1547 = 32'sh000001bc;
	assign w_sys_tmp1551 = (w_sys_tmp1552 + r_run_k_11);
	assign w_sys_tmp1552 = 32'sh000001db;
	assign w_sys_tmp1556 = (w_sys_tmp1557 + r_run_k_11);
	assign w_sys_tmp1557 = 32'sh000001fa;
	assign w_sys_tmp1561 = (w_sys_tmp1562 + r_run_k_11);
	assign w_sys_tmp1562 = 32'sh00000219;
	assign w_sys_tmp1566 = (w_sys_tmp1567 + r_run_k_11);
	assign w_sys_tmp1567 = 32'sh00000238;
	assign w_sys_tmp1571 = (w_sys_tmp1572 + r_run_k_11);
	assign w_sys_tmp1572 = 32'sh00000257;
	assign w_sys_tmp1576 = (w_sys_tmp1577 + r_run_k_11);
	assign w_sys_tmp1577 = 32'sh00000276;
	assign w_sys_tmp1581 = (w_sys_tmp1582 + r_run_k_11);
	assign w_sys_tmp1582 = 32'sh00000295;
	assign w_sys_tmp1586 = (w_sys_tmp1587 + r_run_k_11);
	assign w_sys_tmp1587 = 32'sh000002b4;
	assign w_sys_tmp1591 = (w_sys_tmp1592 + r_run_k_11);
	assign w_sys_tmp1592 = 32'sh000002d3;
	assign w_sys_tmp1596 = (w_sys_tmp1597 + r_run_k_11);
	assign w_sys_tmp1597 = 32'sh000002f2;
	assign w_sys_tmp1601 = (w_sys_tmp1602 + r_run_k_11);
	assign w_sys_tmp1602 = 32'sh00000311;
	assign w_sys_tmp1606 = (w_sys_tmp1607 + r_run_k_11);
	assign w_sys_tmp1607 = 32'sh00000330;
	assign w_sys_tmp1611 = (w_sys_tmp1612 + r_run_k_11);
	assign w_sys_tmp1612 = 32'sh0000034f;
	assign w_sys_tmp1616 = (w_sys_tmp1617 + r_run_k_11);
	assign w_sys_tmp1617 = 32'sh0000036e;
	assign w_sys_tmp1621 = (w_sys_tmp1622 + r_run_k_11);
	assign w_sys_tmp1622 = 32'sh0000038d;
	assign w_sys_tmp1626 = (w_sys_tmp1627 + r_run_k_11);
	assign w_sys_tmp1627 = 32'sh000003ac;
	assign w_sys_tmp1630 = (r_run_k_11 + w_sys_intOne);
	assign w_sys_tmp1631 = 32'sh00000016;
	assign w_sys_tmp1632 = ( !w_sys_tmp1633 );
	assign w_sys_tmp1633 = (w_sys_tmp1634 < r_run_k_11);
	assign w_sys_tmp1634 = 32'sh0000001e;
	assign w_sys_tmp1637 = (w_sys_tmp1638 + r_run_k_11);
	assign w_sys_tmp1638 = 32'sh0000003e;
	assign w_sys_tmp1639 = w_sub06_result_dataout;
	assign w_sys_tmp1643 = (w_sys_tmp1644 + r_run_k_11);
	assign w_sys_tmp1644 = 32'sh0000005d;
	assign w_sys_tmp1649 = (w_sys_tmp1650 + r_run_k_11);
	assign w_sys_tmp1650 = 32'sh0000007c;
	assign w_sys_tmp1655 = (w_sys_tmp1656 + r_run_k_11);
	assign w_sys_tmp1656 = 32'sh0000009b;
	assign w_sys_tmp1661 = (w_sys_tmp1662 + r_run_k_11);
	assign w_sys_tmp1662 = 32'sh000000ba;
	assign w_sys_tmp1667 = (w_sys_tmp1668 + r_run_k_11);
	assign w_sys_tmp1668 = 32'sh000000d9;
	assign w_sys_tmp1673 = (w_sys_tmp1674 + r_run_k_11);
	assign w_sys_tmp1674 = 32'sh000000f8;
	assign w_sys_tmp1679 = (w_sys_tmp1680 + r_run_k_11);
	assign w_sys_tmp1680 = 32'sh00000117;
	assign w_sys_tmp1685 = (w_sys_tmp1686 + r_run_k_11);
	assign w_sys_tmp1686 = 32'sh00000136;
	assign w_sys_tmp1691 = (w_sys_tmp1692 + r_run_k_11);
	assign w_sys_tmp1692 = 32'sh00000155;
	assign w_sys_tmp1697 = (w_sys_tmp1698 + r_run_k_11);
	assign w_sys_tmp1698 = 32'sh00000174;
	assign w_sys_tmp1702 = (w_sys_tmp1703 + r_run_k_11);
	assign w_sys_tmp1703 = 32'sh00000193;
	assign w_sys_tmp1707 = (w_sys_tmp1708 + r_run_k_11);
	assign w_sys_tmp1708 = 32'sh000001b2;
	assign w_sys_tmp1712 = (w_sys_tmp1713 + r_run_k_11);
	assign w_sys_tmp1713 = 32'sh000001d1;
	assign w_sys_tmp1717 = (w_sys_tmp1718 + r_run_k_11);
	assign w_sys_tmp1718 = 32'sh000001f0;
	assign w_sys_tmp1722 = (w_sys_tmp1723 + r_run_k_11);
	assign w_sys_tmp1723 = 32'sh0000020f;
	assign w_sys_tmp1727 = (w_sys_tmp1728 + r_run_k_11);
	assign w_sys_tmp1728 = 32'sh0000022e;
	assign w_sys_tmp1732 = (w_sys_tmp1733 + r_run_k_11);
	assign w_sys_tmp1733 = 32'sh0000024d;
	assign w_sys_tmp1737 = (w_sys_tmp1738 + r_run_k_11);
	assign w_sys_tmp1738 = 32'sh0000026c;
	assign w_sys_tmp1742 = (w_sys_tmp1743 + r_run_k_11);
	assign w_sys_tmp1743 = 32'sh0000028b;
	assign w_sys_tmp1747 = (w_sys_tmp1748 + r_run_k_11);
	assign w_sys_tmp1748 = 32'sh000002aa;
	assign w_sys_tmp1757 = (w_sys_tmp1758 + r_run_k_11);
	assign w_sys_tmp1758 = 32'sh000002c9;
	assign w_sys_tmp1762 = (w_sys_tmp1763 + r_run_k_11);
	assign w_sys_tmp1763 = 32'sh000002e8;
	assign w_sys_tmp1767 = (w_sys_tmp1768 + r_run_k_11);
	assign w_sys_tmp1768 = 32'sh00000307;
	assign w_sys_tmp1772 = (w_sys_tmp1773 + r_run_k_11);
	assign w_sys_tmp1773 = 32'sh00000326;
	assign w_sys_tmp1777 = (w_sys_tmp1778 + r_run_k_11);
	assign w_sys_tmp1778 = 32'sh00000345;
	assign w_sys_tmp1782 = (w_sys_tmp1783 + r_run_k_11);
	assign w_sys_tmp1783 = 32'sh00000364;
	assign w_sys_tmp1787 = (w_sys_tmp1788 + r_run_k_11);
	assign w_sys_tmp1788 = 32'sh00000383;
	assign w_sys_tmp1792 = (w_sys_tmp1793 + r_run_k_11);
	assign w_sys_tmp1793 = 32'sh000003a2;
	assign w_sys_tmp1796 = (r_run_k_11 + w_sys_intOne);


	sub08
		sub08_inst(
			.i_fld_result_1_addr_0 (w_sub08_result_addr),
			.i_fld_result_1_datain_0 (w_sub08_result_datain),
			.o_fld_result_1_dataout_0 (w_sub08_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub08_result_r_w),
			.i_fld_u_0_addr_0 (w_sub08_u_addr),
			.i_fld_u_0_datain_0 (w_sub08_u_datain),
			.o_fld_u_0_dataout_0 (w_sub08_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub08_u_r_w),
			.o_run_busy (w_sub08_run_busy),
			.i_run_req (r_sub08_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub03
		sub03_inst(
			.i_fld_result_1_addr_0 (w_sub03_result_addr),
			.i_fld_result_1_datain_0 (w_sub03_result_datain),
			.o_fld_result_1_dataout_0 (w_sub03_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub03_result_r_w),
			.i_fld_u_0_addr_0 (w_sub03_u_addr),
			.i_fld_u_0_datain_0 (w_sub03_u_datain),
			.o_fld_u_0_dataout_0 (w_sub03_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub03_u_r_w),
			.o_run_busy (w_sub03_run_busy),
			.i_run_req (r_sub03_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub02
		sub02_inst(
			.i_fld_result_1_addr_0 (w_sub02_result_addr),
			.i_fld_result_1_datain_0 (w_sub02_result_datain),
			.o_fld_result_1_dataout_0 (w_sub02_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub02_result_r_w),
			.i_fld_u_0_addr_0 (w_sub02_u_addr),
			.i_fld_u_0_datain_0 (w_sub02_u_datain),
			.o_fld_u_0_dataout_0 (w_sub02_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub02_u_r_w),
			.o_run_busy (w_sub02_run_busy),
			.i_run_req (r_sub02_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub01
		sub01_inst(
			.i_fld_result_1_addr_0 (w_sub01_result_addr),
			.i_fld_result_1_datain_0 (w_sub01_result_datain),
			.o_fld_result_1_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub01_result_r_w),
			.i_fld_u_0_addr_0 (w_sub01_u_addr),
			.i_fld_u_0_datain_0 (w_sub01_u_datain),
			.o_fld_u_0_dataout_0 (w_sub01_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub01_u_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub00
		sub00_inst(
			.i_fld_result_1_addr_0 (w_sub00_result_addr),
			.i_fld_result_1_datain_0 (w_sub00_result_datain),
			.o_fld_result_1_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub00_result_r_w),
			.i_fld_u_0_addr_0 (w_sub00_u_addr),
			.i_fld_u_0_datain_0 (w_sub00_u_datain),
			.o_fld_u_0_dataout_0 (w_sub00_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub00_u_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub07
		sub07_inst(
			.i_fld_result_1_addr_0 (w_sub07_result_addr),
			.i_fld_result_1_datain_0 (w_sub07_result_datain),
			.o_fld_result_1_dataout_0 (w_sub07_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub07_result_r_w),
			.i_fld_u_0_addr_0 (w_sub07_u_addr),
			.i_fld_u_0_datain_0 (w_sub07_u_datain),
			.o_fld_u_0_dataout_0 (w_sub07_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub07_u_r_w),
			.o_run_busy (w_sub07_run_busy),
			.i_run_req (r_sub07_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub06
		sub06_inst(
			.i_fld_result_1_addr_0 (w_sub06_result_addr),
			.i_fld_result_1_datain_0 (w_sub06_result_datain),
			.o_fld_result_1_dataout_0 (w_sub06_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub06_result_r_w),
			.i_fld_u_0_addr_0 (w_sub06_u_addr),
			.i_fld_u_0_datain_0 (w_sub06_u_datain),
			.o_fld_u_0_dataout_0 (w_sub06_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub06_u_r_w),
			.o_run_busy (w_sub06_run_busy),
			.i_run_req (r_sub06_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub05
		sub05_inst(
			.i_fld_result_1_addr_0 (w_sub05_result_addr),
			.i_fld_result_1_datain_0 (w_sub05_result_datain),
			.o_fld_result_1_dataout_0 (w_sub05_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub05_result_r_w),
			.i_fld_u_0_addr_0 (w_sub05_u_addr),
			.i_fld_u_0_datain_0 (w_sub05_u_datain),
			.o_fld_u_0_dataout_0 (w_sub05_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub05_u_r_w),
			.o_run_busy (w_sub05_run_busy),
			.i_run_req (r_sub05_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub04
		sub04_inst(
			.i_fld_result_1_addr_0 (w_sub04_result_addr),
			.i_fld_result_1_datain_0 (w_sub04_result_datain),
			.o_fld_result_1_dataout_0 (w_sub04_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub04_result_r_w),
			.i_fld_u_0_addr_0 (w_sub04_u_addr),
			.i_fld_u_0_datain_0 (w_sub04_u_datain),
			.o_fld_u_0_dataout_0 (w_sub04_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub04_u_r_w),
			.o_run_busy (w_sub04_run_busy),
			.i_run_req (r_sub04_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(9), .WORDS(484) )
		dpram_u_0(
			.clk (clock),
			.ce_0 (w_fld_u_0_ce_0),
			.addr_0 (w_fld_u_0_addr_0),
			.datain_0 (w_fld_u_0_datain_0),
			.dataout_0 (w_fld_u_0_dataout_0),
			.r_w_0 (w_fld_u_0_r_w_0),
			.ce_1 (w_fld_u_0_ce_1),
			.addr_1 (r_fld_u_0_addr_1),
			.datain_1 (r_fld_u_0_datain_1),
			.dataout_1 (w_fld_u_0_dataout_1),
			.r_w_1 (r_fld_u_0_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(9), .WORDS(484) )
		dpram_uu_1(
			.clk (clock),
			.ce_0 (w_fld_uu_1_ce_0),
			.addr_0 (w_fld_uu_1_addr_0),
			.datain_0 (w_fld_uu_1_datain_0),
			.dataout_0 (w_fld_uu_1_dataout_0),
			.r_w_0 (w_fld_uu_1_r_w_0),
			.ce_1 (w_fld_uu_1_ce_1),
			.addr_1 (r_fld_uu_1_addr_1),
			.datain_1 (r_fld_uu_1_datain_1),
			.dataout_1 (w_fld_uu_1_dataout_1),
			.r_w_1 (r_fld_uu_1_r_w_1)
		);

	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h35: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 6'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_phase <= 6'h2;
						end

						6'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h4;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4) ? 6'h9 : 6'hf);

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'ha;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7) ? 6'hd : 6'h6);

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h13)) begin
										r_sys_run_phase <= 6'ha;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h10;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp250) ? 6'h14 : 6'h35);

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h10;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h15;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp253) ? 6'h18 : 6'h1a);

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4f)) begin
										r_sys_run_phase <= 6'h15;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h1b;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp696) ? 6'h1e : 6'h20);

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h47)) begin
										r_sys_run_phase <= 6'h1b;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h21;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1122) ? 6'h24 : 6'h25);

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h22)) begin
										r_sys_run_phase <= 6'h21;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_phase <= 6'h27;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								4'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_phase <= 6'h29;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h2a;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1326) ? 6'h2d : 6'h2f);

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3b)) begin
										r_sys_run_phase <= 6'h2a;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h30;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1632) ? 6'h33 : 6'h11);

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1f)) begin
										r_sys_run_phase <= 6'h30;

									end
								end

							endcase
						end

						6'h35: begin
							r_sys_run_phase <= 6'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 4'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h13)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4f)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h47)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h22)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3b)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1f)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 7'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h13)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h12)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4f)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h4e)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h47)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h46)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h22)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h21)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub00_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub01_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub02_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub03_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub04_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub05_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub06_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub07_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub08_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3b)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3a)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1f)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h1e)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						6'h35: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_addr_1 <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp11[8:0] );

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1) || (r_sys_run_step==7'h5) || (r_sys_run_step==7'h9) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h45) || (r_sys_run_step==7'h49) || (r_sys_run_step==7'h4d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp261[8:0] );

									end
									else
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h3e) || (r_sys_run_step==7'h42) || (r_sys_run_step==7'h46) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h4e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp265[8:0] );

									end
									else
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h2b) || (r_sys_run_step==7'h2f) || (r_sys_run_step==7'h33) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h3b) || (r_sys_run_step==7'h3f) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h47) || (r_sys_run_step==7'h4b) || (r_sys_run_step==7'h4f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp270[8:0] );

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h4) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h38) || (r_sys_run_step==7'h3c) || (r_sys_run_step==7'h40) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h48) || (r_sys_run_step==7'h4c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp257[8:0] );

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h38)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1037[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp743[8:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp875[8:0] );

									end
									else
									if((r_sys_run_step==7'h39) || (r_sys_run_step==7'h3b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1043[8:0] );

									end
									else
									if((r_sys_run_step==7'h22)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp905[8:0] );

									end
									else
									if((r_sys_run_step==7'h2b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp959[8:0] );

									end
									else
									if((r_sys_run_step==7'h17) || (r_sys_run_step==7'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp839[8:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp869[8:0] );

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1019[8:0] );

									end
									else
									if((r_sys_run_step==7'h3f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1079[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp731[8:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp893[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp749[8:0] );

									end
									else
									if((r_sys_run_step==7'h27)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp935[8:0] );

									end
									else
									if((r_sys_run_step==7'h29)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp947[8:0] );

									end
									else
									if((r_sys_run_step==7'h24)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp917[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp719[8:0] );

									end
									else
									if((r_sys_run_step==7'h3d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1067[8:0] );

									end
									else
									if((r_sys_run_step==7'h34)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1013[8:0] );

									end
									else
									if((r_sys_run_step==7'h41)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1091[8:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp881[8:0] );

									end
									else
									if((r_sys_run_step==7'h2d) || (r_sys_run_step==7'h2f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp971[8:0] );

									end
									else
									if((r_sys_run_step==7'h16) || (r_sys_run_step==7'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp833[8:0] );

									end
									else
									if((r_sys_run_step==7'hb) || (r_sys_run_step==7'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp767[8:0] );

									end
									else
									if((r_sys_run_step==7'h32)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1001[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp815[8:0] );

									end
									else
									if((r_sys_run_step==7'h45)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1115[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp701[8:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp887[8:0] );

									end
									else
									if((r_sys_run_step==7'h44)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1109[8:0] );

									end
									else
									if((r_sys_run_step==7'h36)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1025[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp857[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp803[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp725[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp863[8:0] );

									end
									else
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp761[8:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp827[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp737[8:0] );

									end
									else
									if((r_sys_run_step==7'h37)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1031[8:0] );

									end
									else
									if((r_sys_run_step==7'h23)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp911[8:0] );

									end
									else
									if((r_sys_run_step==7'h25)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp923[8:0] );

									end
									else
									if((r_sys_run_step==7'h31)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp995[8:0] );

									end
									else
									if((r_sys_run_step==7'h42)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1097[8:0] );

									end
									else
									if((r_sys_run_step==7'h40)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1085[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp809[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp707[8:0] );

									end
									else
									if((r_sys_run_step==7'h2a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp953[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp785[8:0] );

									end
									else
									if((r_sys_run_step==7'h2e) || (r_sys_run_step==7'h30)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp977[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp755[8:0] );

									end
									else
									if((r_sys_run_step==7'h26)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp929[8:0] );

									end
									else
									if((r_sys_run_step==7'h33)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1007[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp791[8:0] );

									end
									else
									if((r_sys_run_step==7'h3a) || (r_sys_run_step==7'h3c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1049[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp821[8:0] );

									end
									else
									if((r_sys_run_step==7'h43)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1103[8:0] );

									end
									else
									if((r_sys_run_step==7'h28)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp941[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp713[8:0] );

									end
									else
									if((r_sys_run_step==7'h3e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1073[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp797[8:0] );

									end
									else
									if((r_sys_run_step==7'h2c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp965[8:0] );

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp899[8:0] );

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1229[8:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1253[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1235[8:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1301[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1175[8:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1313[8:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1295[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1127[8:0] );

									end
									else
									if((r_sys_run_step==7'h16) || (r_sys_run_step==7'h17)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1259[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1289[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1223[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1157[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1133[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1217[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1247[8:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1319[8:0] );

									end
									else
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1187[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1211[8:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1271[8:0] );

									end
									else
									if((r_sys_run_step==7'hb) || (r_sys_run_step==7'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1193[8:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1277[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1283[8:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1307[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1163[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1139[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1241[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1181[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1169[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1151[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1145[8:0] );

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h17)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1446[8:0] );

									end
									else
									if((r_sys_run_step==7'h2e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1561[8:0] );

									end
									else
									if((r_sys_run_step==7'h27)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1526[8:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1486[8:0] );

									end
									else
									if((r_sys_run_step==7'h2b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1546[8:0] );

									end
									else
									if((r_sys_run_step==7'h25)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1516[8:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1436[8:0] );

									end
									else
									if((r_sys_run_step==7'h34)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1591[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1343[8:0] );

									end
									else
									if((r_sys_run_step==7'h39)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1616[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1416[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1331[8:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1471[8:0] );

									end
									else
									if((r_sys_run_step==7'h33)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1586[8:0] );

									end
									else
									if((r_sys_run_step==7'h22)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1501[8:0] );

									end
									else
									if((r_sys_run_step==7'h28)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1531[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1411[8:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1385[8:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1476[8:0] );

									end
									else
									if((r_sys_run_step==7'h32)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1581[8:0] );

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1596[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1406[8:0] );

									end
									else
									if((r_sys_run_step==7'h26)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1521[8:0] );

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1496[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1466[8:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1481[8:0] );

									end
									else
									if((r_sys_run_step==7'h2a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1541[8:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1456[8:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1379[8:0] );

									end
									else
									if((r_sys_run_step==7'h37)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1606[8:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1396[8:0] );

									end
									else
									if((r_sys_run_step==7'h3b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1626[8:0] );

									end
									else
									if((r_sys_run_step==7'h30)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1571[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1367[8:0] );

									end
									else
									if((r_sys_run_step==7'h36)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1601[8:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1451[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1349[8:0] );

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1441[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1431[8:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1391[8:0] );

									end
									else
									if((r_sys_run_step==7'h24)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1511[8:0] );

									end
									else
									if((r_sys_run_step==7'h31)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1576[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1355[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1337[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1426[8:0] );

									end
									else
									if((r_sys_run_step==7'h2f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1566[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1361[8:0] );

									end
									else
									if((r_sys_run_step==7'h2d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1556[8:0] );

									end
									else
									if((r_sys_run_step==7'h3a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1621[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1461[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1373[8:0] );

									end
									else
									if((r_sys_run_step==7'h29)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1536[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1421[8:0] );

									end
									else
									if((r_sys_run_step==7'h23)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1506[8:0] );

									end
									else
									if((r_sys_run_step==7'h2c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1551[8:0] );

									end
									else
									if((r_sys_run_step==7'h38)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1611[8:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1491[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1401[8:0] );

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1717[8:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1702[8:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1792[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1679[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1707[8:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1685[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1722[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1767[8:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1757[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1712[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1673[8:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1697[8:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1742[8:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1787[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1643[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1732[8:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1691[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1661[8:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1782[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1649[8:0] );

									end
									else
									if((r_sys_run_step==7'h16) || (r_sys_run_step==7'h17)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1747[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1655[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1667[8:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1762[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1737[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1727[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1772[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1637[8:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1777[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp14;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h4) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h38) || (r_sys_run_step==7'h3c) || (r_sys_run_step==7'h40) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h48) || (r_sys_run_step==7'h4c)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp259;

									end
									else
									if((r_sys_run_step==7'h1) || (r_sys_run_step==7'h3) || (r_sys_run_step==7'h5) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'h9) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h2b) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h2f) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h33) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h3b) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h3f) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h45) || (r_sys_run_step==7'h47) || (r_sys_run_step==7'h49) || (r_sys_run_step==7'h4b) || (r_sys_run_step==7'h4d) || (r_sys_run_step==7'h4f)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp263;

									end
									else
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h3e) || (r_sys_run_step==7'h42) || (r_sys_run_step==7'h46) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h4e)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp268;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h38)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp21_float;

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==7'h31)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp19_float;

									end
									else
									if((r_sys_run_step==7'h32)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==7'h36)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp30_float;

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp42_float;

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp24_float;

									end
									else
									if((r_sys_run_step==7'h27)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp28_float;

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp38_float;

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==7'h2b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp35_float;

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp32_float;

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp34_float;

									end
									else
									if((r_sys_run_step==7'h39)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp14_float;

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp40_float;

									end
									else
									if((r_sys_run_step==7'h2c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp31_float;

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp23_float;

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp43_float;

									end
									else
									if((r_sys_run_step==7'h2e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp22_float;

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp37_float;

									end
									else
									if((r_sys_run_step==7'h34)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp41_float;

									end
									else
									if((r_sys_run_step==7'h23)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp25_float;

									end
									else
									if((r_sys_run_step==7'h26)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==7'h30)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==7'h2a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp39_float;

									end
									else
									if((r_sys_run_step==7'h2d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp27_float;

									end
									else
									if((r_sys_run_step==7'h37)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp26_float;

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp18_float;

									end
									else
									if((r_sys_run_step==7'h22)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp29_float;

									end
									else
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'hb)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp1333;

									end
									else
									if((r_sys_run_step==7'h2f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp45_float;

									end
									else
									if((r_sys_run_step==7'h29)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp44_float;

									end
									else
									if((r_sys_run_step==7'h33)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp46_float;

									end
									else
									if((r_sys_run_step==7'h24)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp20_float;

									end
									else
									if((r_sys_run_step==7'h3a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==7'h28)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp36_float;

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp33_float;

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp47_float;

									end
									else
									if((r_sys_run_step==7'h3b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==7'h25)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp17_float;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'he)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==7'hc) || (r_sys_run_step==7'h16)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp19_float;

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp14_float;

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp10_float;

									end
									else
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'hb)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp1639;

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp17_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h4f)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h45)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h20)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h3b)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h1f)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h35: begin
							r_fld_u_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_uu_1_addr_1 <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_fld_uu_1_addr_1 <= $signed( w_sys_tmp16[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_fld_uu_1_datain_1 <= w_sys_tmp14;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_uu_1_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_fld_uu_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h35: begin
							r_fld_uu_1_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h4: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_11 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_11 <= w_sys_tmp6;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_11 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h47)) begin
										r_run_k_11 <= w_sys_tmp1120;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_11 <= w_sys_tmp1121;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h22)) begin
										r_run_k_11 <= w_sys_tmp1324;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_11 <= w_sys_tmp1325;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3b)) begin
										r_run_k_11 <= w_sys_tmp1630;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_11 <= w_sys_tmp1631;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1f)) begin
										r_run_k_11 <= w_sys_tmp1796;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_12 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_run_j_12 <= w_sys_tmp21;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_12 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h4) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h38) || (r_sys_run_step==7'h3c) || (r_sys_run_step==7'h40) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h48) || (r_sys_run_step==7'h4c)) begin
										r_run_j_12 <= w_sys_tmp277;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_n_13 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_n_13 <= w_sys_tmp252;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_mx_14 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_my_15 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_nlast_16 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_17 <= r_run_j_12;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_run_copy0_j_17 <= w_sys_tmp20;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_18 <= r_run_j_12;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h2b) || (r_sys_run_step==7'h2f) || (r_sys_run_step==7'h33) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h3b) || (r_sys_run_step==7'h3f) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h47) || (r_sys_run_step==7'h4b) || (r_sys_run_step==7'h4f)) begin
										r_run_copy0_j_18 <= w_sys_tmp274;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_19 <= r_run_j_12;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h3e) || (r_sys_run_step==7'h42) || (r_sys_run_step==7'h46) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h4e)) begin
										r_run_copy1_j_19 <= w_sys_tmp275;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy2_j_20 <= r_run_j_12;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1) || (r_sys_run_step==7'h5) || (r_sys_run_step==7'h9) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h45) || (r_sys_run_step==7'h49) || (r_sys_run_step==7'h4d)) begin
										r_run_copy2_j_20 <= w_sys_tmp276;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub08_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h19)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1259[9:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1289[9:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1271[9:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1301[9:0] );

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1313[9:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1277[9:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1283[9:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1307[9:0] );

									end
									else
									if((r_sys_run_step==7'h22)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1319[9:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1295[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h19<=r_sys_run_step && r_sys_run_step<=7'h22)) begin
										r_sub08_u_datain <= w_sys_tmp1129;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h19<=r_sys_run_step && r_sys_run_step<=7'h22)) begin
										r_sub08_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub08_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1757[9:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1747[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1762[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1792[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1772[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1782[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1787[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1767[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1777[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub08_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h2b)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp947[9:0] );

									end
									else
									if((r_sys_run_step==7'h29)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp935[9:0] );

									end
									else
									if((r_sys_run_step==7'h25)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp911[9:0] );

									end
									else
									if((r_sys_run_step==7'h26)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp917[9:0] );

									end
									else
									if((r_sys_run_step==7'h27)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp923[9:0] );

									end
									else
									if((r_sys_run_step==7'h28)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp929[9:0] );

									end
									else
									if((r_sys_run_step==7'h2f)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp971[9:0] );

									end
									else
									if((r_sys_run_step==7'h2a)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp941[9:0] );

									end
									else
									if((r_sys_run_step==7'h2d)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp959[9:0] );

									end
									else
									if((r_sys_run_step==7'h2c)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp953[9:0] );

									end
									else
									if((r_sys_run_step==7'h2e)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp965[9:0] );

									end
									else
									if((r_sys_run_step==7'h30)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp977[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h25<=r_sys_run_step && r_sys_run_step<=7'h30)) begin
										r_sub03_u_datain <= w_sys_tmp703;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h25<=r_sys_run_step && r_sys_run_step<=7'h30)) begin
										r_sub03_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub03_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1516[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1501[9:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1531[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1511[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1496[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1526[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1506[9:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1491[9:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1486[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1521[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h9)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub03_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1b)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp839[9:0] );

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp887[9:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp881[9:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp869[9:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp857[9:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp875[9:0] );

									end
									else
									if((r_sys_run_step==7'h24)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp905[9:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp833[9:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp863[9:0] );

									end
									else
									if((r_sys_run_step==7'h23)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp899[9:0] );

									end
									else
									if((r_sys_run_step==7'h22)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp893[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h1a<=r_sys_run_step && r_sys_run_step<=7'h24)) begin
										r_sub02_u_datain <= w_sys_tmp703;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h1a<=r_sys_run_step && r_sys_run_step<=7'h24)) begin
										r_sub02_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub02_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1446[9:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1441[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1461[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1476[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1466[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1481[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1451[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1471[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1456[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub02_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h19)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp839[9:0] );

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp821[9:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp809[9:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp803[9:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp833[9:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp791[9:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp767[9:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp797[9:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp815[9:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp785[9:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp761[9:0] );

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp827[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h19)) begin
										r_sub01_u_datain <= w_sys_tmp703;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h19)) begin
										r_sub01_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub01_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1431[9:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1396[9:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1436[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1411[9:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1391[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1421[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1406[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1416[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1401[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1426[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h9)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'hb)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp755[9:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp749[9:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp743[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp719[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp707[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp725[9:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp767[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp713[9:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp761[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp731[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp737[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp701[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub00_u_datain <= w_sys_tmp703;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub00_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub00_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1361[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1373[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1367[9:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1385[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1379[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1355[9:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1337[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1343[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1349[9:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1331[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h9)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub07_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h13)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1229[9:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1259[9:0] );

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1253[9:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1187[9:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1235[9:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1211[9:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1241[9:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1223[9:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1193[9:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1217[9:0] );

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1247[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h18)) begin
										r_sub07_u_datain <= w_sys_tmp1129;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h18)) begin
										r_sub07_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub07_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1717[9:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1747[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1712[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1732[9:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1702[9:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1697[9:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1742[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1737[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1727[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1707[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1722[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'ha)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub07_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub06_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'hc)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1187[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1139[9:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1193[9:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1181[9:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1175[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1157[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1133[9:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1169[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1163[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1127[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1151[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1145[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub06_u_datain <= w_sys_tmp1129;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub06_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub06_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1649[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1655[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1673[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1667[9:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1691[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1661[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1679[9:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1637[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1685[9:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1643[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h9)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub06_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub05_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h43)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1091[9:0] );

									end
									else
									if((r_sys_run_step==7'h3e)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1049[9:0] );

									end
									else
									if((r_sys_run_step==7'h46)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1109[9:0] );

									end
									else
									if((r_sys_run_step==7'h45)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1103[9:0] );

									end
									else
									if((r_sys_run_step==7'h44)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1097[9:0] );

									end
									else
									if((r_sys_run_step==7'h42)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1085[9:0] );

									end
									else
									if((r_sys_run_step==7'h3d)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1043[9:0] );

									end
									else
									if((r_sys_run_step==7'h40)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1073[9:0] );

									end
									else
									if((r_sys_run_step==7'h41)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1079[9:0] );

									end
									else
									if((r_sys_run_step==7'h3f)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1067[9:0] );

									end
									else
									if((r_sys_run_step==7'h47)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1115[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h3d<=r_sys_run_step && r_sys_run_step<=7'h47)) begin
										r_sub05_u_datain <= w_sys_tmp703;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h3d<=r_sys_run_step && r_sys_run_step<=7'h47)) begin
										r_sub05_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub05_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1586[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1621[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1626[9:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1591[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1601[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1606[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1596[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1616[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1611[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub05_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub04_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3a)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1037[9:0] );

									end
									else
									if((r_sys_run_step==7'h39)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1031[9:0] );

									end
									else
									if((r_sys_run_step==7'h36)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1013[9:0] );

									end
									else
									if((r_sys_run_step==7'h3c)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1049[9:0] );

									end
									else
									if((r_sys_run_step==7'h38)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1025[9:0] );

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1007[9:0] );

									end
									else
									if((r_sys_run_step==7'h33)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp995[9:0] );

									end
									else
									if((r_sys_run_step==7'h31)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp971[9:0] );

									end
									else
									if((r_sys_run_step==7'h3b)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1043[9:0] );

									end
									else
									if((r_sys_run_step==7'h37)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1019[9:0] );

									end
									else
									if((r_sys_run_step==7'h34)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1001[9:0] );

									end
									else
									if((r_sys_run_step==7'h32)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp977[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h31<=r_sys_run_step && r_sys_run_step<=7'h3c)) begin
										r_sub04_u_datain <= w_sys_tmp703;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h31<=r_sys_run_step && r_sys_run_step<=7'h3c)) begin
										r_sub04_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub04_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1556[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1571[9:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1536[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1576[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1561[9:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1581[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1551[9:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1541[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1546[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1566[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h9)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub04_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'hb)) begin
										r_sys_tmp0_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'hb)) begin
										r_sys_tmp0_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'hb)) begin
										r_sys_tmp1_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sys_tmp1_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'hb)) begin
										r_sys_tmp2_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sys_tmp2_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sys_tmp3_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sys_tmp3_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sys_tmp4_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sys_tmp4_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sys_tmp5_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_tmp5_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sys_tmp6_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_tmp6_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sys_tmp7_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sys_tmp7_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sys_tmp8_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sys_tmp8_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sys_tmp9_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_tmp9_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sys_tmp10_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_tmp10_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sys_tmp11_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp11_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sys_tmp12_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp12_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_tmp13_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp13_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_tmp14_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp14_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_tmp15_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp15_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_tmp16_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp16_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_tmp17_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp17_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sys_tmp18_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sys_tmp19_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'hc)) begin
										r_sys_tmp19_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sys_tmp20_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sys_tmp21_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sys_tmp22_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_tmp23_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_tmp24_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_tmp25_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_tmp26_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_tmp27_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp28_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp29_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp30_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp31_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp32_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp33_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp34_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp35_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp36_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp37_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp38_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp39_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp40_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp41_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp42_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp43_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp44_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp45_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp46_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp47_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
