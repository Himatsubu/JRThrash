/*
TimeStamp:	2013/12/16		12:59
*/


module FiltersJRT(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_main_req,	
	output                o_main_busy,	
	input  signed  [11:0] i_filter15_inputWave_addr,	
	input  signed  [15:0] i_filter15_inputWave_datain,	
	output signed  [15:0] o_filter15_inputWave_dataout,	
	input                 i_filter15_inputWave_r_w,	
	input  signed  [10:0] i_filter15_outputWave_addr,	
	input  signed  [15:0] i_filter15_outputWave_datain,	
	output signed  [15:0] o_filter15_outputWave_dataout,	
	input                 i_filter15_outputWave_r_w,	
	input  signed  [11:0] i_filter14_inputWave_addr,	
	input  signed  [15:0] i_filter14_inputWave_datain,	
	output signed  [15:0] o_filter14_inputWave_dataout,	
	input                 i_filter14_inputWave_r_w,	
	input  signed  [10:0] i_filter14_outputWave_addr,	
	input  signed  [15:0] i_filter14_outputWave_datain,	
	output signed  [15:0] o_filter14_outputWave_dataout,	
	input                 i_filter14_outputWave_r_w,	
	input  signed  [11:0] i_filter13_inputWave_addr,	
	input  signed  [15:0] i_filter13_inputWave_datain,	
	output signed  [15:0] o_filter13_inputWave_dataout,	
	input                 i_filter13_inputWave_r_w,	
	input  signed  [10:0] i_filter13_outputWave_addr,	
	input  signed  [15:0] i_filter13_outputWave_datain,	
	output signed  [15:0] o_filter13_outputWave_dataout,	
	input                 i_filter13_outputWave_r_w,	
	input  signed  [11:0] i_filter8_inputWave_addr,	
	input  signed  [15:0] i_filter8_inputWave_datain,	
	output signed  [15:0] o_filter8_inputWave_dataout,	
	input                 i_filter8_inputWave_r_w,	
	input  signed  [10:0] i_filter8_outputWave_addr,	
	input  signed  [15:0] i_filter8_outputWave_datain,	
	output signed  [15:0] o_filter8_outputWave_dataout,	
	input                 i_filter8_outputWave_r_w,	
	input  signed  [11:0] i_filter12_inputWave_addr,	
	input  signed  [15:0] i_filter12_inputWave_datain,	
	output signed  [15:0] o_filter12_inputWave_dataout,	
	input                 i_filter12_inputWave_r_w,	
	input  signed  [10:0] i_filter12_outputWave_addr,	
	input  signed  [15:0] i_filter12_outputWave_datain,	
	output signed  [15:0] o_filter12_outputWave_dataout,	
	input                 i_filter12_outputWave_r_w,	
	input  signed  [11:0] i_filter11_inputWave_addr,	
	input  signed  [15:0] i_filter11_inputWave_datain,	
	output signed  [15:0] o_filter11_inputWave_dataout,	
	input                 i_filter11_inputWave_r_w,	
	input  signed  [10:0] i_filter11_outputWave_addr,	
	input  signed  [15:0] i_filter11_outputWave_datain,	
	output signed  [15:0] o_filter11_outputWave_dataout,	
	input                 i_filter11_outputWave_r_w,	
	input  signed  [11:0] i_filter9_inputWave_addr,	
	input  signed  [15:0] i_filter9_inputWave_datain,	
	output signed  [15:0] o_filter9_inputWave_dataout,	
	input                 i_filter9_inputWave_r_w,	
	input  signed  [10:0] i_filter9_outputWave_addr,	
	input  signed  [15:0] i_filter9_outputWave_datain,	
	output signed  [15:0] o_filter9_outputWave_dataout,	
	input                 i_filter9_outputWave_r_w,	
	input  signed  [11:0] i_filter1_inputWave_addr,	
	input  signed  [15:0] i_filter1_inputWave_datain,	
	output signed  [15:0] o_filter1_inputWave_dataout,	
	input                 i_filter1_inputWave_r_w,	
	input  signed  [10:0] i_filter1_outputWave_addr,	
	input  signed  [15:0] i_filter1_outputWave_datain,	
	output signed  [15:0] o_filter1_outputWave_dataout,	
	input                 i_filter1_outputWave_r_w,	
	input  signed  [11:0] i_filter10_inputWave_addr,	
	input  signed  [15:0] i_filter10_inputWave_datain,	
	output signed  [15:0] o_filter10_inputWave_dataout,	
	input                 i_filter10_inputWave_r_w,	
	input  signed  [10:0] i_filter10_outputWave_addr,	
	input  signed  [15:0] i_filter10_outputWave_datain,	
	output signed  [15:0] o_filter10_outputWave_dataout,	
	input                 i_filter10_outputWave_r_w,	
	input  signed  [11:0] i_filter0_inputWave_addr,	
	input  signed  [15:0] i_filter0_inputWave_datain,	
	output signed  [15:0] o_filter0_inputWave_dataout,	
	input                 i_filter0_inputWave_r_w,	
	input  signed  [10:0] i_filter0_outputWave_addr,	
	input  signed  [15:0] i_filter0_outputWave_datain,	
	output signed  [15:0] o_filter0_outputWave_dataout,	
	input                 i_filter0_outputWave_r_w,	
	input  signed  [11:0] i_filter3_inputWave_addr,	
	input  signed  [15:0] i_filter3_inputWave_datain,	
	output signed  [15:0] o_filter3_inputWave_dataout,	
	input                 i_filter3_inputWave_r_w,	
	input  signed  [10:0] i_filter3_outputWave_addr,	
	input  signed  [15:0] i_filter3_outputWave_datain,	
	output signed  [15:0] o_filter3_outputWave_dataout,	
	input                 i_filter3_outputWave_r_w,	
	input  signed  [11:0] i_filter2_inputWave_addr,	
	input  signed  [15:0] i_filter2_inputWave_datain,	
	output signed  [15:0] o_filter2_inputWave_dataout,	
	input                 i_filter2_inputWave_r_w,	
	input  signed  [10:0] i_filter2_outputWave_addr,	
	input  signed  [15:0] i_filter2_outputWave_datain,	
	output signed  [15:0] o_filter2_outputWave_dataout,	
	input                 i_filter2_outputWave_r_w,	
	input  signed  [11:0] i_filter5_inputWave_addr,	
	input  signed  [15:0] i_filter5_inputWave_datain,	
	output signed  [15:0] o_filter5_inputWave_dataout,	
	input                 i_filter5_inputWave_r_w,	
	input  signed  [10:0] i_filter5_outputWave_addr,	
	input  signed  [15:0] i_filter5_outputWave_datain,	
	output signed  [15:0] o_filter5_outputWave_dataout,	
	input                 i_filter5_outputWave_r_w,	
	input  signed  [11:0] i_filter4_inputWave_addr,	
	input  signed  [15:0] i_filter4_inputWave_datain,	
	output signed  [15:0] o_filter4_inputWave_dataout,	
	input                 i_filter4_inputWave_r_w,	
	input  signed  [10:0] i_filter4_outputWave_addr,	
	input  signed  [15:0] i_filter4_outputWave_datain,	
	output signed  [15:0] o_filter4_outputWave_dataout,	
	input                 i_filter4_outputWave_r_w,	
	input  signed  [11:0] i_filter7_inputWave_addr,	
	input  signed  [15:0] i_filter7_inputWave_datain,	
	output signed  [15:0] o_filter7_inputWave_dataout,	
	input                 i_filter7_inputWave_r_w,	
	input  signed  [10:0] i_filter7_outputWave_addr,	
	input  signed  [15:0] i_filter7_outputWave_datain,	
	output signed  [15:0] o_filter7_outputWave_dataout,	
	input                 i_filter7_outputWave_r_w,	
	input  signed  [11:0] i_filter6_inputWave_addr,	
	input  signed  [15:0] i_filter6_inputWave_datain,	
	output signed  [15:0] o_filter6_inputWave_dataout,	
	input                 i_filter6_inputWave_r_w,	
	input  signed  [10:0] i_filter6_outputWave_addr,	
	input  signed  [15:0] i_filter6_outputWave_datain,	
	output signed  [15:0] o_filter6_outputWave_dataout,	
	input                 i_filter6_outputWave_r_w	
);

	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_main_caller;
	reg                r_sys_main_req;
	reg         [ 2:0] r_sys_main_phase;
	reg         [ 4:0] r_sys_main_stage;
	reg         [ 1:0] r_sys_main_step;
	reg                r_sys_main_busy;
	wire        [ 4:0] w_sys_main_stage_p1;
	wire        [ 1:0] w_sys_main_step_p1;
	reg                r_filter15_run_req;
	wire               w_filter15_run_busy;
	wire signed [11:0] w_filter15_inputWave_addr;
	reg  signed [11:0] r_filter15_inputWave_addr;
	wire signed [15:0] w_filter15_inputWave_datain;
	reg  signed [15:0] r_filter15_inputWave_datain;
	wire signed [15:0] w_filter15_inputWave_dataout;
	wire               w_filter15_inputWave_r_w;
	reg                r_filter15_inputWave_r_w;
	wire signed [10:0] w_filter15_outputWave_addr;
	reg  signed [10:0] r_filter15_outputWave_addr;
	wire signed [15:0] w_filter15_outputWave_datain;
	reg  signed [15:0] r_filter15_outputWave_datain;
	wire signed [15:0] w_filter15_outputWave_dataout;
	wire               w_filter15_outputWave_r_w;
	reg                r_filter15_outputWave_r_w;
	wire signed [ 8:0] w_filter15_filterCoef_addr;
	reg  signed [ 8:0] r_filter15_filterCoef_addr;
	wire signed [15:0] w_filter15_filterCoef_datain;
	reg  signed [15:0] r_filter15_filterCoef_datain;
	wire signed [15:0] w_filter15_filterCoef_dataout;
	wire               w_filter15_filterCoef_r_w;
	reg                r_filter15_filterCoef_r_w;
	reg                r_filter14_run_req;
	wire               w_filter14_run_busy;
	wire signed [11:0] w_filter14_inputWave_addr;
	reg  signed [11:0] r_filter14_inputWave_addr;
	wire signed [15:0] w_filter14_inputWave_datain;
	reg  signed [15:0] r_filter14_inputWave_datain;
	wire signed [15:0] w_filter14_inputWave_dataout;
	wire               w_filter14_inputWave_r_w;
	reg                r_filter14_inputWave_r_w;
	wire signed [10:0] w_filter14_outputWave_addr;
	reg  signed [10:0] r_filter14_outputWave_addr;
	wire signed [15:0] w_filter14_outputWave_datain;
	reg  signed [15:0] r_filter14_outputWave_datain;
	wire signed [15:0] w_filter14_outputWave_dataout;
	wire               w_filter14_outputWave_r_w;
	reg                r_filter14_outputWave_r_w;
	wire signed [ 8:0] w_filter14_filterCoef_addr;
	reg  signed [ 8:0] r_filter14_filterCoef_addr;
	wire signed [15:0] w_filter14_filterCoef_datain;
	reg  signed [15:0] r_filter14_filterCoef_datain;
	wire signed [15:0] w_filter14_filterCoef_dataout;
	wire               w_filter14_filterCoef_r_w;
	reg                r_filter14_filterCoef_r_w;
	reg                r_filter13_run_req;
	wire               w_filter13_run_busy;
	wire signed [11:0] w_filter13_inputWave_addr;
	reg  signed [11:0] r_filter13_inputWave_addr;
	wire signed [15:0] w_filter13_inputWave_datain;
	reg  signed [15:0] r_filter13_inputWave_datain;
	wire signed [15:0] w_filter13_inputWave_dataout;
	wire               w_filter13_inputWave_r_w;
	reg                r_filter13_inputWave_r_w;
	wire signed [10:0] w_filter13_outputWave_addr;
	reg  signed [10:0] r_filter13_outputWave_addr;
	wire signed [15:0] w_filter13_outputWave_datain;
	reg  signed [15:0] r_filter13_outputWave_datain;
	wire signed [15:0] w_filter13_outputWave_dataout;
	wire               w_filter13_outputWave_r_w;
	reg                r_filter13_outputWave_r_w;
	wire signed [ 8:0] w_filter13_filterCoef_addr;
	reg  signed [ 8:0] r_filter13_filterCoef_addr;
	wire signed [15:0] w_filter13_filterCoef_datain;
	reg  signed [15:0] r_filter13_filterCoef_datain;
	wire signed [15:0] w_filter13_filterCoef_dataout;
	wire               w_filter13_filterCoef_r_w;
	reg                r_filter13_filterCoef_r_w;
	reg                r_filter8_run_req;
	wire               w_filter8_run_busy;
	wire signed [11:0] w_filter8_inputWave_addr;
	reg  signed [11:0] r_filter8_inputWave_addr;
	wire signed [15:0] w_filter8_inputWave_datain;
	reg  signed [15:0] r_filter8_inputWave_datain;
	wire signed [15:0] w_filter8_inputWave_dataout;
	wire               w_filter8_inputWave_r_w;
	reg                r_filter8_inputWave_r_w;
	wire signed [10:0] w_filter8_outputWave_addr;
	reg  signed [10:0] r_filter8_outputWave_addr;
	wire signed [15:0] w_filter8_outputWave_datain;
	reg  signed [15:0] r_filter8_outputWave_datain;
	wire signed [15:0] w_filter8_outputWave_dataout;
	wire               w_filter8_outputWave_r_w;
	reg                r_filter8_outputWave_r_w;
	wire signed [ 8:0] w_filter8_filterCoef_addr;
	reg  signed [ 8:0] r_filter8_filterCoef_addr;
	wire signed [15:0] w_filter8_filterCoef_datain;
	reg  signed [15:0] r_filter8_filterCoef_datain;
	wire signed [15:0] w_filter8_filterCoef_dataout;
	wire               w_filter8_filterCoef_r_w;
	reg                r_filter8_filterCoef_r_w;
	reg                r_filter12_run_req;
	wire               w_filter12_run_busy;
	wire signed [11:0] w_filter12_inputWave_addr;
	reg  signed [11:0] r_filter12_inputWave_addr;
	wire signed [15:0] w_filter12_inputWave_datain;
	reg  signed [15:0] r_filter12_inputWave_datain;
	wire signed [15:0] w_filter12_inputWave_dataout;
	wire               w_filter12_inputWave_r_w;
	reg                r_filter12_inputWave_r_w;
	wire signed [10:0] w_filter12_outputWave_addr;
	reg  signed [10:0] r_filter12_outputWave_addr;
	wire signed [15:0] w_filter12_outputWave_datain;
	reg  signed [15:0] r_filter12_outputWave_datain;
	wire signed [15:0] w_filter12_outputWave_dataout;
	wire               w_filter12_outputWave_r_w;
	reg                r_filter12_outputWave_r_w;
	wire signed [ 8:0] w_filter12_filterCoef_addr;
	reg  signed [ 8:0] r_filter12_filterCoef_addr;
	wire signed [15:0] w_filter12_filterCoef_datain;
	reg  signed [15:0] r_filter12_filterCoef_datain;
	wire signed [15:0] w_filter12_filterCoef_dataout;
	wire               w_filter12_filterCoef_r_w;
	reg                r_filter12_filterCoef_r_w;
	reg                r_filter11_run_req;
	wire               w_filter11_run_busy;
	wire signed [11:0] w_filter11_inputWave_addr;
	reg  signed [11:0] r_filter11_inputWave_addr;
	wire signed [15:0] w_filter11_inputWave_datain;
	reg  signed [15:0] r_filter11_inputWave_datain;
	wire signed [15:0] w_filter11_inputWave_dataout;
	wire               w_filter11_inputWave_r_w;
	reg                r_filter11_inputWave_r_w;
	wire signed [10:0] w_filter11_outputWave_addr;
	reg  signed [10:0] r_filter11_outputWave_addr;
	wire signed [15:0] w_filter11_outputWave_datain;
	reg  signed [15:0] r_filter11_outputWave_datain;
	wire signed [15:0] w_filter11_outputWave_dataout;
	wire               w_filter11_outputWave_r_w;
	reg                r_filter11_outputWave_r_w;
	wire signed [ 8:0] w_filter11_filterCoef_addr;
	reg  signed [ 8:0] r_filter11_filterCoef_addr;
	wire signed [15:0] w_filter11_filterCoef_datain;
	reg  signed [15:0] r_filter11_filterCoef_datain;
	wire signed [15:0] w_filter11_filterCoef_dataout;
	wire               w_filter11_filterCoef_r_w;
	reg                r_filter11_filterCoef_r_w;
	reg                r_filter9_run_req;
	wire               w_filter9_run_busy;
	wire signed [11:0] w_filter9_inputWave_addr;
	reg  signed [11:0] r_filter9_inputWave_addr;
	wire signed [15:0] w_filter9_inputWave_datain;
	reg  signed [15:0] r_filter9_inputWave_datain;
	wire signed [15:0] w_filter9_inputWave_dataout;
	wire               w_filter9_inputWave_r_w;
	reg                r_filter9_inputWave_r_w;
	wire signed [10:0] w_filter9_outputWave_addr;
	reg  signed [10:0] r_filter9_outputWave_addr;
	wire signed [15:0] w_filter9_outputWave_datain;
	reg  signed [15:0] r_filter9_outputWave_datain;
	wire signed [15:0] w_filter9_outputWave_dataout;
	wire               w_filter9_outputWave_r_w;
	reg                r_filter9_outputWave_r_w;
	wire signed [ 8:0] w_filter9_filterCoef_addr;
	reg  signed [ 8:0] r_filter9_filterCoef_addr;
	wire signed [15:0] w_filter9_filterCoef_datain;
	reg  signed [15:0] r_filter9_filterCoef_datain;
	wire signed [15:0] w_filter9_filterCoef_dataout;
	wire               w_filter9_filterCoef_r_w;
	reg                r_filter9_filterCoef_r_w;
	reg                r_filter1_run_req;
	wire               w_filter1_run_busy;
	wire signed [11:0] w_filter1_inputWave_addr;
	reg  signed [11:0] r_filter1_inputWave_addr;
	wire signed [15:0] w_filter1_inputWave_datain;
	reg  signed [15:0] r_filter1_inputWave_datain;
	wire signed [15:0] w_filter1_inputWave_dataout;
	wire               w_filter1_inputWave_r_w;
	reg                r_filter1_inputWave_r_w;
	wire signed [10:0] w_filter1_outputWave_addr;
	reg  signed [10:0] r_filter1_outputWave_addr;
	wire signed [15:0] w_filter1_outputWave_datain;
	reg  signed [15:0] r_filter1_outputWave_datain;
	wire signed [15:0] w_filter1_outputWave_dataout;
	wire               w_filter1_outputWave_r_w;
	reg                r_filter1_outputWave_r_w;
	wire signed [ 8:0] w_filter1_filterCoef_addr;
	reg  signed [ 8:0] r_filter1_filterCoef_addr;
	wire signed [15:0] w_filter1_filterCoef_datain;
	reg  signed [15:0] r_filter1_filterCoef_datain;
	wire signed [15:0] w_filter1_filterCoef_dataout;
	wire               w_filter1_filterCoef_r_w;
	reg                r_filter1_filterCoef_r_w;
	reg                r_filter10_run_req;
	wire               w_filter10_run_busy;
	wire signed [11:0] w_filter10_inputWave_addr;
	reg  signed [11:0] r_filter10_inputWave_addr;
	wire signed [15:0] w_filter10_inputWave_datain;
	reg  signed [15:0] r_filter10_inputWave_datain;
	wire signed [15:0] w_filter10_inputWave_dataout;
	wire               w_filter10_inputWave_r_w;
	reg                r_filter10_inputWave_r_w;
	wire signed [10:0] w_filter10_outputWave_addr;
	reg  signed [10:0] r_filter10_outputWave_addr;
	wire signed [15:0] w_filter10_outputWave_datain;
	reg  signed [15:0] r_filter10_outputWave_datain;
	wire signed [15:0] w_filter10_outputWave_dataout;
	wire               w_filter10_outputWave_r_w;
	reg                r_filter10_outputWave_r_w;
	wire signed [ 8:0] w_filter10_filterCoef_addr;
	reg  signed [ 8:0] r_filter10_filterCoef_addr;
	wire signed [15:0] w_filter10_filterCoef_datain;
	reg  signed [15:0] r_filter10_filterCoef_datain;
	wire signed [15:0] w_filter10_filterCoef_dataout;
	wire               w_filter10_filterCoef_r_w;
	reg                r_filter10_filterCoef_r_w;
	reg                r_filter0_run_req;
	wire               w_filter0_run_busy;
	wire signed [11:0] w_filter0_inputWave_addr;
	reg  signed [11:0] r_filter0_inputWave_addr;
	wire signed [15:0] w_filter0_inputWave_datain;
	reg  signed [15:0] r_filter0_inputWave_datain;
	wire signed [15:0] w_filter0_inputWave_dataout;
	wire               w_filter0_inputWave_r_w;
	reg                r_filter0_inputWave_r_w;
	wire signed [10:0] w_filter0_outputWave_addr;
	reg  signed [10:0] r_filter0_outputWave_addr;
	wire signed [15:0] w_filter0_outputWave_datain;
	reg  signed [15:0] r_filter0_outputWave_datain;
	wire signed [15:0] w_filter0_outputWave_dataout;
	wire               w_filter0_outputWave_r_w;
	reg                r_filter0_outputWave_r_w;
	wire signed [ 8:0] w_filter0_filterCoef_addr;
	reg  signed [ 8:0] r_filter0_filterCoef_addr;
	wire signed [15:0] w_filter0_filterCoef_datain;
	reg  signed [15:0] r_filter0_filterCoef_datain;
	wire signed [15:0] w_filter0_filterCoef_dataout;
	wire               w_filter0_filterCoef_r_w;
	reg                r_filter0_filterCoef_r_w;
	reg                r_filter3_run_req;
	wire               w_filter3_run_busy;
	wire signed [11:0] w_filter3_inputWave_addr;
	reg  signed [11:0] r_filter3_inputWave_addr;
	wire signed [15:0] w_filter3_inputWave_datain;
	reg  signed [15:0] r_filter3_inputWave_datain;
	wire signed [15:0] w_filter3_inputWave_dataout;
	wire               w_filter3_inputWave_r_w;
	reg                r_filter3_inputWave_r_w;
	wire signed [10:0] w_filter3_outputWave_addr;
	reg  signed [10:0] r_filter3_outputWave_addr;
	wire signed [15:0] w_filter3_outputWave_datain;
	reg  signed [15:0] r_filter3_outputWave_datain;
	wire signed [15:0] w_filter3_outputWave_dataout;
	wire               w_filter3_outputWave_r_w;
	reg                r_filter3_outputWave_r_w;
	wire signed [ 8:0] w_filter3_filterCoef_addr;
	reg  signed [ 8:0] r_filter3_filterCoef_addr;
	wire signed [15:0] w_filter3_filterCoef_datain;
	reg  signed [15:0] r_filter3_filterCoef_datain;
	wire signed [15:0] w_filter3_filterCoef_dataout;
	wire               w_filter3_filterCoef_r_w;
	reg                r_filter3_filterCoef_r_w;
	reg                r_filter2_run_req;
	wire               w_filter2_run_busy;
	wire signed [11:0] w_filter2_inputWave_addr;
	reg  signed [11:0] r_filter2_inputWave_addr;
	wire signed [15:0] w_filter2_inputWave_datain;
	reg  signed [15:0] r_filter2_inputWave_datain;
	wire signed [15:0] w_filter2_inputWave_dataout;
	wire               w_filter2_inputWave_r_w;
	reg                r_filter2_inputWave_r_w;
	wire signed [10:0] w_filter2_outputWave_addr;
	reg  signed [10:0] r_filter2_outputWave_addr;
	wire signed [15:0] w_filter2_outputWave_datain;
	reg  signed [15:0] r_filter2_outputWave_datain;
	wire signed [15:0] w_filter2_outputWave_dataout;
	wire               w_filter2_outputWave_r_w;
	reg                r_filter2_outputWave_r_w;
	wire signed [ 8:0] w_filter2_filterCoef_addr;
	reg  signed [ 8:0] r_filter2_filterCoef_addr;
	wire signed [15:0] w_filter2_filterCoef_datain;
	reg  signed [15:0] r_filter2_filterCoef_datain;
	wire signed [15:0] w_filter2_filterCoef_dataout;
	wire               w_filter2_filterCoef_r_w;
	reg                r_filter2_filterCoef_r_w;
	reg                r_filter5_run_req;
	wire               w_filter5_run_busy;
	wire signed [11:0] w_filter5_inputWave_addr;
	reg  signed [11:0] r_filter5_inputWave_addr;
	wire signed [15:0] w_filter5_inputWave_datain;
	reg  signed [15:0] r_filter5_inputWave_datain;
	wire signed [15:0] w_filter5_inputWave_dataout;
	wire               w_filter5_inputWave_r_w;
	reg                r_filter5_inputWave_r_w;
	wire signed [10:0] w_filter5_outputWave_addr;
	reg  signed [10:0] r_filter5_outputWave_addr;
	wire signed [15:0] w_filter5_outputWave_datain;
	reg  signed [15:0] r_filter5_outputWave_datain;
	wire signed [15:0] w_filter5_outputWave_dataout;
	wire               w_filter5_outputWave_r_w;
	reg                r_filter5_outputWave_r_w;
	wire signed [ 8:0] w_filter5_filterCoef_addr;
	reg  signed [ 8:0] r_filter5_filterCoef_addr;
	wire signed [15:0] w_filter5_filterCoef_datain;
	reg  signed [15:0] r_filter5_filterCoef_datain;
	wire signed [15:0] w_filter5_filterCoef_dataout;
	wire               w_filter5_filterCoef_r_w;
	reg                r_filter5_filterCoef_r_w;
	reg                r_filter4_run_req;
	wire               w_filter4_run_busy;
	wire signed [11:0] w_filter4_inputWave_addr;
	reg  signed [11:0] r_filter4_inputWave_addr;
	wire signed [15:0] w_filter4_inputWave_datain;
	reg  signed [15:0] r_filter4_inputWave_datain;
	wire signed [15:0] w_filter4_inputWave_dataout;
	wire               w_filter4_inputWave_r_w;
	reg                r_filter4_inputWave_r_w;
	wire signed [10:0] w_filter4_outputWave_addr;
	reg  signed [10:0] r_filter4_outputWave_addr;
	wire signed [15:0] w_filter4_outputWave_datain;
	reg  signed [15:0] r_filter4_outputWave_datain;
	wire signed [15:0] w_filter4_outputWave_dataout;
	wire               w_filter4_outputWave_r_w;
	reg                r_filter4_outputWave_r_w;
	wire signed [ 8:0] w_filter4_filterCoef_addr;
	reg  signed [ 8:0] r_filter4_filterCoef_addr;
	wire signed [15:0] w_filter4_filterCoef_datain;
	reg  signed [15:0] r_filter4_filterCoef_datain;
	wire signed [15:0] w_filter4_filterCoef_dataout;
	wire               w_filter4_filterCoef_r_w;
	reg                r_filter4_filterCoef_r_w;
	reg                r_filter7_run_req;
	wire               w_filter7_run_busy;
	wire signed [11:0] w_filter7_inputWave_addr;
	reg  signed [11:0] r_filter7_inputWave_addr;
	wire signed [15:0] w_filter7_inputWave_datain;
	reg  signed [15:0] r_filter7_inputWave_datain;
	wire signed [15:0] w_filter7_inputWave_dataout;
	wire               w_filter7_inputWave_r_w;
	reg                r_filter7_inputWave_r_w;
	wire signed [10:0] w_filter7_outputWave_addr;
	reg  signed [10:0] r_filter7_outputWave_addr;
	wire signed [15:0] w_filter7_outputWave_datain;
	reg  signed [15:0] r_filter7_outputWave_datain;
	wire signed [15:0] w_filter7_outputWave_dataout;
	wire               w_filter7_outputWave_r_w;
	reg                r_filter7_outputWave_r_w;
	wire signed [ 8:0] w_filter7_filterCoef_addr;
	reg  signed [ 8:0] r_filter7_filterCoef_addr;
	wire signed [15:0] w_filter7_filterCoef_datain;
	reg  signed [15:0] r_filter7_filterCoef_datain;
	wire signed [15:0] w_filter7_filterCoef_dataout;
	wire               w_filter7_filterCoef_r_w;
	reg                r_filter7_filterCoef_r_w;
	reg                r_filter6_run_req;
	wire               w_filter6_run_busy;
	wire signed [11:0] w_filter6_inputWave_addr;
	reg  signed [11:0] r_filter6_inputWave_addr;
	wire signed [15:0] w_filter6_inputWave_datain;
	reg  signed [15:0] r_filter6_inputWave_datain;
	wire signed [15:0] w_filter6_inputWave_dataout;
	wire               w_filter6_inputWave_r_w;
	reg                r_filter6_inputWave_r_w;
	wire signed [10:0] w_filter6_outputWave_addr;
	reg  signed [10:0] r_filter6_outputWave_addr;
	wire signed [15:0] w_filter6_outputWave_datain;
	reg  signed [15:0] r_filter6_outputWave_datain;
	wire signed [15:0] w_filter6_outputWave_dataout;
	wire               w_filter6_outputWave_r_w;
	reg                r_filter6_outputWave_r_w;
	wire signed [ 8:0] w_filter6_filterCoef_addr;
	reg  signed [ 8:0] r_filter6_filterCoef_addr;
	wire signed [15:0] w_filter6_filterCoef_datain;
	reg  signed [15:0] r_filter6_filterCoef_datain;
	wire signed [15:0] w_filter6_filterCoef_dataout;
	wire               w_filter6_filterCoef_r_w;
	reg                r_filter6_filterCoef_r_w;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_main_busy = r_sys_main_busy;
	assign w_sys_main_stage_p1 = (r_sys_main_stage + 5'h1);
	assign w_sys_main_step_p1 = (r_sys_main_step + 2'h1);
	assign w_filter15_inputWave_addr = ( (|r_sys_processing_methodID) ? r_filter15_inputWave_addr : i_filter15_inputWave_addr ) ;
	assign w_filter15_inputWave_datain = ( (|r_sys_processing_methodID) ? r_filter15_inputWave_datain : i_filter15_inputWave_datain ) ;
	assign o_filter15_inputWave_dataout = w_filter15_inputWave_dataout;
	assign w_filter15_inputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter15_inputWave_r_w : i_filter15_inputWave_r_w ) ;
	assign w_filter15_outputWave_addr = ( (|r_sys_processing_methodID) ? r_filter15_outputWave_addr : i_filter15_outputWave_addr ) ;
	assign w_filter15_outputWave_datain = ( (|r_sys_processing_methodID) ? r_filter15_outputWave_datain : i_filter15_outputWave_datain ) ;
	assign o_filter15_outputWave_dataout = w_filter15_outputWave_dataout;
	assign w_filter15_outputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter15_outputWave_r_w : i_filter15_outputWave_r_w ) ;
	assign w_filter15_filterCoef_addr = ( (|r_sys_processing_methodID) ? r_filter15_filterCoef_addr : 9'sh0 ) ;
	assign w_filter15_filterCoef_datain = ( (|r_sys_processing_methodID) ? r_filter15_filterCoef_datain : 16'sh0 ) ;
	assign w_filter15_filterCoef_r_w = ( (|r_sys_processing_methodID) ? r_filter15_filterCoef_r_w : 1'h0 ) ;
	assign w_filter14_inputWave_addr = ( (|r_sys_processing_methodID) ? r_filter14_inputWave_addr : i_filter14_inputWave_addr ) ;
	assign w_filter14_inputWave_datain = ( (|r_sys_processing_methodID) ? r_filter14_inputWave_datain : i_filter14_inputWave_datain ) ;
	assign o_filter14_inputWave_dataout = w_filter14_inputWave_dataout;
	assign w_filter14_inputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter14_inputWave_r_w : i_filter14_inputWave_r_w ) ;
	assign w_filter14_outputWave_addr = ( (|r_sys_processing_methodID) ? r_filter14_outputWave_addr : i_filter14_outputWave_addr ) ;
	assign w_filter14_outputWave_datain = ( (|r_sys_processing_methodID) ? r_filter14_outputWave_datain : i_filter14_outputWave_datain ) ;
	assign o_filter14_outputWave_dataout = w_filter14_outputWave_dataout;
	assign w_filter14_outputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter14_outputWave_r_w : i_filter14_outputWave_r_w ) ;
	assign w_filter14_filterCoef_addr = ( (|r_sys_processing_methodID) ? r_filter14_filterCoef_addr : 9'sh0 ) ;
	assign w_filter14_filterCoef_datain = ( (|r_sys_processing_methodID) ? r_filter14_filterCoef_datain : 16'sh0 ) ;
	assign w_filter14_filterCoef_r_w = ( (|r_sys_processing_methodID) ? r_filter14_filterCoef_r_w : 1'h0 ) ;
	assign w_filter13_inputWave_addr = ( (|r_sys_processing_methodID) ? r_filter13_inputWave_addr : i_filter13_inputWave_addr ) ;
	assign w_filter13_inputWave_datain = ( (|r_sys_processing_methodID) ? r_filter13_inputWave_datain : i_filter13_inputWave_datain ) ;
	assign o_filter13_inputWave_dataout = w_filter13_inputWave_dataout;
	assign w_filter13_inputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter13_inputWave_r_w : i_filter13_inputWave_r_w ) ;
	assign w_filter13_outputWave_addr = ( (|r_sys_processing_methodID) ? r_filter13_outputWave_addr : i_filter13_outputWave_addr ) ;
	assign w_filter13_outputWave_datain = ( (|r_sys_processing_methodID) ? r_filter13_outputWave_datain : i_filter13_outputWave_datain ) ;
	assign o_filter13_outputWave_dataout = w_filter13_outputWave_dataout;
	assign w_filter13_outputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter13_outputWave_r_w : i_filter13_outputWave_r_w ) ;
	assign w_filter13_filterCoef_addr = ( (|r_sys_processing_methodID) ? r_filter13_filterCoef_addr : 9'sh0 ) ;
	assign w_filter13_filterCoef_datain = ( (|r_sys_processing_methodID) ? r_filter13_filterCoef_datain : 16'sh0 ) ;
	assign w_filter13_filterCoef_r_w = ( (|r_sys_processing_methodID) ? r_filter13_filterCoef_r_w : 1'h0 ) ;
	assign w_filter8_inputWave_addr = ( (|r_sys_processing_methodID) ? r_filter8_inputWave_addr : i_filter8_inputWave_addr ) ;
	assign w_filter8_inputWave_datain = ( (|r_sys_processing_methodID) ? r_filter8_inputWave_datain : i_filter8_inputWave_datain ) ;
	assign o_filter8_inputWave_dataout = w_filter8_inputWave_dataout;
	assign w_filter8_inputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter8_inputWave_r_w : i_filter8_inputWave_r_w ) ;
	assign w_filter8_outputWave_addr = ( (|r_sys_processing_methodID) ? r_filter8_outputWave_addr : i_filter8_outputWave_addr ) ;
	assign w_filter8_outputWave_datain = ( (|r_sys_processing_methodID) ? r_filter8_outputWave_datain : i_filter8_outputWave_datain ) ;
	assign o_filter8_outputWave_dataout = w_filter8_outputWave_dataout;
	assign w_filter8_outputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter8_outputWave_r_w : i_filter8_outputWave_r_w ) ;
	assign w_filter8_filterCoef_addr = ( (|r_sys_processing_methodID) ? r_filter8_filterCoef_addr : 9'sh0 ) ;
	assign w_filter8_filterCoef_datain = ( (|r_sys_processing_methodID) ? r_filter8_filterCoef_datain : 16'sh0 ) ;
	assign w_filter8_filterCoef_r_w = ( (|r_sys_processing_methodID) ? r_filter8_filterCoef_r_w : 1'h0 ) ;
	assign w_filter12_inputWave_addr = ( (|r_sys_processing_methodID) ? r_filter12_inputWave_addr : i_filter12_inputWave_addr ) ;
	assign w_filter12_inputWave_datain = ( (|r_sys_processing_methodID) ? r_filter12_inputWave_datain : i_filter12_inputWave_datain ) ;
	assign o_filter12_inputWave_dataout = w_filter12_inputWave_dataout;
	assign w_filter12_inputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter12_inputWave_r_w : i_filter12_inputWave_r_w ) ;
	assign w_filter12_outputWave_addr = ( (|r_sys_processing_methodID) ? r_filter12_outputWave_addr : i_filter12_outputWave_addr ) ;
	assign w_filter12_outputWave_datain = ( (|r_sys_processing_methodID) ? r_filter12_outputWave_datain : i_filter12_outputWave_datain ) ;
	assign o_filter12_outputWave_dataout = w_filter12_outputWave_dataout;
	assign w_filter12_outputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter12_outputWave_r_w : i_filter12_outputWave_r_w ) ;
	assign w_filter12_filterCoef_addr = ( (|r_sys_processing_methodID) ? r_filter12_filterCoef_addr : 9'sh0 ) ;
	assign w_filter12_filterCoef_datain = ( (|r_sys_processing_methodID) ? r_filter12_filterCoef_datain : 16'sh0 ) ;
	assign w_filter12_filterCoef_r_w = ( (|r_sys_processing_methodID) ? r_filter12_filterCoef_r_w : 1'h0 ) ;
	assign w_filter11_inputWave_addr = ( (|r_sys_processing_methodID) ? r_filter11_inputWave_addr : i_filter11_inputWave_addr ) ;
	assign w_filter11_inputWave_datain = ( (|r_sys_processing_methodID) ? r_filter11_inputWave_datain : i_filter11_inputWave_datain ) ;
	assign o_filter11_inputWave_dataout = w_filter11_inputWave_dataout;
	assign w_filter11_inputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter11_inputWave_r_w : i_filter11_inputWave_r_w ) ;
	assign w_filter11_outputWave_addr = ( (|r_sys_processing_methodID) ? r_filter11_outputWave_addr : i_filter11_outputWave_addr ) ;
	assign w_filter11_outputWave_datain = ( (|r_sys_processing_methodID) ? r_filter11_outputWave_datain : i_filter11_outputWave_datain ) ;
	assign o_filter11_outputWave_dataout = w_filter11_outputWave_dataout;
	assign w_filter11_outputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter11_outputWave_r_w : i_filter11_outputWave_r_w ) ;
	assign w_filter11_filterCoef_addr = ( (|r_sys_processing_methodID) ? r_filter11_filterCoef_addr : 9'sh0 ) ;
	assign w_filter11_filterCoef_datain = ( (|r_sys_processing_methodID) ? r_filter11_filterCoef_datain : 16'sh0 ) ;
	assign w_filter11_filterCoef_r_w = ( (|r_sys_processing_methodID) ? r_filter11_filterCoef_r_w : 1'h0 ) ;
	assign w_filter9_inputWave_addr = ( (|r_sys_processing_methodID) ? r_filter9_inputWave_addr : i_filter9_inputWave_addr ) ;
	assign w_filter9_inputWave_datain = ( (|r_sys_processing_methodID) ? r_filter9_inputWave_datain : i_filter9_inputWave_datain ) ;
	assign o_filter9_inputWave_dataout = w_filter9_inputWave_dataout;
	assign w_filter9_inputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter9_inputWave_r_w : i_filter9_inputWave_r_w ) ;
	assign w_filter9_outputWave_addr = ( (|r_sys_processing_methodID) ? r_filter9_outputWave_addr : i_filter9_outputWave_addr ) ;
	assign w_filter9_outputWave_datain = ( (|r_sys_processing_methodID) ? r_filter9_outputWave_datain : i_filter9_outputWave_datain ) ;
	assign o_filter9_outputWave_dataout = w_filter9_outputWave_dataout;
	assign w_filter9_outputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter9_outputWave_r_w : i_filter9_outputWave_r_w ) ;
	assign w_filter9_filterCoef_addr = ( (|r_sys_processing_methodID) ? r_filter9_filterCoef_addr : 9'sh0 ) ;
	assign w_filter9_filterCoef_datain = ( (|r_sys_processing_methodID) ? r_filter9_filterCoef_datain : 16'sh0 ) ;
	assign w_filter9_filterCoef_r_w = ( (|r_sys_processing_methodID) ? r_filter9_filterCoef_r_w : 1'h0 ) ;
	assign w_filter1_inputWave_addr = ( (|r_sys_processing_methodID) ? r_filter1_inputWave_addr : i_filter1_inputWave_addr ) ;
	assign w_filter1_inputWave_datain = ( (|r_sys_processing_methodID) ? r_filter1_inputWave_datain : i_filter1_inputWave_datain ) ;
	assign o_filter1_inputWave_dataout = w_filter1_inputWave_dataout;
	assign w_filter1_inputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter1_inputWave_r_w : i_filter1_inputWave_r_w ) ;
	assign w_filter1_outputWave_addr = ( (|r_sys_processing_methodID) ? r_filter1_outputWave_addr : i_filter1_outputWave_addr ) ;
	assign w_filter1_outputWave_datain = ( (|r_sys_processing_methodID) ? r_filter1_outputWave_datain : i_filter1_outputWave_datain ) ;
	assign o_filter1_outputWave_dataout = w_filter1_outputWave_dataout;
	assign w_filter1_outputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter1_outputWave_r_w : i_filter1_outputWave_r_w ) ;
	assign w_filter1_filterCoef_addr = ( (|r_sys_processing_methodID) ? r_filter1_filterCoef_addr : 9'sh0 ) ;
	assign w_filter1_filterCoef_datain = ( (|r_sys_processing_methodID) ? r_filter1_filterCoef_datain : 16'sh0 ) ;
	assign w_filter1_filterCoef_r_w = ( (|r_sys_processing_methodID) ? r_filter1_filterCoef_r_w : 1'h0 ) ;
	assign w_filter10_inputWave_addr = ( (|r_sys_processing_methodID) ? r_filter10_inputWave_addr : i_filter10_inputWave_addr ) ;
	assign w_filter10_inputWave_datain = ( (|r_sys_processing_methodID) ? r_filter10_inputWave_datain : i_filter10_inputWave_datain ) ;
	assign o_filter10_inputWave_dataout = w_filter10_inputWave_dataout;
	assign w_filter10_inputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter10_inputWave_r_w : i_filter10_inputWave_r_w ) ;
	assign w_filter10_outputWave_addr = ( (|r_sys_processing_methodID) ? r_filter10_outputWave_addr : i_filter10_outputWave_addr ) ;
	assign w_filter10_outputWave_datain = ( (|r_sys_processing_methodID) ? r_filter10_outputWave_datain : i_filter10_outputWave_datain ) ;
	assign o_filter10_outputWave_dataout = w_filter10_outputWave_dataout;
	assign w_filter10_outputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter10_outputWave_r_w : i_filter10_outputWave_r_w ) ;
	assign w_filter10_filterCoef_addr = ( (|r_sys_processing_methodID) ? r_filter10_filterCoef_addr : 9'sh0 ) ;
	assign w_filter10_filterCoef_datain = ( (|r_sys_processing_methodID) ? r_filter10_filterCoef_datain : 16'sh0 ) ;
	assign w_filter10_filterCoef_r_w = ( (|r_sys_processing_methodID) ? r_filter10_filterCoef_r_w : 1'h0 ) ;
	assign w_filter0_inputWave_addr = ( (|r_sys_processing_methodID) ? r_filter0_inputWave_addr : i_filter0_inputWave_addr ) ;
	assign w_filter0_inputWave_datain = ( (|r_sys_processing_methodID) ? r_filter0_inputWave_datain : i_filter0_inputWave_datain ) ;
	assign o_filter0_inputWave_dataout = w_filter0_inputWave_dataout;
	assign w_filter0_inputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter0_inputWave_r_w : i_filter0_inputWave_r_w ) ;
	assign w_filter0_outputWave_addr = ( (|r_sys_processing_methodID) ? r_filter0_outputWave_addr : i_filter0_outputWave_addr ) ;
	assign w_filter0_outputWave_datain = ( (|r_sys_processing_methodID) ? r_filter0_outputWave_datain : i_filter0_outputWave_datain ) ;
	assign o_filter0_outputWave_dataout = w_filter0_outputWave_dataout;
	assign w_filter0_outputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter0_outputWave_r_w : i_filter0_outputWave_r_w ) ;
	assign w_filter0_filterCoef_addr = ( (|r_sys_processing_methodID) ? r_filter0_filterCoef_addr : 9'sh0 ) ;
	assign w_filter0_filterCoef_datain = ( (|r_sys_processing_methodID) ? r_filter0_filterCoef_datain : 16'sh0 ) ;
	assign w_filter0_filterCoef_r_w = ( (|r_sys_processing_methodID) ? r_filter0_filterCoef_r_w : 1'h0 ) ;
	assign w_filter3_inputWave_addr = ( (|r_sys_processing_methodID) ? r_filter3_inputWave_addr : i_filter3_inputWave_addr ) ;
	assign w_filter3_inputWave_datain = ( (|r_sys_processing_methodID) ? r_filter3_inputWave_datain : i_filter3_inputWave_datain ) ;
	assign o_filter3_inputWave_dataout = w_filter3_inputWave_dataout;
	assign w_filter3_inputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter3_inputWave_r_w : i_filter3_inputWave_r_w ) ;
	assign w_filter3_outputWave_addr = ( (|r_sys_processing_methodID) ? r_filter3_outputWave_addr : i_filter3_outputWave_addr ) ;
	assign w_filter3_outputWave_datain = ( (|r_sys_processing_methodID) ? r_filter3_outputWave_datain : i_filter3_outputWave_datain ) ;
	assign o_filter3_outputWave_dataout = w_filter3_outputWave_dataout;
	assign w_filter3_outputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter3_outputWave_r_w : i_filter3_outputWave_r_w ) ;
	assign w_filter3_filterCoef_addr = ( (|r_sys_processing_methodID) ? r_filter3_filterCoef_addr : 9'sh0 ) ;
	assign w_filter3_filterCoef_datain = ( (|r_sys_processing_methodID) ? r_filter3_filterCoef_datain : 16'sh0 ) ;
	assign w_filter3_filterCoef_r_w = ( (|r_sys_processing_methodID) ? r_filter3_filterCoef_r_w : 1'h0 ) ;
	assign w_filter2_inputWave_addr = ( (|r_sys_processing_methodID) ? r_filter2_inputWave_addr : i_filter2_inputWave_addr ) ;
	assign w_filter2_inputWave_datain = ( (|r_sys_processing_methodID) ? r_filter2_inputWave_datain : i_filter2_inputWave_datain ) ;
	assign o_filter2_inputWave_dataout = w_filter2_inputWave_dataout;
	assign w_filter2_inputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter2_inputWave_r_w : i_filter2_inputWave_r_w ) ;
	assign w_filter2_outputWave_addr = ( (|r_sys_processing_methodID) ? r_filter2_outputWave_addr : i_filter2_outputWave_addr ) ;
	assign w_filter2_outputWave_datain = ( (|r_sys_processing_methodID) ? r_filter2_outputWave_datain : i_filter2_outputWave_datain ) ;
	assign o_filter2_outputWave_dataout = w_filter2_outputWave_dataout;
	assign w_filter2_outputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter2_outputWave_r_w : i_filter2_outputWave_r_w ) ;
	assign w_filter2_filterCoef_addr = ( (|r_sys_processing_methodID) ? r_filter2_filterCoef_addr : 9'sh0 ) ;
	assign w_filter2_filterCoef_datain = ( (|r_sys_processing_methodID) ? r_filter2_filterCoef_datain : 16'sh0 ) ;
	assign w_filter2_filterCoef_r_w = ( (|r_sys_processing_methodID) ? r_filter2_filterCoef_r_w : 1'h0 ) ;
	assign w_filter5_inputWave_addr = ( (|r_sys_processing_methodID) ? r_filter5_inputWave_addr : i_filter5_inputWave_addr ) ;
	assign w_filter5_inputWave_datain = ( (|r_sys_processing_methodID) ? r_filter5_inputWave_datain : i_filter5_inputWave_datain ) ;
	assign o_filter5_inputWave_dataout = w_filter5_inputWave_dataout;
	assign w_filter5_inputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter5_inputWave_r_w : i_filter5_inputWave_r_w ) ;
	assign w_filter5_outputWave_addr = ( (|r_sys_processing_methodID) ? r_filter5_outputWave_addr : i_filter5_outputWave_addr ) ;
	assign w_filter5_outputWave_datain = ( (|r_sys_processing_methodID) ? r_filter5_outputWave_datain : i_filter5_outputWave_datain ) ;
	assign o_filter5_outputWave_dataout = w_filter5_outputWave_dataout;
	assign w_filter5_outputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter5_outputWave_r_w : i_filter5_outputWave_r_w ) ;
	assign w_filter5_filterCoef_addr = ( (|r_sys_processing_methodID) ? r_filter5_filterCoef_addr : 9'sh0 ) ;
	assign w_filter5_filterCoef_datain = ( (|r_sys_processing_methodID) ? r_filter5_filterCoef_datain : 16'sh0 ) ;
	assign w_filter5_filterCoef_r_w = ( (|r_sys_processing_methodID) ? r_filter5_filterCoef_r_w : 1'h0 ) ;
	assign w_filter4_inputWave_addr = ( (|r_sys_processing_methodID) ? r_filter4_inputWave_addr : i_filter4_inputWave_addr ) ;
	assign w_filter4_inputWave_datain = ( (|r_sys_processing_methodID) ? r_filter4_inputWave_datain : i_filter4_inputWave_datain ) ;
	assign o_filter4_inputWave_dataout = w_filter4_inputWave_dataout;
	assign w_filter4_inputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter4_inputWave_r_w : i_filter4_inputWave_r_w ) ;
	assign w_filter4_outputWave_addr = ( (|r_sys_processing_methodID) ? r_filter4_outputWave_addr : i_filter4_outputWave_addr ) ;
	assign w_filter4_outputWave_datain = ( (|r_sys_processing_methodID) ? r_filter4_outputWave_datain : i_filter4_outputWave_datain ) ;
	assign o_filter4_outputWave_dataout = w_filter4_outputWave_dataout;
	assign w_filter4_outputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter4_outputWave_r_w : i_filter4_outputWave_r_w ) ;
	assign w_filter4_filterCoef_addr = ( (|r_sys_processing_methodID) ? r_filter4_filterCoef_addr : 9'sh0 ) ;
	assign w_filter4_filterCoef_datain = ( (|r_sys_processing_methodID) ? r_filter4_filterCoef_datain : 16'sh0 ) ;
	assign w_filter4_filterCoef_r_w = ( (|r_sys_processing_methodID) ? r_filter4_filterCoef_r_w : 1'h0 ) ;
	assign w_filter7_inputWave_addr = ( (|r_sys_processing_methodID) ? r_filter7_inputWave_addr : i_filter7_inputWave_addr ) ;
	assign w_filter7_inputWave_datain = ( (|r_sys_processing_methodID) ? r_filter7_inputWave_datain : i_filter7_inputWave_datain ) ;
	assign o_filter7_inputWave_dataout = w_filter7_inputWave_dataout;
	assign w_filter7_inputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter7_inputWave_r_w : i_filter7_inputWave_r_w ) ;
	assign w_filter7_outputWave_addr = ( (|r_sys_processing_methodID) ? r_filter7_outputWave_addr : i_filter7_outputWave_addr ) ;
	assign w_filter7_outputWave_datain = ( (|r_sys_processing_methodID) ? r_filter7_outputWave_datain : i_filter7_outputWave_datain ) ;
	assign o_filter7_outputWave_dataout = w_filter7_outputWave_dataout;
	assign w_filter7_outputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter7_outputWave_r_w : i_filter7_outputWave_r_w ) ;
	assign w_filter7_filterCoef_addr = ( (|r_sys_processing_methodID) ? r_filter7_filterCoef_addr : 9'sh0 ) ;
	assign w_filter7_filterCoef_datain = ( (|r_sys_processing_methodID) ? r_filter7_filterCoef_datain : 16'sh0 ) ;
	assign w_filter7_filterCoef_r_w = ( (|r_sys_processing_methodID) ? r_filter7_filterCoef_r_w : 1'h0 ) ;
	assign w_filter6_inputWave_addr = ( (|r_sys_processing_methodID) ? r_filter6_inputWave_addr : i_filter6_inputWave_addr ) ;
	assign w_filter6_inputWave_datain = ( (|r_sys_processing_methodID) ? r_filter6_inputWave_datain : i_filter6_inputWave_datain ) ;
	assign o_filter6_inputWave_dataout = w_filter6_inputWave_dataout;
	assign w_filter6_inputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter6_inputWave_r_w : i_filter6_inputWave_r_w ) ;
	assign w_filter6_outputWave_addr = ( (|r_sys_processing_methodID) ? r_filter6_outputWave_addr : i_filter6_outputWave_addr ) ;
	assign w_filter6_outputWave_datain = ( (|r_sys_processing_methodID) ? r_filter6_outputWave_datain : i_filter6_outputWave_datain ) ;
	assign o_filter6_outputWave_dataout = w_filter6_outputWave_dataout;
	assign w_filter6_outputWave_r_w = ( (|r_sys_processing_methodID) ? r_filter6_outputWave_r_w : i_filter6_outputWave_r_w ) ;
	assign w_filter6_filterCoef_addr = ( (|r_sys_processing_methodID) ? r_filter6_filterCoef_addr : 9'sh0 ) ;
	assign w_filter6_filterCoef_datain = ( (|r_sys_processing_methodID) ? r_filter6_filterCoef_datain : 16'sh0 ) ;
	assign w_filter6_filterCoef_r_w = ( (|r_sys_processing_methodID) ? r_filter6_filterCoef_r_w : 1'h0 ) ;


	FixedFilterThread
		filter15_inst(
			.i_fld_filterCoef_2_addr_0 (w_filter15_filterCoef_addr),
			.i_fld_filterCoef_2_datain_0 (w_filter15_filterCoef_datain),
			.o_fld_filterCoef_2_dataout_0 (w_filter15_filterCoef_dataout),
			.i_fld_filterCoef_2_r_w_0 (w_filter15_filterCoef_r_w),
			.i_fld_inputWave_0_addr_0 (w_filter15_inputWave_addr),
			.i_fld_inputWave_0_datain_0 (w_filter15_inputWave_datain),
			.o_fld_inputWave_0_dataout_0 (w_filter15_inputWave_dataout),
			.i_fld_inputWave_0_r_w_0 (w_filter15_inputWave_r_w),
			.i_fld_outputWave_1_addr_0 (w_filter15_outputWave_addr),
			.i_fld_outputWave_1_datain_0 (w_filter15_outputWave_datain),
			.o_fld_outputWave_1_dataout_0 (w_filter15_outputWave_dataout),
			.i_fld_outputWave_1_r_w_0 (w_filter15_outputWave_r_w),
			.o_run_busy (w_filter15_run_busy),
			.i_run_req (r_filter15_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	FixedFilterThread
		filter14_inst(
			.i_fld_filterCoef_2_addr_0 (w_filter14_filterCoef_addr),
			.i_fld_filterCoef_2_datain_0 (w_filter14_filterCoef_datain),
			.o_fld_filterCoef_2_dataout_0 (w_filter14_filterCoef_dataout),
			.i_fld_filterCoef_2_r_w_0 (w_filter14_filterCoef_r_w),
			.i_fld_inputWave_0_addr_0 (w_filter14_inputWave_addr),
			.i_fld_inputWave_0_datain_0 (w_filter14_inputWave_datain),
			.o_fld_inputWave_0_dataout_0 (w_filter14_inputWave_dataout),
			.i_fld_inputWave_0_r_w_0 (w_filter14_inputWave_r_w),
			.i_fld_outputWave_1_addr_0 (w_filter14_outputWave_addr),
			.i_fld_outputWave_1_datain_0 (w_filter14_outputWave_datain),
			.o_fld_outputWave_1_dataout_0 (w_filter14_outputWave_dataout),
			.i_fld_outputWave_1_r_w_0 (w_filter14_outputWave_r_w),
			.o_run_busy (w_filter14_run_busy),
			.i_run_req (r_filter14_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	FixedFilterThread
		filter13_inst(
			.i_fld_filterCoef_2_addr_0 (w_filter13_filterCoef_addr),
			.i_fld_filterCoef_2_datain_0 (w_filter13_filterCoef_datain),
			.o_fld_filterCoef_2_dataout_0 (w_filter13_filterCoef_dataout),
			.i_fld_filterCoef_2_r_w_0 (w_filter13_filterCoef_r_w),
			.i_fld_inputWave_0_addr_0 (w_filter13_inputWave_addr),
			.i_fld_inputWave_0_datain_0 (w_filter13_inputWave_datain),
			.o_fld_inputWave_0_dataout_0 (w_filter13_inputWave_dataout),
			.i_fld_inputWave_0_r_w_0 (w_filter13_inputWave_r_w),
			.i_fld_outputWave_1_addr_0 (w_filter13_outputWave_addr),
			.i_fld_outputWave_1_datain_0 (w_filter13_outputWave_datain),
			.o_fld_outputWave_1_dataout_0 (w_filter13_outputWave_dataout),
			.i_fld_outputWave_1_r_w_0 (w_filter13_outputWave_r_w),
			.o_run_busy (w_filter13_run_busy),
			.i_run_req (r_filter13_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	FixedFilterThread
		filter8_inst(
			.i_fld_filterCoef_2_addr_0 (w_filter8_filterCoef_addr),
			.i_fld_filterCoef_2_datain_0 (w_filter8_filterCoef_datain),
			.o_fld_filterCoef_2_dataout_0 (w_filter8_filterCoef_dataout),
			.i_fld_filterCoef_2_r_w_0 (w_filter8_filterCoef_r_w),
			.i_fld_inputWave_0_addr_0 (w_filter8_inputWave_addr),
			.i_fld_inputWave_0_datain_0 (w_filter8_inputWave_datain),
			.o_fld_inputWave_0_dataout_0 (w_filter8_inputWave_dataout),
			.i_fld_inputWave_0_r_w_0 (w_filter8_inputWave_r_w),
			.i_fld_outputWave_1_addr_0 (w_filter8_outputWave_addr),
			.i_fld_outputWave_1_datain_0 (w_filter8_outputWave_datain),
			.o_fld_outputWave_1_dataout_0 (w_filter8_outputWave_dataout),
			.i_fld_outputWave_1_r_w_0 (w_filter8_outputWave_r_w),
			.o_run_busy (w_filter8_run_busy),
			.i_run_req (r_filter8_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	FixedFilterThread
		filter12_inst(
			.i_fld_filterCoef_2_addr_0 (w_filter12_filterCoef_addr),
			.i_fld_filterCoef_2_datain_0 (w_filter12_filterCoef_datain),
			.o_fld_filterCoef_2_dataout_0 (w_filter12_filterCoef_dataout),
			.i_fld_filterCoef_2_r_w_0 (w_filter12_filterCoef_r_w),
			.i_fld_inputWave_0_addr_0 (w_filter12_inputWave_addr),
			.i_fld_inputWave_0_datain_0 (w_filter12_inputWave_datain),
			.o_fld_inputWave_0_dataout_0 (w_filter12_inputWave_dataout),
			.i_fld_inputWave_0_r_w_0 (w_filter12_inputWave_r_w),
			.i_fld_outputWave_1_addr_0 (w_filter12_outputWave_addr),
			.i_fld_outputWave_1_datain_0 (w_filter12_outputWave_datain),
			.o_fld_outputWave_1_dataout_0 (w_filter12_outputWave_dataout),
			.i_fld_outputWave_1_r_w_0 (w_filter12_outputWave_r_w),
			.o_run_busy (w_filter12_run_busy),
			.i_run_req (r_filter12_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	FixedFilterThread
		filter11_inst(
			.i_fld_filterCoef_2_addr_0 (w_filter11_filterCoef_addr),
			.i_fld_filterCoef_2_datain_0 (w_filter11_filterCoef_datain),
			.o_fld_filterCoef_2_dataout_0 (w_filter11_filterCoef_dataout),
			.i_fld_filterCoef_2_r_w_0 (w_filter11_filterCoef_r_w),
			.i_fld_inputWave_0_addr_0 (w_filter11_inputWave_addr),
			.i_fld_inputWave_0_datain_0 (w_filter11_inputWave_datain),
			.o_fld_inputWave_0_dataout_0 (w_filter11_inputWave_dataout),
			.i_fld_inputWave_0_r_w_0 (w_filter11_inputWave_r_w),
			.i_fld_outputWave_1_addr_0 (w_filter11_outputWave_addr),
			.i_fld_outputWave_1_datain_0 (w_filter11_outputWave_datain),
			.o_fld_outputWave_1_dataout_0 (w_filter11_outputWave_dataout),
			.i_fld_outputWave_1_r_w_0 (w_filter11_outputWave_r_w),
			.o_run_busy (w_filter11_run_busy),
			.i_run_req (r_filter11_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	FixedFilterThread
		filter9_inst(
			.i_fld_filterCoef_2_addr_0 (w_filter9_filterCoef_addr),
			.i_fld_filterCoef_2_datain_0 (w_filter9_filterCoef_datain),
			.o_fld_filterCoef_2_dataout_0 (w_filter9_filterCoef_dataout),
			.i_fld_filterCoef_2_r_w_0 (w_filter9_filterCoef_r_w),
			.i_fld_inputWave_0_addr_0 (w_filter9_inputWave_addr),
			.i_fld_inputWave_0_datain_0 (w_filter9_inputWave_datain),
			.o_fld_inputWave_0_dataout_0 (w_filter9_inputWave_dataout),
			.i_fld_inputWave_0_r_w_0 (w_filter9_inputWave_r_w),
			.i_fld_outputWave_1_addr_0 (w_filter9_outputWave_addr),
			.i_fld_outputWave_1_datain_0 (w_filter9_outputWave_datain),
			.o_fld_outputWave_1_dataout_0 (w_filter9_outputWave_dataout),
			.i_fld_outputWave_1_r_w_0 (w_filter9_outputWave_r_w),
			.o_run_busy (w_filter9_run_busy),
			.i_run_req (r_filter9_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	FixedFilterThread
		filter1_inst(
			.i_fld_filterCoef_2_addr_0 (w_filter1_filterCoef_addr),
			.i_fld_filterCoef_2_datain_0 (w_filter1_filterCoef_datain),
			.o_fld_filterCoef_2_dataout_0 (w_filter1_filterCoef_dataout),
			.i_fld_filterCoef_2_r_w_0 (w_filter1_filterCoef_r_w),
			.i_fld_inputWave_0_addr_0 (w_filter1_inputWave_addr),
			.i_fld_inputWave_0_datain_0 (w_filter1_inputWave_datain),
			.o_fld_inputWave_0_dataout_0 (w_filter1_inputWave_dataout),
			.i_fld_inputWave_0_r_w_0 (w_filter1_inputWave_r_w),
			.i_fld_outputWave_1_addr_0 (w_filter1_outputWave_addr),
			.i_fld_outputWave_1_datain_0 (w_filter1_outputWave_datain),
			.o_fld_outputWave_1_dataout_0 (w_filter1_outputWave_dataout),
			.i_fld_outputWave_1_r_w_0 (w_filter1_outputWave_r_w),
			.o_run_busy (w_filter1_run_busy),
			.i_run_req (r_filter1_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	FixedFilterThread
		filter10_inst(
			.i_fld_filterCoef_2_addr_0 (w_filter10_filterCoef_addr),
			.i_fld_filterCoef_2_datain_0 (w_filter10_filterCoef_datain),
			.o_fld_filterCoef_2_dataout_0 (w_filter10_filterCoef_dataout),
			.i_fld_filterCoef_2_r_w_0 (w_filter10_filterCoef_r_w),
			.i_fld_inputWave_0_addr_0 (w_filter10_inputWave_addr),
			.i_fld_inputWave_0_datain_0 (w_filter10_inputWave_datain),
			.o_fld_inputWave_0_dataout_0 (w_filter10_inputWave_dataout),
			.i_fld_inputWave_0_r_w_0 (w_filter10_inputWave_r_w),
			.i_fld_outputWave_1_addr_0 (w_filter10_outputWave_addr),
			.i_fld_outputWave_1_datain_0 (w_filter10_outputWave_datain),
			.o_fld_outputWave_1_dataout_0 (w_filter10_outputWave_dataout),
			.i_fld_outputWave_1_r_w_0 (w_filter10_outputWave_r_w),
			.o_run_busy (w_filter10_run_busy),
			.i_run_req (r_filter10_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	FixedFilterThread
		filter0_inst(
			.i_fld_filterCoef_2_addr_0 (w_filter0_filterCoef_addr),
			.i_fld_filterCoef_2_datain_0 (w_filter0_filterCoef_datain),
			.o_fld_filterCoef_2_dataout_0 (w_filter0_filterCoef_dataout),
			.i_fld_filterCoef_2_r_w_0 (w_filter0_filterCoef_r_w),
			.i_fld_inputWave_0_addr_0 (w_filter0_inputWave_addr),
			.i_fld_inputWave_0_datain_0 (w_filter0_inputWave_datain),
			.o_fld_inputWave_0_dataout_0 (w_filter0_inputWave_dataout),
			.i_fld_inputWave_0_r_w_0 (w_filter0_inputWave_r_w),
			.i_fld_outputWave_1_addr_0 (w_filter0_outputWave_addr),
			.i_fld_outputWave_1_datain_0 (w_filter0_outputWave_datain),
			.o_fld_outputWave_1_dataout_0 (w_filter0_outputWave_dataout),
			.i_fld_outputWave_1_r_w_0 (w_filter0_outputWave_r_w),
			.o_run_busy (w_filter0_run_busy),
			.i_run_req (r_filter0_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	FixedFilterThread
		filter3_inst(
			.i_fld_filterCoef_2_addr_0 (w_filter3_filterCoef_addr),
			.i_fld_filterCoef_2_datain_0 (w_filter3_filterCoef_datain),
			.o_fld_filterCoef_2_dataout_0 (w_filter3_filterCoef_dataout),
			.i_fld_filterCoef_2_r_w_0 (w_filter3_filterCoef_r_w),
			.i_fld_inputWave_0_addr_0 (w_filter3_inputWave_addr),
			.i_fld_inputWave_0_datain_0 (w_filter3_inputWave_datain),
			.o_fld_inputWave_0_dataout_0 (w_filter3_inputWave_dataout),
			.i_fld_inputWave_0_r_w_0 (w_filter3_inputWave_r_w),
			.i_fld_outputWave_1_addr_0 (w_filter3_outputWave_addr),
			.i_fld_outputWave_1_datain_0 (w_filter3_outputWave_datain),
			.o_fld_outputWave_1_dataout_0 (w_filter3_outputWave_dataout),
			.i_fld_outputWave_1_r_w_0 (w_filter3_outputWave_r_w),
			.o_run_busy (w_filter3_run_busy),
			.i_run_req (r_filter3_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	FixedFilterThread
		filter2_inst(
			.i_fld_filterCoef_2_addr_0 (w_filter2_filterCoef_addr),
			.i_fld_filterCoef_2_datain_0 (w_filter2_filterCoef_datain),
			.o_fld_filterCoef_2_dataout_0 (w_filter2_filterCoef_dataout),
			.i_fld_filterCoef_2_r_w_0 (w_filter2_filterCoef_r_w),
			.i_fld_inputWave_0_addr_0 (w_filter2_inputWave_addr),
			.i_fld_inputWave_0_datain_0 (w_filter2_inputWave_datain),
			.o_fld_inputWave_0_dataout_0 (w_filter2_inputWave_dataout),
			.i_fld_inputWave_0_r_w_0 (w_filter2_inputWave_r_w),
			.i_fld_outputWave_1_addr_0 (w_filter2_outputWave_addr),
			.i_fld_outputWave_1_datain_0 (w_filter2_outputWave_datain),
			.o_fld_outputWave_1_dataout_0 (w_filter2_outputWave_dataout),
			.i_fld_outputWave_1_r_w_0 (w_filter2_outputWave_r_w),
			.o_run_busy (w_filter2_run_busy),
			.i_run_req (r_filter2_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	FixedFilterThread
		filter5_inst(
			.i_fld_filterCoef_2_addr_0 (w_filter5_filterCoef_addr),
			.i_fld_filterCoef_2_datain_0 (w_filter5_filterCoef_datain),
			.o_fld_filterCoef_2_dataout_0 (w_filter5_filterCoef_dataout),
			.i_fld_filterCoef_2_r_w_0 (w_filter5_filterCoef_r_w),
			.i_fld_inputWave_0_addr_0 (w_filter5_inputWave_addr),
			.i_fld_inputWave_0_datain_0 (w_filter5_inputWave_datain),
			.o_fld_inputWave_0_dataout_0 (w_filter5_inputWave_dataout),
			.i_fld_inputWave_0_r_w_0 (w_filter5_inputWave_r_w),
			.i_fld_outputWave_1_addr_0 (w_filter5_outputWave_addr),
			.i_fld_outputWave_1_datain_0 (w_filter5_outputWave_datain),
			.o_fld_outputWave_1_dataout_0 (w_filter5_outputWave_dataout),
			.i_fld_outputWave_1_r_w_0 (w_filter5_outputWave_r_w),
			.o_run_busy (w_filter5_run_busy),
			.i_run_req (r_filter5_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	FixedFilterThread
		filter4_inst(
			.i_fld_filterCoef_2_addr_0 (w_filter4_filterCoef_addr),
			.i_fld_filterCoef_2_datain_0 (w_filter4_filterCoef_datain),
			.o_fld_filterCoef_2_dataout_0 (w_filter4_filterCoef_dataout),
			.i_fld_filterCoef_2_r_w_0 (w_filter4_filterCoef_r_w),
			.i_fld_inputWave_0_addr_0 (w_filter4_inputWave_addr),
			.i_fld_inputWave_0_datain_0 (w_filter4_inputWave_datain),
			.o_fld_inputWave_0_dataout_0 (w_filter4_inputWave_dataout),
			.i_fld_inputWave_0_r_w_0 (w_filter4_inputWave_r_w),
			.i_fld_outputWave_1_addr_0 (w_filter4_outputWave_addr),
			.i_fld_outputWave_1_datain_0 (w_filter4_outputWave_datain),
			.o_fld_outputWave_1_dataout_0 (w_filter4_outputWave_dataout),
			.i_fld_outputWave_1_r_w_0 (w_filter4_outputWave_r_w),
			.o_run_busy (w_filter4_run_busy),
			.i_run_req (r_filter4_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	FixedFilterThread
		filter7_inst(
			.i_fld_filterCoef_2_addr_0 (w_filter7_filterCoef_addr),
			.i_fld_filterCoef_2_datain_0 (w_filter7_filterCoef_datain),
			.o_fld_filterCoef_2_dataout_0 (w_filter7_filterCoef_dataout),
			.i_fld_filterCoef_2_r_w_0 (w_filter7_filterCoef_r_w),
			.i_fld_inputWave_0_addr_0 (w_filter7_inputWave_addr),
			.i_fld_inputWave_0_datain_0 (w_filter7_inputWave_datain),
			.o_fld_inputWave_0_dataout_0 (w_filter7_inputWave_dataout),
			.i_fld_inputWave_0_r_w_0 (w_filter7_inputWave_r_w),
			.i_fld_outputWave_1_addr_0 (w_filter7_outputWave_addr),
			.i_fld_outputWave_1_datain_0 (w_filter7_outputWave_datain),
			.o_fld_outputWave_1_dataout_0 (w_filter7_outputWave_dataout),
			.i_fld_outputWave_1_r_w_0 (w_filter7_outputWave_r_w),
			.o_run_busy (w_filter7_run_busy),
			.i_run_req (r_filter7_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	FixedFilterThread
		filter6_inst(
			.i_fld_filterCoef_2_addr_0 (w_filter6_filterCoef_addr),
			.i_fld_filterCoef_2_datain_0 (w_filter6_filterCoef_datain),
			.o_fld_filterCoef_2_dataout_0 (w_filter6_filterCoef_dataout),
			.i_fld_filterCoef_2_r_w_0 (w_filter6_filterCoef_r_w),
			.i_fld_inputWave_0_addr_0 (w_filter6_inputWave_addr),
			.i_fld_inputWave_0_datain_0 (w_filter6_inputWave_datain),
			.o_fld_inputWave_0_dataout_0 (w_filter6_inputWave_dataout),
			.i_fld_inputWave_0_r_w_0 (w_filter6_inputWave_r_w),
			.i_fld_outputWave_1_addr_0 (w_filter6_outputWave_addr),
			.i_fld_outputWave_1_datain_0 (w_filter6_outputWave_datain),
			.o_fld_outputWave_1_dataout_0 (w_filter6_outputWave_dataout),
			.i_fld_outputWave_1_r_w_0 (w_filter6_outputWave_r_w),
			.o_run_busy (w_filter6_run_busy),
			.i_run_req (r_filter6_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_main_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_main_phase) 
						3'h6: begin
							r_sys_processing_methodID <= r_sys_main_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_main_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_main_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_main_phase <= 3'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h0: begin
							r_sys_main_phase <= 3'h2;
						end

						3'h2: begin

							case(r_sys_main_stage) 
								5'hf: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_phase <= 3'h4;

									end
								end

							endcase
						end

						3'h4: begin

							case(r_sys_main_stage) 
								5'hf: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_phase <= 3'h6;

									end
								end

							endcase
						end

						3'h6: begin
							r_sys_main_phase <= 3'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_main_stage <= 5'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= 5'h0;

									end
								end

							endcase
						end

						3'h4: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= w_sys_main_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_stage <= 5'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_main_step <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
									else
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= w_sys_main_step_p1;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
									else
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= w_sys_main_step_p1;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= w_sys_main_step_p1;

									end
									else
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
									else
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= w_sys_main_step_p1;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
									else
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= w_sys_main_step_p1;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= w_sys_main_step_p1;

									end
									else
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
									else
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= w_sys_main_step_p1;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= w_sys_main_step_p1;

									end
									else
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
									else
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= w_sys_main_step_p1;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
									else
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= w_sys_main_step_p1;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
									else
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= w_sys_main_step_p1;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= w_sys_main_step_p1;

									end
									else
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= w_sys_main_step_p1;

									end
									else
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
									else
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= w_sys_main_step_p1;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
									else
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= w_sys_main_step_p1;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
									else
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= w_sys_main_step_p1;

									end
								end

							endcase
						end

						3'h4: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= ((w_filter0_run_busy) ? r_sys_main_step : w_sys_main_step_p1);

									end
									else
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
									else
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= ((w_filter1_run_busy) ? r_sys_main_step : w_sys_main_step_p1);

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= ((w_filter2_run_busy) ? r_sys_main_step : w_sys_main_step_p1);

									end
									else
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= ((w_filter3_run_busy) ? r_sys_main_step : w_sys_main_step_p1);

									end
									else
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
									else
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= ((w_filter4_run_busy) ? r_sys_main_step : w_sys_main_step_p1);

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
									else
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= ((w_filter5_run_busy) ? r_sys_main_step : w_sys_main_step_p1);

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= ((w_filter6_run_busy) ? r_sys_main_step : w_sys_main_step_p1);

									end
									else
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
									else
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= ((w_filter7_run_busy) ? r_sys_main_step : w_sys_main_step_p1);

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
									else
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= ((w_filter8_run_busy) ? r_sys_main_step : w_sys_main_step_p1);

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
									else
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= ((w_filter9_run_busy) ? r_sys_main_step : w_sys_main_step_p1);

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
									else
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= ((w_filter10_run_busy) ? r_sys_main_step : w_sys_main_step_p1);

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
									else
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= ((w_filter11_run_busy) ? r_sys_main_step : w_sys_main_step_p1);

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
									else
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= ((w_filter12_run_busy) ? r_sys_main_step : w_sys_main_step_p1);

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
									else
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= ((w_filter13_run_busy) ? r_sys_main_step : w_sys_main_step_p1);

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
									else
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= ((w_filter14_run_busy) ? r_sys_main_step : w_sys_main_step_p1);

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_sys_main_step <= ((w_filter15_run_busy) ? r_sys_main_step : w_sys_main_step_p1);

									end
									else
									if((r_sys_main_step==2'h1)) begin
										r_sys_main_step <= 2'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_main_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_main_busy <= ((i_main_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_main_phase) 
						3'h0: begin
							r_sys_main_busy <= w_sys_boolTrue;
						end

						3'h6: begin
							r_sys_main_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter15_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_main_step==2'h1)) begin
										r_filter15_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter15_inputWave_addr <= 12'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter15_inputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_inputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter15_inputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter15_outputWave_addr <= 11'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter15_outputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_outputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter15_outputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter15_filterCoef_addr <= 9'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter15_filterCoef_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter15_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter15_filterCoef_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter14_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_main_step==2'h1)) begin
										r_filter14_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter14_inputWave_addr <= 12'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter14_inputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_inputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter14_inputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter14_outputWave_addr <= 11'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter14_outputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_outputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter14_outputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter14_filterCoef_addr <= 9'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter14_filterCoef_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter14_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter14_filterCoef_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter13_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_main_step==2'h1)) begin
										r_filter13_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter13_inputWave_addr <= 12'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter13_inputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_inputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter13_inputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter13_outputWave_addr <= 11'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter13_outputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_outputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter13_outputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter13_filterCoef_addr <= 9'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter13_filterCoef_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter13_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter13_filterCoef_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter8_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_main_step==2'h1)) begin
										r_filter8_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter8_inputWave_addr <= 12'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter8_inputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_inputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter8_inputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter8_outputWave_addr <= 11'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter8_outputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_outputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter8_outputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter8_filterCoef_addr <= 9'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter8_filterCoef_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter8_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter8_filterCoef_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter12_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_main_step==2'h1)) begin
										r_filter12_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter12_inputWave_addr <= 12'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter12_inputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_inputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter12_inputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter12_outputWave_addr <= 11'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter12_outputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_outputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter12_outputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter12_filterCoef_addr <= 9'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter12_filterCoef_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter12_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter12_filterCoef_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter11_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_main_step==2'h1)) begin
										r_filter11_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter11_inputWave_addr <= 12'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter11_inputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_inputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter11_inputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter11_outputWave_addr <= 11'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter11_outputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_outputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter11_outputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter11_filterCoef_addr <= 9'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter11_filterCoef_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter11_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter11_filterCoef_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter9_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_main_step==2'h1)) begin
										r_filter9_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter9_inputWave_addr <= 12'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter9_inputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_inputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter9_inputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter9_outputWave_addr <= 11'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter9_outputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_outputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter9_outputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter9_filterCoef_addr <= 9'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter9_filterCoef_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter9_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter9_filterCoef_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter1_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_main_step==2'h1)) begin
										r_filter1_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter1_inputWave_addr <= 12'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter1_inputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_inputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter1_inputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter1_outputWave_addr <= 11'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter1_outputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_outputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter1_outputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter1_filterCoef_addr <= 9'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter1_filterCoef_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter1_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter1_filterCoef_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter10_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_main_step==2'h1)) begin
										r_filter10_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter10_inputWave_addr <= 12'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter10_inputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_inputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter10_inputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter10_outputWave_addr <= 11'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter10_outputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_outputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter10_outputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter10_filterCoef_addr <= 9'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter10_filterCoef_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter10_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter10_filterCoef_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter0_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_main_step==2'h1)) begin
										r_filter0_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter0_inputWave_addr <= 12'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter0_inputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_inputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter0_inputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter0_outputWave_addr <= 11'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter0_outputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_outputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter0_outputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter0_filterCoef_addr <= 9'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter0_filterCoef_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter0_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter0_filterCoef_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter3_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_main_step==2'h1)) begin
										r_filter3_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter3_inputWave_addr <= 12'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter3_inputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_inputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter3_inputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter3_outputWave_addr <= 11'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter3_outputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_outputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter3_outputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter3_filterCoef_addr <= 9'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter3_filterCoef_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter3_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter3_filterCoef_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter2_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_main_step==2'h1)) begin
										r_filter2_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter2_inputWave_addr <= 12'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter2_inputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_inputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter2_inputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter2_outputWave_addr <= 11'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter2_outputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_outputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter2_outputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter2_filterCoef_addr <= 9'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter2_filterCoef_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter2_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter2_filterCoef_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter5_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_main_step==2'h1)) begin
										r_filter5_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter5_inputWave_addr <= 12'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter5_inputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_inputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter5_inputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter5_outputWave_addr <= 11'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter5_outputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_outputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter5_outputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter5_filterCoef_addr <= 9'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter5_filterCoef_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter5_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter5_filterCoef_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter4_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_main_step==2'h1)) begin
										r_filter4_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter4_inputWave_addr <= 12'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter4_inputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_inputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter4_inputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter4_outputWave_addr <= 11'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter4_outputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_outputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter4_outputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter4_filterCoef_addr <= 9'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter4_filterCoef_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter4_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter4_filterCoef_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter7_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_main_step==2'h1)) begin
										r_filter7_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter7_inputWave_addr <= 12'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter7_inputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_inputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter7_inputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter7_outputWave_addr <= 11'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter7_outputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_outputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter7_outputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter7_filterCoef_addr <= 9'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter7_filterCoef_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter7_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter7_filterCoef_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter6_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_main_step==2'h1)) begin
										r_filter6_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter6_inputWave_addr <= 12'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter6_inputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_inputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_inputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter6_inputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter6_outputWave_addr <= 11'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter6_outputWave_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_outputWave_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_outputWave_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter6_outputWave_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter6_filterCoef_addr <= 9'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_filter6_filterCoef_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_main_phase) 
						3'h2: begin

							case(r_sys_main_stage) 
								5'h0: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_main_step==2'h0)) begin
										r_filter6_filterCoef_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_filter6_filterCoef_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


endmodule
