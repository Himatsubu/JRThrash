/*
TimeStamp:	2016/6/26		16:26
*/


module c1(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy	
);

	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 5:0] r_sys_run_phase;
	reg         [ 3:0] r_sys_run_stage;
	reg         [ 6:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 3:0] w_sys_run_stage_p1;
	wire        [ 6:0] w_sys_run_step_p1;
	wire signed [ 8:0] w_fld_u_0_addr_0;
	wire        [31:0] w_fld_u_0_datain_0;
	wire        [31:0] w_fld_u_0_dataout_0;
	wire               w_fld_u_0_r_w_0;
	wire               w_fld_u_0_ce_0;
	reg  signed [ 8:0] r_fld_u_0_addr_1;
	reg         [31:0] r_fld_u_0_datain_1;
	wire        [31:0] w_fld_u_0_dataout_1;
	reg                r_fld_u_0_r_w_1;
	wire               w_fld_u_0_ce_1;
	wire signed [ 8:0] w_fld_uu_1_addr_0;
	wire        [31:0] w_fld_uu_1_datain_0;
	wire        [31:0] w_fld_uu_1_dataout_0;
	wire               w_fld_uu_1_r_w_0;
	wire               w_fld_uu_1_ce_0;
	reg  signed [ 8:0] r_fld_uu_1_addr_1;
	reg         [31:0] r_fld_uu_1_datain_1;
	wire        [31:0] w_fld_uu_1_dataout_1;
	reg                r_fld_uu_1_r_w_1;
	wire               w_fld_uu_1_ce_1;
	reg  signed [31:0] r_run_k_11;
	reg  signed [31:0] r_run_j_12;
	reg  signed [31:0] r_run_n_13;
	reg  signed [31:0] r_run_mx_14;
	reg  signed [31:0] r_run_my_15;
	reg  signed [31:0] r_run_nlast_16;
	reg  signed [31:0] r_run_copy0_j_17;
	reg  signed [31:0] r_run_copy0_j_18;
	reg  signed [31:0] r_run_copy1_j_19;
	reg  signed [31:0] r_run_copy2_j_20;
	reg                r_sub08_run_req;
	wire               w_sub08_run_busy;
	wire signed [ 9:0] w_sub08_u_addr;
	reg  signed [ 9:0] r_sub08_u_addr;
	wire        [31:0] w_sub08_u_datain;
	reg         [31:0] r_sub08_u_datain;
	wire        [31:0] w_sub08_u_dataout;
	wire               w_sub08_u_r_w;
	reg                r_sub08_u_r_w;
	wire signed [ 9:0] w_sub08_result_addr;
	reg  signed [ 9:0] r_sub08_result_addr;
	wire        [31:0] w_sub08_result_datain;
	reg         [31:0] r_sub08_result_datain;
	wire        [31:0] w_sub08_result_dataout;
	wire               w_sub08_result_r_w;
	reg                r_sub08_result_r_w;
	reg                r_sub03_run_req;
	wire               w_sub03_run_busy;
	wire signed [ 9:0] w_sub03_u_addr;
	reg  signed [ 9:0] r_sub03_u_addr;
	wire        [31:0] w_sub03_u_datain;
	reg         [31:0] r_sub03_u_datain;
	wire        [31:0] w_sub03_u_dataout;
	wire               w_sub03_u_r_w;
	reg                r_sub03_u_r_w;
	wire signed [ 9:0] w_sub03_result_addr;
	reg  signed [ 9:0] r_sub03_result_addr;
	wire        [31:0] w_sub03_result_datain;
	reg         [31:0] r_sub03_result_datain;
	wire        [31:0] w_sub03_result_dataout;
	wire               w_sub03_result_r_w;
	reg                r_sub03_result_r_w;
	reg                r_sub02_run_req;
	wire               w_sub02_run_busy;
	wire signed [ 9:0] w_sub02_u_addr;
	reg  signed [ 9:0] r_sub02_u_addr;
	wire        [31:0] w_sub02_u_datain;
	reg         [31:0] r_sub02_u_datain;
	wire        [31:0] w_sub02_u_dataout;
	wire               w_sub02_u_r_w;
	reg                r_sub02_u_r_w;
	wire signed [ 9:0] w_sub02_result_addr;
	reg  signed [ 9:0] r_sub02_result_addr;
	wire        [31:0] w_sub02_result_datain;
	reg         [31:0] r_sub02_result_datain;
	wire        [31:0] w_sub02_result_dataout;
	wire               w_sub02_result_r_w;
	reg                r_sub02_result_r_w;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [ 9:0] w_sub01_u_addr;
	reg  signed [ 9:0] r_sub01_u_addr;
	wire        [31:0] w_sub01_u_datain;
	reg         [31:0] r_sub01_u_datain;
	wire        [31:0] w_sub01_u_dataout;
	wire               w_sub01_u_r_w;
	reg                r_sub01_u_r_w;
	wire signed [ 9:0] w_sub01_result_addr;
	reg  signed [ 9:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [ 9:0] w_sub00_u_addr;
	reg  signed [ 9:0] r_sub00_u_addr;
	wire        [31:0] w_sub00_u_datain;
	reg         [31:0] r_sub00_u_datain;
	wire        [31:0] w_sub00_u_dataout;
	wire               w_sub00_u_r_w;
	reg                r_sub00_u_r_w;
	wire signed [ 9:0] w_sub00_result_addr;
	reg  signed [ 9:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	reg                r_sub07_run_req;
	wire               w_sub07_run_busy;
	wire signed [ 9:0] w_sub07_u_addr;
	reg  signed [ 9:0] r_sub07_u_addr;
	wire        [31:0] w_sub07_u_datain;
	reg         [31:0] r_sub07_u_datain;
	wire        [31:0] w_sub07_u_dataout;
	wire               w_sub07_u_r_w;
	reg                r_sub07_u_r_w;
	wire signed [ 9:0] w_sub07_result_addr;
	reg  signed [ 9:0] r_sub07_result_addr;
	wire        [31:0] w_sub07_result_datain;
	reg         [31:0] r_sub07_result_datain;
	wire        [31:0] w_sub07_result_dataout;
	wire               w_sub07_result_r_w;
	reg                r_sub07_result_r_w;
	reg                r_sub06_run_req;
	wire               w_sub06_run_busy;
	wire signed [ 9:0] w_sub06_u_addr;
	reg  signed [ 9:0] r_sub06_u_addr;
	wire        [31:0] w_sub06_u_datain;
	reg         [31:0] r_sub06_u_datain;
	wire        [31:0] w_sub06_u_dataout;
	wire               w_sub06_u_r_w;
	reg                r_sub06_u_r_w;
	wire signed [ 9:0] w_sub06_result_addr;
	reg  signed [ 9:0] r_sub06_result_addr;
	wire        [31:0] w_sub06_result_datain;
	reg         [31:0] r_sub06_result_datain;
	wire        [31:0] w_sub06_result_dataout;
	wire               w_sub06_result_r_w;
	reg                r_sub06_result_r_w;
	reg                r_sub05_run_req;
	wire               w_sub05_run_busy;
	wire signed [ 9:0] w_sub05_u_addr;
	reg  signed [ 9:0] r_sub05_u_addr;
	wire        [31:0] w_sub05_u_datain;
	reg         [31:0] r_sub05_u_datain;
	wire        [31:0] w_sub05_u_dataout;
	wire               w_sub05_u_r_w;
	reg                r_sub05_u_r_w;
	wire signed [ 9:0] w_sub05_result_addr;
	reg  signed [ 9:0] r_sub05_result_addr;
	wire        [31:0] w_sub05_result_datain;
	reg         [31:0] r_sub05_result_datain;
	wire        [31:0] w_sub05_result_dataout;
	wire               w_sub05_result_r_w;
	reg                r_sub05_result_r_w;
	reg                r_sub04_run_req;
	wire               w_sub04_run_busy;
	wire signed [ 9:0] w_sub04_u_addr;
	reg  signed [ 9:0] r_sub04_u_addr;
	wire        [31:0] w_sub04_u_datain;
	reg         [31:0] r_sub04_u_datain;
	wire        [31:0] w_sub04_u_dataout;
	wire               w_sub04_u_r_w;
	reg                r_sub04_u_r_w;
	wire signed [ 9:0] w_sub04_result_addr;
	reg  signed [ 9:0] r_sub04_result_addr;
	wire        [31:0] w_sub04_result_datain;
	reg         [31:0] r_sub04_result_datain;
	wire        [31:0] w_sub04_result_dataout;
	wire               w_sub04_result_r_w;
	reg                r_sub04_result_r_w;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg         [31:0] r_sys_tmp4_float;
	reg         [31:0] r_sys_tmp5_float;
	reg         [31:0] r_sys_tmp6_float;
	reg         [31:0] r_sys_tmp7_float;
	reg         [31:0] r_sys_tmp8_float;
	reg         [31:0] r_sys_tmp9_float;
	reg         [31:0] r_sys_tmp10_float;
	reg         [31:0] r_sys_tmp11_float;
	reg         [31:0] r_sys_tmp12_float;
	reg         [31:0] r_sys_tmp13_float;
	reg         [31:0] r_sys_tmp14_float;
	reg         [31:0] r_sys_tmp15_float;
	reg         [31:0] r_sys_tmp16_float;
	reg         [31:0] r_sys_tmp17_float;
	reg         [31:0] r_sys_tmp18_float;
	reg         [31:0] r_sys_tmp19_float;
	reg         [31:0] r_sys_tmp20_float;
	reg         [31:0] r_sys_tmp21_float;
	reg         [31:0] r_sys_tmp22_float;
	reg         [31:0] r_sys_tmp23_float;
	reg         [31:0] r_sys_tmp24_float;
	reg         [31:0] r_sys_tmp25_float;
	reg         [31:0] r_sys_tmp26_float;
	reg         [31:0] r_sys_tmp27_float;
	reg         [31:0] r_sys_tmp28_float;
	reg         [31:0] r_sys_tmp29_float;
	reg         [31:0] r_sys_tmp30_float;
	reg         [31:0] r_sys_tmp31_float;
	reg         [31:0] r_sys_tmp32_float;
	reg         [31:0] r_sys_tmp33_float;
	reg         [31:0] r_sys_tmp34_float;
	reg         [31:0] r_sys_tmp35_float;
	reg         [31:0] r_sys_tmp36_float;
	reg         [31:0] r_sys_tmp37_float;
	reg         [31:0] r_sys_tmp38_float;
	reg         [31:0] r_sys_tmp39_float;
	reg         [31:0] r_sys_tmp40_float;
	reg         [31:0] r_sys_tmp41_float;
	reg         [31:0] r_sys_tmp42_float;
	reg         [31:0] r_sys_tmp43_float;
	reg         [31:0] r_sys_tmp44_float;
	reg         [31:0] r_sys_tmp45_float;
	reg         [31:0] r_sys_tmp46_float;
	reg         [31:0] r_sys_tmp47_float;
	wire signed [31:0] w_sys_tmp1;
	wire signed [31:0] w_sys_tmp3;
	wire               w_sys_tmp4;
	wire               w_sys_tmp5;
	wire signed [31:0] w_sys_tmp6;
	wire               w_sys_tmp7;
	wire               w_sys_tmp8;
	wire signed [31:0] w_sys_tmp11;
	wire signed [31:0] w_sys_tmp12;
	wire signed [31:0] w_sys_tmp13;
	wire        [31:0] w_sys_tmp14;
	wire signed [31:0] w_sys_tmp16;
	wire signed [31:0] w_sys_tmp17;
	wire signed [31:0] w_sys_tmp20;
	wire signed [31:0] w_sys_tmp21;
	wire               w_sys_tmp94;
	wire               w_sys_tmp95;
	wire signed [31:0] w_sys_tmp96;
	wire               w_sys_tmp97;
	wire               w_sys_tmp98;
	wire signed [31:0] w_sys_tmp101;
	wire signed [31:0] w_sys_tmp102;
	wire        [31:0] w_sys_tmp103;
	wire signed [31:0] w_sys_tmp105;
	wire signed [31:0] w_sys_tmp106;
	wire        [31:0] w_sys_tmp107;
	wire signed [31:0] w_sys_tmp109;
	wire signed [31:0] w_sys_tmp110;
	wire        [31:0] w_sys_tmp112;
	wire signed [31:0] w_sys_tmp114;
	wire signed [31:0] w_sys_tmp115;
	wire signed [31:0] w_sys_tmp118;
	wire signed [31:0] w_sys_tmp119;
	wire signed [31:0] w_sys_tmp120;
	wire signed [31:0] w_sys_tmp121;
	wire               w_sys_tmp254;
	wire               w_sys_tmp255;
	wire signed [31:0] w_sys_tmp256;
	wire signed [31:0] w_sys_tmp259;
	wire signed [31:0] w_sys_tmp260;
	wire        [31:0] w_sys_tmp261;
	wire signed [31:0] w_sys_tmp265;
	wire signed [31:0] w_sys_tmp266;
	wire signed [31:0] w_sys_tmp271;
	wire signed [31:0] w_sys_tmp272;
	wire signed [31:0] w_sys_tmp277;
	wire signed [31:0] w_sys_tmp278;
	wire signed [31:0] w_sys_tmp283;
	wire signed [31:0] w_sys_tmp284;
	wire signed [31:0] w_sys_tmp289;
	wire signed [31:0] w_sys_tmp290;
	wire signed [31:0] w_sys_tmp295;
	wire signed [31:0] w_sys_tmp296;
	wire signed [31:0] w_sys_tmp301;
	wire signed [31:0] w_sys_tmp302;
	wire signed [31:0] w_sys_tmp307;
	wire signed [31:0] w_sys_tmp308;
	wire signed [31:0] w_sys_tmp313;
	wire signed [31:0] w_sys_tmp314;
	wire signed [31:0] w_sys_tmp319;
	wire signed [31:0] w_sys_tmp320;
	wire signed [31:0] w_sys_tmp325;
	wire signed [31:0] w_sys_tmp326;
	wire signed [31:0] w_sys_tmp343;
	wire signed [31:0] w_sys_tmp344;
	wire signed [31:0] w_sys_tmp349;
	wire signed [31:0] w_sys_tmp350;
	wire signed [31:0] w_sys_tmp355;
	wire signed [31:0] w_sys_tmp356;
	wire signed [31:0] w_sys_tmp361;
	wire signed [31:0] w_sys_tmp362;
	wire signed [31:0] w_sys_tmp367;
	wire signed [31:0] w_sys_tmp368;
	wire signed [31:0] w_sys_tmp373;
	wire signed [31:0] w_sys_tmp374;
	wire signed [31:0] w_sys_tmp379;
	wire signed [31:0] w_sys_tmp380;
	wire signed [31:0] w_sys_tmp385;
	wire signed [31:0] w_sys_tmp386;
	wire signed [31:0] w_sys_tmp391;
	wire signed [31:0] w_sys_tmp392;
	wire signed [31:0] w_sys_tmp397;
	wire signed [31:0] w_sys_tmp398;
	wire signed [31:0] w_sys_tmp415;
	wire signed [31:0] w_sys_tmp416;
	wire signed [31:0] w_sys_tmp421;
	wire signed [31:0] w_sys_tmp422;
	wire signed [31:0] w_sys_tmp427;
	wire signed [31:0] w_sys_tmp428;
	wire signed [31:0] w_sys_tmp433;
	wire signed [31:0] w_sys_tmp434;
	wire signed [31:0] w_sys_tmp439;
	wire signed [31:0] w_sys_tmp440;
	wire signed [31:0] w_sys_tmp445;
	wire signed [31:0] w_sys_tmp446;
	wire signed [31:0] w_sys_tmp451;
	wire signed [31:0] w_sys_tmp452;
	wire signed [31:0] w_sys_tmp457;
	wire signed [31:0] w_sys_tmp458;
	wire signed [31:0] w_sys_tmp463;
	wire signed [31:0] w_sys_tmp464;
	wire signed [31:0] w_sys_tmp469;
	wire signed [31:0] w_sys_tmp470;
	wire signed [31:0] w_sys_tmp475;
	wire signed [31:0] w_sys_tmp476;
	wire signed [31:0] w_sys_tmp481;
	wire signed [31:0] w_sys_tmp482;
	wire signed [31:0] w_sys_tmp487;
	wire signed [31:0] w_sys_tmp488;
	wire signed [31:0] w_sys_tmp493;
	wire signed [31:0] w_sys_tmp494;
	wire signed [31:0] w_sys_tmp499;
	wire signed [31:0] w_sys_tmp500;
	wire signed [31:0] w_sys_tmp505;
	wire signed [31:0] w_sys_tmp506;
	wire signed [31:0] w_sys_tmp511;
	wire signed [31:0] w_sys_tmp512;
	wire signed [31:0] w_sys_tmp517;
	wire signed [31:0] w_sys_tmp518;
	wire signed [31:0] w_sys_tmp523;
	wire signed [31:0] w_sys_tmp524;
	wire signed [31:0] w_sys_tmp529;
	wire signed [31:0] w_sys_tmp530;
	wire signed [31:0] w_sys_tmp535;
	wire signed [31:0] w_sys_tmp536;
	wire signed [31:0] w_sys_tmp553;
	wire signed [31:0] w_sys_tmp554;
	wire signed [31:0] w_sys_tmp559;
	wire signed [31:0] w_sys_tmp560;
	wire signed [31:0] w_sys_tmp565;
	wire signed [31:0] w_sys_tmp566;
	wire signed [31:0] w_sys_tmp571;
	wire signed [31:0] w_sys_tmp572;
	wire signed [31:0] w_sys_tmp577;
	wire signed [31:0] w_sys_tmp578;
	wire signed [31:0] w_sys_tmp583;
	wire signed [31:0] w_sys_tmp584;
	wire signed [31:0] w_sys_tmp589;
	wire signed [31:0] w_sys_tmp590;
	wire signed [31:0] w_sys_tmp595;
	wire signed [31:0] w_sys_tmp596;
	wire signed [31:0] w_sys_tmp601;
	wire signed [31:0] w_sys_tmp602;
	wire signed [31:0] w_sys_tmp607;
	wire signed [31:0] w_sys_tmp608;
	wire signed [31:0] w_sys_tmp625;
	wire signed [31:0] w_sys_tmp626;
	wire signed [31:0] w_sys_tmp631;
	wire signed [31:0] w_sys_tmp632;
	wire signed [31:0] w_sys_tmp637;
	wire signed [31:0] w_sys_tmp638;
	wire signed [31:0] w_sys_tmp643;
	wire signed [31:0] w_sys_tmp644;
	wire signed [31:0] w_sys_tmp649;
	wire signed [31:0] w_sys_tmp650;
	wire signed [31:0] w_sys_tmp655;
	wire signed [31:0] w_sys_tmp656;
	wire signed [31:0] w_sys_tmp661;
	wire signed [31:0] w_sys_tmp662;
	wire signed [31:0] w_sys_tmp667;
	wire signed [31:0] w_sys_tmp668;
	wire signed [31:0] w_sys_tmp673;
	wire signed [31:0] w_sys_tmp674;
	wire signed [31:0] w_sys_tmp678;
	wire signed [31:0] w_sys_tmp679;
	wire               w_sys_tmp680;
	wire               w_sys_tmp681;
	wire signed [31:0] w_sys_tmp682;
	wire signed [31:0] w_sys_tmp685;
	wire signed [31:0] w_sys_tmp686;
	wire        [31:0] w_sys_tmp687;
	wire signed [31:0] w_sys_tmp691;
	wire signed [31:0] w_sys_tmp692;
	wire signed [31:0] w_sys_tmp697;
	wire signed [31:0] w_sys_tmp698;
	wire signed [31:0] w_sys_tmp703;
	wire signed [31:0] w_sys_tmp704;
	wire signed [31:0] w_sys_tmp709;
	wire signed [31:0] w_sys_tmp710;
	wire signed [31:0] w_sys_tmp715;
	wire signed [31:0] w_sys_tmp716;
	wire signed [31:0] w_sys_tmp721;
	wire signed [31:0] w_sys_tmp722;
	wire signed [31:0] w_sys_tmp727;
	wire signed [31:0] w_sys_tmp728;
	wire signed [31:0] w_sys_tmp733;
	wire signed [31:0] w_sys_tmp734;
	wire signed [31:0] w_sys_tmp739;
	wire signed [31:0] w_sys_tmp740;
	wire signed [31:0] w_sys_tmp745;
	wire signed [31:0] w_sys_tmp746;
	wire signed [31:0] w_sys_tmp751;
	wire signed [31:0] w_sys_tmp752;
	wire signed [31:0] w_sys_tmp769;
	wire signed [31:0] w_sys_tmp770;
	wire signed [31:0] w_sys_tmp775;
	wire signed [31:0] w_sys_tmp776;
	wire signed [31:0] w_sys_tmp781;
	wire signed [31:0] w_sys_tmp782;
	wire signed [31:0] w_sys_tmp787;
	wire signed [31:0] w_sys_tmp788;
	wire signed [31:0] w_sys_tmp793;
	wire signed [31:0] w_sys_tmp794;
	wire signed [31:0] w_sys_tmp799;
	wire signed [31:0] w_sys_tmp800;
	wire signed [31:0] w_sys_tmp805;
	wire signed [31:0] w_sys_tmp806;
	wire signed [31:0] w_sys_tmp811;
	wire signed [31:0] w_sys_tmp812;
	wire signed [31:0] w_sys_tmp817;
	wire signed [31:0] w_sys_tmp818;
	wire signed [31:0] w_sys_tmp829;
	wire signed [31:0] w_sys_tmp830;
	wire signed [31:0] w_sys_tmp835;
	wire signed [31:0] w_sys_tmp836;
	wire signed [31:0] w_sys_tmp841;
	wire signed [31:0] w_sys_tmp842;
	wire signed [31:0] w_sys_tmp847;
	wire signed [31:0] w_sys_tmp848;
	wire signed [31:0] w_sys_tmp853;
	wire signed [31:0] w_sys_tmp854;
	wire signed [31:0] w_sys_tmp859;
	wire signed [31:0] w_sys_tmp860;
	wire signed [31:0] w_sys_tmp865;
	wire signed [31:0] w_sys_tmp866;
	wire signed [31:0] w_sys_tmp871;
	wire signed [31:0] w_sys_tmp872;
	wire signed [31:0] w_sys_tmp877;
	wire signed [31:0] w_sys_tmp878;
	wire signed [31:0] w_sys_tmp882;
	wire signed [31:0] w_sys_tmp883;
	wire               w_sys_tmp884;
	wire               w_sys_tmp885;
	wire signed [31:0] w_sys_tmp886;
	wire signed [31:0] w_sys_tmp889;
	wire signed [31:0] w_sys_tmp890;
	wire        [31:0] w_sys_tmp891;
	wire signed [31:0] w_sys_tmp895;
	wire signed [31:0] w_sys_tmp896;
	wire signed [31:0] w_sys_tmp901;
	wire signed [31:0] w_sys_tmp902;
	wire signed [31:0] w_sys_tmp907;
	wire signed [31:0] w_sys_tmp908;
	wire signed [31:0] w_sys_tmp913;
	wire signed [31:0] w_sys_tmp914;
	wire signed [31:0] w_sys_tmp919;
	wire signed [31:0] w_sys_tmp920;
	wire signed [31:0] w_sys_tmp925;
	wire signed [31:0] w_sys_tmp926;
	wire signed [31:0] w_sys_tmp931;
	wire signed [31:0] w_sys_tmp932;
	wire signed [31:0] w_sys_tmp937;
	wire signed [31:0] w_sys_tmp938;
	wire signed [31:0] w_sys_tmp943;
	wire signed [31:0] w_sys_tmp944;
	wire signed [31:0] w_sys_tmp949;
	wire signed [31:0] w_sys_tmp950;
	wire signed [31:0] w_sys_tmp954;
	wire signed [31:0] w_sys_tmp955;
	wire signed [31:0] w_sys_tmp959;
	wire signed [31:0] w_sys_tmp960;
	wire signed [31:0] w_sys_tmp964;
	wire signed [31:0] w_sys_tmp965;
	wire signed [31:0] w_sys_tmp969;
	wire signed [31:0] w_sys_tmp970;
	wire signed [31:0] w_sys_tmp974;
	wire signed [31:0] w_sys_tmp975;
	wire signed [31:0] w_sys_tmp979;
	wire signed [31:0] w_sys_tmp980;
	wire signed [31:0] w_sys_tmp984;
	wire signed [31:0] w_sys_tmp985;
	wire signed [31:0] w_sys_tmp989;
	wire signed [31:0] w_sys_tmp990;
	wire signed [31:0] w_sys_tmp994;
	wire signed [31:0] w_sys_tmp995;
	wire signed [31:0] w_sys_tmp999;
	wire signed [31:0] w_sys_tmp1000;
	wire signed [31:0] w_sys_tmp1004;
	wire signed [31:0] w_sys_tmp1005;
	wire signed [31:0] w_sys_tmp1009;
	wire signed [31:0] w_sys_tmp1010;
	wire signed [31:0] w_sys_tmp1014;
	wire signed [31:0] w_sys_tmp1015;
	wire signed [31:0] w_sys_tmp1019;
	wire signed [31:0] w_sys_tmp1020;
	wire signed [31:0] w_sys_tmp1024;
	wire signed [31:0] w_sys_tmp1025;
	wire signed [31:0] w_sys_tmp1029;
	wire signed [31:0] w_sys_tmp1030;
	wire signed [31:0] w_sys_tmp1034;
	wire signed [31:0] w_sys_tmp1035;
	wire signed [31:0] w_sys_tmp1039;
	wire signed [31:0] w_sys_tmp1040;
	wire signed [31:0] w_sys_tmp1044;
	wire signed [31:0] w_sys_tmp1045;
	wire signed [31:0] w_sys_tmp1049;
	wire signed [31:0] w_sys_tmp1050;
	wire signed [31:0] w_sys_tmp1054;
	wire signed [31:0] w_sys_tmp1055;
	wire signed [31:0] w_sys_tmp1059;
	wire signed [31:0] w_sys_tmp1060;
	wire signed [31:0] w_sys_tmp1064;
	wire signed [31:0] w_sys_tmp1065;
	wire signed [31:0] w_sys_tmp1069;
	wire signed [31:0] w_sys_tmp1070;
	wire signed [31:0] w_sys_tmp1074;
	wire signed [31:0] w_sys_tmp1075;
	wire signed [31:0] w_sys_tmp1079;
	wire signed [31:0] w_sys_tmp1080;
	wire signed [31:0] w_sys_tmp1084;
	wire signed [31:0] w_sys_tmp1085;
	wire signed [31:0] w_sys_tmp1089;
	wire signed [31:0] w_sys_tmp1090;
	wire signed [31:0] w_sys_tmp1094;
	wire signed [31:0] w_sys_tmp1095;
	wire signed [31:0] w_sys_tmp1099;
	wire signed [31:0] w_sys_tmp1100;
	wire signed [31:0] w_sys_tmp1104;
	wire signed [31:0] w_sys_tmp1105;
	wire signed [31:0] w_sys_tmp1109;
	wire signed [31:0] w_sys_tmp1110;
	wire signed [31:0] w_sys_tmp1114;
	wire signed [31:0] w_sys_tmp1115;
	wire signed [31:0] w_sys_tmp1119;
	wire signed [31:0] w_sys_tmp1120;
	wire signed [31:0] w_sys_tmp1124;
	wire signed [31:0] w_sys_tmp1125;
	wire signed [31:0] w_sys_tmp1129;
	wire signed [31:0] w_sys_tmp1130;
	wire signed [31:0] w_sys_tmp1134;
	wire signed [31:0] w_sys_tmp1135;
	wire signed [31:0] w_sys_tmp1139;
	wire signed [31:0] w_sys_tmp1140;
	wire signed [31:0] w_sys_tmp1144;
	wire signed [31:0] w_sys_tmp1145;
	wire signed [31:0] w_sys_tmp1149;
	wire signed [31:0] w_sys_tmp1150;
	wire signed [31:0] w_sys_tmp1154;
	wire signed [31:0] w_sys_tmp1155;
	wire signed [31:0] w_sys_tmp1159;
	wire signed [31:0] w_sys_tmp1160;
	wire signed [31:0] w_sys_tmp1164;
	wire signed [31:0] w_sys_tmp1165;
	wire signed [31:0] w_sys_tmp1169;
	wire signed [31:0] w_sys_tmp1170;
	wire signed [31:0] w_sys_tmp1174;
	wire signed [31:0] w_sys_tmp1175;
	wire signed [31:0] w_sys_tmp1179;
	wire signed [31:0] w_sys_tmp1180;
	wire signed [31:0] w_sys_tmp1184;
	wire signed [31:0] w_sys_tmp1185;
	wire signed [31:0] w_sys_tmp1188;
	wire signed [31:0] w_sys_tmp1189;
	wire               w_sys_tmp1190;
	wire               w_sys_tmp1191;
	wire signed [31:0] w_sys_tmp1192;
	wire signed [31:0] w_sys_tmp1195;
	wire signed [31:0] w_sys_tmp1196;
	wire        [31:0] w_sys_tmp1197;
	wire signed [31:0] w_sys_tmp1201;
	wire signed [31:0] w_sys_tmp1202;
	wire signed [31:0] w_sys_tmp1207;
	wire signed [31:0] w_sys_tmp1208;
	wire signed [31:0] w_sys_tmp1213;
	wire signed [31:0] w_sys_tmp1214;
	wire signed [31:0] w_sys_tmp1219;
	wire signed [31:0] w_sys_tmp1220;
	wire signed [31:0] w_sys_tmp1225;
	wire signed [31:0] w_sys_tmp1226;
	wire signed [31:0] w_sys_tmp1231;
	wire signed [31:0] w_sys_tmp1232;
	wire signed [31:0] w_sys_tmp1237;
	wire signed [31:0] w_sys_tmp1238;
	wire signed [31:0] w_sys_tmp1243;
	wire signed [31:0] w_sys_tmp1244;
	wire signed [31:0] w_sys_tmp1249;
	wire signed [31:0] w_sys_tmp1250;
	wire signed [31:0] w_sys_tmp1255;
	wire signed [31:0] w_sys_tmp1256;
	wire signed [31:0] w_sys_tmp1260;
	wire signed [31:0] w_sys_tmp1261;
	wire signed [31:0] w_sys_tmp1265;
	wire signed [31:0] w_sys_tmp1266;
	wire signed [31:0] w_sys_tmp1270;
	wire signed [31:0] w_sys_tmp1271;
	wire signed [31:0] w_sys_tmp1275;
	wire signed [31:0] w_sys_tmp1276;
	wire signed [31:0] w_sys_tmp1280;
	wire signed [31:0] w_sys_tmp1281;
	wire signed [31:0] w_sys_tmp1285;
	wire signed [31:0] w_sys_tmp1286;
	wire signed [31:0] w_sys_tmp1290;
	wire signed [31:0] w_sys_tmp1291;
	wire signed [31:0] w_sys_tmp1295;
	wire signed [31:0] w_sys_tmp1296;
	wire signed [31:0] w_sys_tmp1300;
	wire signed [31:0] w_sys_tmp1301;
	wire signed [31:0] w_sys_tmp1305;
	wire signed [31:0] w_sys_tmp1306;
	wire signed [31:0] w_sys_tmp1315;
	wire signed [31:0] w_sys_tmp1316;
	wire signed [31:0] w_sys_tmp1320;
	wire signed [31:0] w_sys_tmp1321;
	wire signed [31:0] w_sys_tmp1325;
	wire signed [31:0] w_sys_tmp1326;
	wire signed [31:0] w_sys_tmp1330;
	wire signed [31:0] w_sys_tmp1331;
	wire signed [31:0] w_sys_tmp1335;
	wire signed [31:0] w_sys_tmp1336;
	wire signed [31:0] w_sys_tmp1340;
	wire signed [31:0] w_sys_tmp1341;
	wire signed [31:0] w_sys_tmp1345;
	wire signed [31:0] w_sys_tmp1346;
	wire signed [31:0] w_sys_tmp1350;
	wire signed [31:0] w_sys_tmp1351;
	wire signed [31:0] w_sys_tmp1354;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 4'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 7'h1);
	assign w_fld_u_0_addr_0 = 9'sh0;
	assign w_fld_u_0_datain_0 = 32'h0;
	assign w_fld_u_0_r_w_0 = 1'h0;
	assign w_fld_u_0_ce_0 = w_sys_ce;
	assign w_fld_u_0_ce_1 = w_sys_ce;
	assign w_fld_uu_1_addr_0 = 9'sh0;
	assign w_fld_uu_1_datain_0 = 32'h0;
	assign w_fld_uu_1_r_w_0 = 1'h0;
	assign w_fld_uu_1_ce_0 = w_sys_ce;
	assign w_fld_uu_1_ce_1 = w_sys_ce;
	assign w_sub08_u_addr = ( (|r_sys_processing_methodID) ? r_sub08_u_addr : 10'sh0 ) ;
	assign w_sub08_u_datain = ( (|r_sys_processing_methodID) ? r_sub08_u_datain : 32'h0 ) ;
	assign w_sub08_u_r_w = ( (|r_sys_processing_methodID) ? r_sub08_u_r_w : 1'h0 ) ;
	assign w_sub08_result_addr = ( (|r_sys_processing_methodID) ? r_sub08_result_addr : 10'sh0 ) ;
	assign w_sub08_result_datain = ( (|r_sys_processing_methodID) ? r_sub08_result_datain : 32'h0 ) ;
	assign w_sub08_result_r_w = ( (|r_sys_processing_methodID) ? r_sub08_result_r_w : 1'h0 ) ;
	assign w_sub03_u_addr = ( (|r_sys_processing_methodID) ? r_sub03_u_addr : 10'sh0 ) ;
	assign w_sub03_u_datain = ( (|r_sys_processing_methodID) ? r_sub03_u_datain : 32'h0 ) ;
	assign w_sub03_u_r_w = ( (|r_sys_processing_methodID) ? r_sub03_u_r_w : 1'h0 ) ;
	assign w_sub03_result_addr = ( (|r_sys_processing_methodID) ? r_sub03_result_addr : 10'sh0 ) ;
	assign w_sub03_result_datain = ( (|r_sys_processing_methodID) ? r_sub03_result_datain : 32'h0 ) ;
	assign w_sub03_result_r_w = ( (|r_sys_processing_methodID) ? r_sub03_result_r_w : 1'h0 ) ;
	assign w_sub02_u_addr = ( (|r_sys_processing_methodID) ? r_sub02_u_addr : 10'sh0 ) ;
	assign w_sub02_u_datain = ( (|r_sys_processing_methodID) ? r_sub02_u_datain : 32'h0 ) ;
	assign w_sub02_u_r_w = ( (|r_sys_processing_methodID) ? r_sub02_u_r_w : 1'h0 ) ;
	assign w_sub02_result_addr = ( (|r_sys_processing_methodID) ? r_sub02_result_addr : 10'sh0 ) ;
	assign w_sub02_result_datain = ( (|r_sys_processing_methodID) ? r_sub02_result_datain : 32'h0 ) ;
	assign w_sub02_result_r_w = ( (|r_sys_processing_methodID) ? r_sub02_result_r_w : 1'h0 ) ;
	assign w_sub01_u_addr = ( (|r_sys_processing_methodID) ? r_sub01_u_addr : 10'sh0 ) ;
	assign w_sub01_u_datain = ( (|r_sys_processing_methodID) ? r_sub01_u_datain : 32'h0 ) ;
	assign w_sub01_u_r_w = ( (|r_sys_processing_methodID) ? r_sub01_u_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 10'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub00_u_addr = ( (|r_sys_processing_methodID) ? r_sub00_u_addr : 10'sh0 ) ;
	assign w_sub00_u_datain = ( (|r_sys_processing_methodID) ? r_sub00_u_datain : 32'h0 ) ;
	assign w_sub00_u_r_w = ( (|r_sys_processing_methodID) ? r_sub00_u_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 10'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sub07_u_addr = ( (|r_sys_processing_methodID) ? r_sub07_u_addr : 10'sh0 ) ;
	assign w_sub07_u_datain = ( (|r_sys_processing_methodID) ? r_sub07_u_datain : 32'h0 ) ;
	assign w_sub07_u_r_w = ( (|r_sys_processing_methodID) ? r_sub07_u_r_w : 1'h0 ) ;
	assign w_sub07_result_addr = ( (|r_sys_processing_methodID) ? r_sub07_result_addr : 10'sh0 ) ;
	assign w_sub07_result_datain = ( (|r_sys_processing_methodID) ? r_sub07_result_datain : 32'h0 ) ;
	assign w_sub07_result_r_w = ( (|r_sys_processing_methodID) ? r_sub07_result_r_w : 1'h0 ) ;
	assign w_sub06_u_addr = ( (|r_sys_processing_methodID) ? r_sub06_u_addr : 10'sh0 ) ;
	assign w_sub06_u_datain = ( (|r_sys_processing_methodID) ? r_sub06_u_datain : 32'h0 ) ;
	assign w_sub06_u_r_w = ( (|r_sys_processing_methodID) ? r_sub06_u_r_w : 1'h0 ) ;
	assign w_sub06_result_addr = ( (|r_sys_processing_methodID) ? r_sub06_result_addr : 10'sh0 ) ;
	assign w_sub06_result_datain = ( (|r_sys_processing_methodID) ? r_sub06_result_datain : 32'h0 ) ;
	assign w_sub06_result_r_w = ( (|r_sys_processing_methodID) ? r_sub06_result_r_w : 1'h0 ) ;
	assign w_sub05_u_addr = ( (|r_sys_processing_methodID) ? r_sub05_u_addr : 10'sh0 ) ;
	assign w_sub05_u_datain = ( (|r_sys_processing_methodID) ? r_sub05_u_datain : 32'h0 ) ;
	assign w_sub05_u_r_w = ( (|r_sys_processing_methodID) ? r_sub05_u_r_w : 1'h0 ) ;
	assign w_sub05_result_addr = ( (|r_sys_processing_methodID) ? r_sub05_result_addr : 10'sh0 ) ;
	assign w_sub05_result_datain = ( (|r_sys_processing_methodID) ? r_sub05_result_datain : 32'h0 ) ;
	assign w_sub05_result_r_w = ( (|r_sys_processing_methodID) ? r_sub05_result_r_w : 1'h0 ) ;
	assign w_sub04_u_addr = ( (|r_sys_processing_methodID) ? r_sub04_u_addr : 10'sh0 ) ;
	assign w_sub04_u_datain = ( (|r_sys_processing_methodID) ? r_sub04_u_datain : 32'h0 ) ;
	assign w_sub04_u_r_w = ( (|r_sys_processing_methodID) ? r_sub04_u_r_w : 1'h0 ) ;
	assign w_sub04_result_addr = ( (|r_sys_processing_methodID) ? r_sub04_result_addr : 10'sh0 ) ;
	assign w_sub04_result_datain = ( (|r_sys_processing_methodID) ? r_sub04_result_datain : 32'h0 ) ;
	assign w_sub04_result_r_w = ( (|r_sys_processing_methodID) ? r_sub04_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh0000001f;
	assign w_sys_tmp3 = 32'sh00000002;
	assign w_sys_tmp4 = ( !w_sys_tmp5 );
	assign w_sys_tmp5 = (r_run_my_15 < r_run_k_11);
	assign w_sys_tmp6 = (r_run_k_11 + w_sys_intOne);
	assign w_sys_tmp7 = ( !w_sys_tmp8 );
	assign w_sys_tmp8 = (r_run_mx_14 < r_run_j_12);
	assign w_sys_tmp11 = (w_sys_tmp12 + r_run_k_11);
	assign w_sys_tmp12 = (r_run_j_12 * w_sys_tmp13);
	assign w_sys_tmp13 = 32'sh0000001f;
	assign w_sys_tmp14 = 32'h0;
	assign w_sys_tmp16 = (w_sys_tmp17 + r_run_k_11);
	assign w_sys_tmp17 = (r_run_copy0_j_17 * w_sys_tmp13);
	assign w_sys_tmp20 = (r_run_copy0_j_17 + w_sys_intOne);
	assign w_sys_tmp21 = (r_run_j_12 + w_sys_intOne);
	assign w_sys_tmp94 = ( !w_sys_tmp95 );
	assign w_sys_tmp95 = (r_run_nlast_16 < r_run_n_13);
	assign w_sys_tmp96 = (r_run_n_13 + w_sys_intOne);
	assign w_sys_tmp97 = ( !w_sys_tmp98 );
	assign w_sys_tmp98 = (r_run_my_15 < r_run_j_12);
	assign w_sys_tmp101 = (w_sys_tmp102 + r_run_j_12);
	assign w_sys_tmp102 = 32'sh0000001f;
	assign w_sys_tmp103 = 32'h3f000000;
	assign w_sys_tmp105 = (w_sys_tmp106 + r_run_copy2_j_20);
	assign w_sys_tmp106 = 32'sh000001b9;
	assign w_sys_tmp107 = 32'h0;
	assign w_sys_tmp109 = (w_sys_tmp110 + w_sys_intOne);
	assign w_sys_tmp110 = (r_run_copy1_j_19 * w_sys_tmp102);
	assign w_sys_tmp112 = 32'h3f800000;
	assign w_sys_tmp114 = (w_sys_tmp115 + r_run_my_15);
	assign w_sys_tmp115 = (r_run_copy0_j_18 * w_sys_tmp102);
	assign w_sys_tmp118 = (r_run_copy0_j_18 + w_sys_intOne);
	assign w_sys_tmp119 = (r_run_copy1_j_19 + w_sys_intOne);
	assign w_sys_tmp120 = (r_run_copy2_j_20 + w_sys_intOne);
	assign w_sys_tmp121 = (r_run_j_12 + w_sys_intOne);
	assign w_sys_tmp254 = ( !w_sys_tmp255 );
	assign w_sys_tmp255 = (w_sys_tmp256 < r_run_k_11);
	assign w_sys_tmp256 = 32'sh0000000c;
	assign w_sys_tmp259 = (w_sys_tmp260 + r_run_k_11);
	assign w_sys_tmp260 = 32'sh0000001f;
	assign w_sys_tmp261 = w_fld_u_0_dataout_1;
	assign w_sys_tmp265 = (w_sys_tmp266 + r_run_k_11);
	assign w_sys_tmp266 = 32'sh0000003e;
	assign w_sys_tmp271 = (w_sys_tmp272 + r_run_k_11);
	assign w_sys_tmp272 = 32'sh0000005d;
	assign w_sys_tmp277 = (w_sys_tmp278 + r_run_k_11);
	assign w_sys_tmp278 = 32'sh0000007c;
	assign w_sys_tmp283 = (w_sys_tmp284 + r_run_k_11);
	assign w_sys_tmp284 = 32'sh0000009b;
	assign w_sys_tmp289 = (w_sys_tmp290 + r_run_k_11);
	assign w_sys_tmp290 = 32'sh000000ba;
	assign w_sys_tmp295 = (w_sys_tmp296 + r_run_k_11);
	assign w_sys_tmp296 = 32'sh000000d9;
	assign w_sys_tmp301 = (w_sys_tmp302 + r_run_k_11);
	assign w_sys_tmp302 = 32'sh000000f8;
	assign w_sys_tmp307 = (w_sys_tmp308 + r_run_k_11);
	assign w_sys_tmp308 = 32'sh00000117;
	assign w_sys_tmp313 = (w_sys_tmp314 + r_run_k_11);
	assign w_sys_tmp314 = 32'sh00000136;
	assign w_sys_tmp319 = (w_sys_tmp320 + r_run_k_11);
	assign w_sys_tmp320 = 32'sh00000155;
	assign w_sys_tmp325 = (w_sys_tmp326 + r_run_k_11);
	assign w_sys_tmp326 = 32'sh00000174;
	assign w_sys_tmp343 = (w_sys_tmp344 + r_run_k_11);
	assign w_sys_tmp344 = 32'sh00000193;
	assign w_sys_tmp349 = (w_sys_tmp350 + r_run_k_11);
	assign w_sys_tmp350 = 32'sh000001b2;
	assign w_sys_tmp355 = (w_sys_tmp356 + r_run_k_11);
	assign w_sys_tmp356 = 32'sh000001d1;
	assign w_sys_tmp361 = (w_sys_tmp362 + r_run_k_11);
	assign w_sys_tmp362 = 32'sh000001f0;
	assign w_sys_tmp367 = (w_sys_tmp368 + r_run_k_11);
	assign w_sys_tmp368 = 32'sh0000020f;
	assign w_sys_tmp373 = (w_sys_tmp374 + r_run_k_11);
	assign w_sys_tmp374 = 32'sh0000022e;
	assign w_sys_tmp379 = (w_sys_tmp380 + r_run_k_11);
	assign w_sys_tmp380 = 32'sh0000024d;
	assign w_sys_tmp385 = (w_sys_tmp386 + r_run_k_11);
	assign w_sys_tmp386 = 32'sh0000026c;
	assign w_sys_tmp391 = (w_sys_tmp392 + r_run_k_11);
	assign w_sys_tmp392 = 32'sh0000028b;
	assign w_sys_tmp397 = (w_sys_tmp398 + r_run_k_11);
	assign w_sys_tmp398 = 32'sh000002aa;
	assign w_sys_tmp415 = (w_sys_tmp416 + r_run_k_11);
	assign w_sys_tmp416 = 32'sh000002c9;
	assign w_sys_tmp421 = (w_sys_tmp422 + r_run_k_11);
	assign w_sys_tmp422 = 32'sh000002e8;
	assign w_sys_tmp427 = (w_sys_tmp428 + r_run_k_11);
	assign w_sys_tmp428 = 32'sh00000307;
	assign w_sys_tmp433 = (w_sys_tmp434 + r_run_k_11);
	assign w_sys_tmp434 = 32'sh00000326;
	assign w_sys_tmp439 = (w_sys_tmp440 + r_run_k_11);
	assign w_sys_tmp440 = 32'sh00000345;
	assign w_sys_tmp445 = (w_sys_tmp446 + r_run_k_11);
	assign w_sys_tmp446 = 32'sh00000364;
	assign w_sys_tmp451 = (w_sys_tmp452 + r_run_k_11);
	assign w_sys_tmp452 = 32'sh00000383;
	assign w_sys_tmp457 = (w_sys_tmp458 + r_run_k_11);
	assign w_sys_tmp458 = 32'sh000003a2;
	assign w_sys_tmp463 = (w_sys_tmp464 + r_run_k_11);
	assign w_sys_tmp464 = 32'sh000003c1;
	assign w_sys_tmp469 = (w_sys_tmp470 + r_run_k_11);
	assign w_sys_tmp470 = 32'sh00000029;
	assign w_sys_tmp475 = (w_sys_tmp476 + r_run_k_11);
	assign w_sys_tmp476 = 32'sh00000048;
	assign w_sys_tmp481 = (w_sys_tmp482 + r_run_k_11);
	assign w_sys_tmp482 = 32'sh00000067;
	assign w_sys_tmp487 = (w_sys_tmp488 + r_run_k_11);
	assign w_sys_tmp488 = 32'sh00000086;
	assign w_sys_tmp493 = (w_sys_tmp494 + r_run_k_11);
	assign w_sys_tmp494 = 32'sh000000a5;
	assign w_sys_tmp499 = (w_sys_tmp500 + r_run_k_11);
	assign w_sys_tmp500 = 32'sh000000c4;
	assign w_sys_tmp505 = (w_sys_tmp506 + r_run_k_11);
	assign w_sys_tmp506 = 32'sh000000e3;
	assign w_sys_tmp511 = (w_sys_tmp512 + r_run_k_11);
	assign w_sys_tmp512 = 32'sh00000102;
	assign w_sys_tmp517 = (w_sys_tmp518 + r_run_k_11);
	assign w_sys_tmp518 = 32'sh00000121;
	assign w_sys_tmp523 = (w_sys_tmp524 + r_run_k_11);
	assign w_sys_tmp524 = 32'sh00000140;
	assign w_sys_tmp529 = (w_sys_tmp530 + r_run_k_11);
	assign w_sys_tmp530 = 32'sh0000015f;
	assign w_sys_tmp535 = (w_sys_tmp536 + r_run_k_11);
	assign w_sys_tmp536 = 32'sh0000017e;
	assign w_sys_tmp553 = (w_sys_tmp554 + r_run_k_11);
	assign w_sys_tmp554 = 32'sh0000019d;
	assign w_sys_tmp559 = (w_sys_tmp560 + r_run_k_11);
	assign w_sys_tmp560 = 32'sh000001bc;
	assign w_sys_tmp565 = (w_sys_tmp566 + r_run_k_11);
	assign w_sys_tmp566 = 32'sh000001db;
	assign w_sys_tmp571 = (w_sys_tmp572 + r_run_k_11);
	assign w_sys_tmp572 = 32'sh000001fa;
	assign w_sys_tmp577 = (w_sys_tmp578 + r_run_k_11);
	assign w_sys_tmp578 = 32'sh00000219;
	assign w_sys_tmp583 = (w_sys_tmp584 + r_run_k_11);
	assign w_sys_tmp584 = 32'sh00000238;
	assign w_sys_tmp589 = (w_sys_tmp590 + r_run_k_11);
	assign w_sys_tmp590 = 32'sh00000257;
	assign w_sys_tmp595 = (w_sys_tmp596 + r_run_k_11);
	assign w_sys_tmp596 = 32'sh00000276;
	assign w_sys_tmp601 = (w_sys_tmp602 + r_run_k_11);
	assign w_sys_tmp602 = 32'sh00000295;
	assign w_sys_tmp607 = (w_sys_tmp608 + r_run_k_11);
	assign w_sys_tmp608 = 32'sh000002b4;
	assign w_sys_tmp625 = (w_sys_tmp626 + r_run_k_11);
	assign w_sys_tmp626 = 32'sh000002d3;
	assign w_sys_tmp631 = (w_sys_tmp632 + r_run_k_11);
	assign w_sys_tmp632 = 32'sh000002f2;
	assign w_sys_tmp637 = (w_sys_tmp638 + r_run_k_11);
	assign w_sys_tmp638 = 32'sh00000311;
	assign w_sys_tmp643 = (w_sys_tmp644 + r_run_k_11);
	assign w_sys_tmp644 = 32'sh00000330;
	assign w_sys_tmp649 = (w_sys_tmp650 + r_run_k_11);
	assign w_sys_tmp650 = 32'sh0000034f;
	assign w_sys_tmp655 = (w_sys_tmp656 + r_run_k_11);
	assign w_sys_tmp656 = 32'sh0000036e;
	assign w_sys_tmp661 = (w_sys_tmp662 + r_run_k_11);
	assign w_sys_tmp662 = 32'sh0000038d;
	assign w_sys_tmp667 = (w_sys_tmp668 + r_run_k_11);
	assign w_sys_tmp668 = 32'sh000003ac;
	assign w_sys_tmp673 = (w_sys_tmp674 + r_run_k_11);
	assign w_sys_tmp674 = 32'sh000003cb;
	assign w_sys_tmp678 = (r_run_k_11 + w_sys_intOne);
	assign w_sys_tmp679 = 32'sh00000015;
	assign w_sys_tmp680 = ( !w_sys_tmp681 );
	assign w_sys_tmp681 = (w_sys_tmp682 < r_run_k_11);
	assign w_sys_tmp682 = 32'sh0000001f;
	assign w_sys_tmp685 = (w_sys_tmp686 + r_run_k_11);
	assign w_sys_tmp686 = 32'sh0000001f;
	assign w_sys_tmp687 = w_fld_u_0_dataout_1;
	assign w_sys_tmp691 = (w_sys_tmp692 + r_run_k_11);
	assign w_sys_tmp692 = 32'sh0000003e;
	assign w_sys_tmp697 = (w_sys_tmp698 + r_run_k_11);
	assign w_sys_tmp698 = 32'sh0000005d;
	assign w_sys_tmp703 = (w_sys_tmp704 + r_run_k_11);
	assign w_sys_tmp704 = 32'sh0000007c;
	assign w_sys_tmp709 = (w_sys_tmp710 + r_run_k_11);
	assign w_sys_tmp710 = 32'sh0000009b;
	assign w_sys_tmp715 = (w_sys_tmp716 + r_run_k_11);
	assign w_sys_tmp716 = 32'sh000000ba;
	assign w_sys_tmp721 = (w_sys_tmp722 + r_run_k_11);
	assign w_sys_tmp722 = 32'sh000000d9;
	assign w_sys_tmp727 = (w_sys_tmp728 + r_run_k_11);
	assign w_sys_tmp728 = 32'sh000000f8;
	assign w_sys_tmp733 = (w_sys_tmp734 + r_run_k_11);
	assign w_sys_tmp734 = 32'sh00000117;
	assign w_sys_tmp739 = (w_sys_tmp740 + r_run_k_11);
	assign w_sys_tmp740 = 32'sh00000136;
	assign w_sys_tmp745 = (w_sys_tmp746 + r_run_k_11);
	assign w_sys_tmp746 = 32'sh00000155;
	assign w_sys_tmp751 = (w_sys_tmp752 + r_run_k_11);
	assign w_sys_tmp752 = 32'sh00000174;
	assign w_sys_tmp769 = (w_sys_tmp770 + r_run_k_11);
	assign w_sys_tmp770 = 32'sh00000193;
	assign w_sys_tmp775 = (w_sys_tmp776 + r_run_k_11);
	assign w_sys_tmp776 = 32'sh000001b2;
	assign w_sys_tmp781 = (w_sys_tmp782 + r_run_k_11);
	assign w_sys_tmp782 = 32'sh000001d1;
	assign w_sys_tmp787 = (w_sys_tmp788 + r_run_k_11);
	assign w_sys_tmp788 = 32'sh000001f0;
	assign w_sys_tmp793 = (w_sys_tmp794 + r_run_k_11);
	assign w_sys_tmp794 = 32'sh0000020f;
	assign w_sys_tmp799 = (w_sys_tmp800 + r_run_k_11);
	assign w_sys_tmp800 = 32'sh0000022e;
	assign w_sys_tmp805 = (w_sys_tmp806 + r_run_k_11);
	assign w_sys_tmp806 = 32'sh0000024d;
	assign w_sys_tmp811 = (w_sys_tmp812 + r_run_k_11);
	assign w_sys_tmp812 = 32'sh0000026c;
	assign w_sys_tmp817 = (w_sys_tmp818 + r_run_k_11);
	assign w_sys_tmp818 = 32'sh0000028b;
	assign w_sys_tmp829 = (w_sys_tmp830 + r_run_k_11);
	assign w_sys_tmp830 = 32'sh000002aa;
	assign w_sys_tmp835 = (w_sys_tmp836 + r_run_k_11);
	assign w_sys_tmp836 = 32'sh000002c9;
	assign w_sys_tmp841 = (w_sys_tmp842 + r_run_k_11);
	assign w_sys_tmp842 = 32'sh000002e8;
	assign w_sys_tmp847 = (w_sys_tmp848 + r_run_k_11);
	assign w_sys_tmp848 = 32'sh00000307;
	assign w_sys_tmp853 = (w_sys_tmp854 + r_run_k_11);
	assign w_sys_tmp854 = 32'sh00000326;
	assign w_sys_tmp859 = (w_sys_tmp860 + r_run_k_11);
	assign w_sys_tmp860 = 32'sh00000345;
	assign w_sys_tmp865 = (w_sys_tmp866 + r_run_k_11);
	assign w_sys_tmp866 = 32'sh00000364;
	assign w_sys_tmp871 = (w_sys_tmp872 + r_run_k_11);
	assign w_sys_tmp872 = 32'sh00000383;
	assign w_sys_tmp877 = (w_sys_tmp878 + r_run_k_11);
	assign w_sys_tmp878 = 32'sh000003a2;
	assign w_sys_tmp882 = (r_run_k_11 + w_sys_intOne);
	assign w_sys_tmp883 = 32'sh00000002;
	assign w_sys_tmp884 = ( !w_sys_tmp885 );
	assign w_sys_tmp885 = (w_sys_tmp886 < r_run_k_11);
	assign w_sys_tmp886 = 32'sh0000000b;
	assign w_sys_tmp889 = (w_sys_tmp890 + r_run_k_11);
	assign w_sys_tmp890 = 32'sh0000003e;
	assign w_sys_tmp891 = w_sub00_result_dataout;
	assign w_sys_tmp895 = (w_sys_tmp896 + r_run_k_11);
	assign w_sys_tmp896 = 32'sh0000005d;
	assign w_sys_tmp901 = (w_sys_tmp902 + r_run_k_11);
	assign w_sys_tmp902 = 32'sh0000007c;
	assign w_sys_tmp907 = (w_sys_tmp908 + r_run_k_11);
	assign w_sys_tmp908 = 32'sh0000009b;
	assign w_sys_tmp913 = (w_sys_tmp914 + r_run_k_11);
	assign w_sys_tmp914 = 32'sh000000ba;
	assign w_sys_tmp919 = (w_sys_tmp920 + r_run_k_11);
	assign w_sys_tmp920 = 32'sh000000d9;
	assign w_sys_tmp925 = (w_sys_tmp926 + r_run_k_11);
	assign w_sys_tmp926 = 32'sh000000f8;
	assign w_sys_tmp931 = (w_sys_tmp932 + r_run_k_11);
	assign w_sys_tmp932 = 32'sh00000117;
	assign w_sys_tmp937 = (w_sys_tmp938 + r_run_k_11);
	assign w_sys_tmp938 = 32'sh00000136;
	assign w_sys_tmp943 = (w_sys_tmp944 + r_run_k_11);
	assign w_sys_tmp944 = 32'sh00000155;
	assign w_sys_tmp949 = (w_sys_tmp950 + r_run_k_11);
	assign w_sys_tmp950 = 32'sh00000174;
	assign w_sys_tmp954 = (w_sys_tmp955 + r_run_k_11);
	assign w_sys_tmp955 = 32'sh00000193;
	assign w_sys_tmp959 = (w_sys_tmp960 + r_run_k_11);
	assign w_sys_tmp960 = 32'sh000001b2;
	assign w_sys_tmp964 = (w_sys_tmp965 + r_run_k_11);
	assign w_sys_tmp965 = 32'sh000001d1;
	assign w_sys_tmp969 = (w_sys_tmp970 + r_run_k_11);
	assign w_sys_tmp970 = 32'sh000001f0;
	assign w_sys_tmp974 = (w_sys_tmp975 + r_run_k_11);
	assign w_sys_tmp975 = 32'sh0000020f;
	assign w_sys_tmp979 = (w_sys_tmp980 + r_run_k_11);
	assign w_sys_tmp980 = 32'sh0000022e;
	assign w_sys_tmp984 = (w_sys_tmp985 + r_run_k_11);
	assign w_sys_tmp985 = 32'sh0000024d;
	assign w_sys_tmp989 = (w_sys_tmp990 + r_run_k_11);
	assign w_sys_tmp990 = 32'sh0000026c;
	assign w_sys_tmp994 = (w_sys_tmp995 + r_run_k_11);
	assign w_sys_tmp995 = 32'sh0000028b;
	assign w_sys_tmp999 = (w_sys_tmp1000 + r_run_k_11);
	assign w_sys_tmp1000 = 32'sh000002aa;
	assign w_sys_tmp1004 = (w_sys_tmp1005 + r_run_k_11);
	assign w_sys_tmp1005 = 32'sh000002c9;
	assign w_sys_tmp1009 = (w_sys_tmp1010 + r_run_k_11);
	assign w_sys_tmp1010 = 32'sh000002e8;
	assign w_sys_tmp1014 = (w_sys_tmp1015 + r_run_k_11);
	assign w_sys_tmp1015 = 32'sh00000307;
	assign w_sys_tmp1019 = (w_sys_tmp1020 + r_run_k_11);
	assign w_sys_tmp1020 = 32'sh00000326;
	assign w_sys_tmp1024 = (w_sys_tmp1025 + r_run_k_11);
	assign w_sys_tmp1025 = 32'sh00000345;
	assign w_sys_tmp1029 = (w_sys_tmp1030 + r_run_k_11);
	assign w_sys_tmp1030 = 32'sh00000364;
	assign w_sys_tmp1034 = (w_sys_tmp1035 + r_run_k_11);
	assign w_sys_tmp1035 = 32'sh00000383;
	assign w_sys_tmp1039 = (w_sys_tmp1040 + r_run_k_11);
	assign w_sys_tmp1040 = 32'sh000003a2;
	assign w_sys_tmp1044 = (w_sys_tmp1045 + r_run_k_11);
	assign w_sys_tmp1045 = 32'sh00000048;
	assign w_sys_tmp1049 = (w_sys_tmp1050 + r_run_k_11);
	assign w_sys_tmp1050 = 32'sh00000067;
	assign w_sys_tmp1054 = (w_sys_tmp1055 + r_run_k_11);
	assign w_sys_tmp1055 = 32'sh00000086;
	assign w_sys_tmp1059 = (w_sys_tmp1060 + r_run_k_11);
	assign w_sys_tmp1060 = 32'sh000000a5;
	assign w_sys_tmp1064 = (w_sys_tmp1065 + r_run_k_11);
	assign w_sys_tmp1065 = 32'sh000000c4;
	assign w_sys_tmp1069 = (w_sys_tmp1070 + r_run_k_11);
	assign w_sys_tmp1070 = 32'sh000000e3;
	assign w_sys_tmp1074 = (w_sys_tmp1075 + r_run_k_11);
	assign w_sys_tmp1075 = 32'sh00000102;
	assign w_sys_tmp1079 = (w_sys_tmp1080 + r_run_k_11);
	assign w_sys_tmp1080 = 32'sh00000121;
	assign w_sys_tmp1084 = (w_sys_tmp1085 + r_run_k_11);
	assign w_sys_tmp1085 = 32'sh00000140;
	assign w_sys_tmp1089 = (w_sys_tmp1090 + r_run_k_11);
	assign w_sys_tmp1090 = 32'sh0000015f;
	assign w_sys_tmp1094 = (w_sys_tmp1095 + r_run_k_11);
	assign w_sys_tmp1095 = 32'sh0000017e;
	assign w_sys_tmp1099 = (w_sys_tmp1100 + r_run_k_11);
	assign w_sys_tmp1100 = 32'sh0000019d;
	assign w_sys_tmp1104 = (w_sys_tmp1105 + r_run_k_11);
	assign w_sys_tmp1105 = 32'sh000001bc;
	assign w_sys_tmp1109 = (w_sys_tmp1110 + r_run_k_11);
	assign w_sys_tmp1110 = 32'sh000001db;
	assign w_sys_tmp1114 = (w_sys_tmp1115 + r_run_k_11);
	assign w_sys_tmp1115 = 32'sh000001fa;
	assign w_sys_tmp1119 = (w_sys_tmp1120 + r_run_k_11);
	assign w_sys_tmp1120 = 32'sh00000219;
	assign w_sys_tmp1124 = (w_sys_tmp1125 + r_run_k_11);
	assign w_sys_tmp1125 = 32'sh00000238;
	assign w_sys_tmp1129 = (w_sys_tmp1130 + r_run_k_11);
	assign w_sys_tmp1130 = 32'sh00000257;
	assign w_sys_tmp1134 = (w_sys_tmp1135 + r_run_k_11);
	assign w_sys_tmp1135 = 32'sh00000276;
	assign w_sys_tmp1139 = (w_sys_tmp1140 + r_run_k_11);
	assign w_sys_tmp1140 = 32'sh00000295;
	assign w_sys_tmp1144 = (w_sys_tmp1145 + r_run_k_11);
	assign w_sys_tmp1145 = 32'sh000002b4;
	assign w_sys_tmp1149 = (w_sys_tmp1150 + r_run_k_11);
	assign w_sys_tmp1150 = 32'sh000002d3;
	assign w_sys_tmp1154 = (w_sys_tmp1155 + r_run_k_11);
	assign w_sys_tmp1155 = 32'sh000002f2;
	assign w_sys_tmp1159 = (w_sys_tmp1160 + r_run_k_11);
	assign w_sys_tmp1160 = 32'sh00000311;
	assign w_sys_tmp1164 = (w_sys_tmp1165 + r_run_k_11);
	assign w_sys_tmp1165 = 32'sh00000330;
	assign w_sys_tmp1169 = (w_sys_tmp1170 + r_run_k_11);
	assign w_sys_tmp1170 = 32'sh0000034f;
	assign w_sys_tmp1174 = (w_sys_tmp1175 + r_run_k_11);
	assign w_sys_tmp1175 = 32'sh0000036e;
	assign w_sys_tmp1179 = (w_sys_tmp1180 + r_run_k_11);
	assign w_sys_tmp1180 = 32'sh0000038d;
	assign w_sys_tmp1184 = (w_sys_tmp1185 + r_run_k_11);
	assign w_sys_tmp1185 = 32'sh000003ac;
	assign w_sys_tmp1188 = (r_run_k_11 + w_sys_intOne);
	assign w_sys_tmp1189 = 32'sh00000016;
	assign w_sys_tmp1190 = ( !w_sys_tmp1191 );
	assign w_sys_tmp1191 = (w_sys_tmp1192 < r_run_k_11);
	assign w_sys_tmp1192 = 32'sh0000001e;
	assign w_sys_tmp1195 = (w_sys_tmp1196 + r_run_k_11);
	assign w_sys_tmp1196 = 32'sh0000003e;
	assign w_sys_tmp1197 = w_sub06_result_dataout;
	assign w_sys_tmp1201 = (w_sys_tmp1202 + r_run_k_11);
	assign w_sys_tmp1202 = 32'sh0000005d;
	assign w_sys_tmp1207 = (w_sys_tmp1208 + r_run_k_11);
	assign w_sys_tmp1208 = 32'sh0000007c;
	assign w_sys_tmp1213 = (w_sys_tmp1214 + r_run_k_11);
	assign w_sys_tmp1214 = 32'sh0000009b;
	assign w_sys_tmp1219 = (w_sys_tmp1220 + r_run_k_11);
	assign w_sys_tmp1220 = 32'sh000000ba;
	assign w_sys_tmp1225 = (w_sys_tmp1226 + r_run_k_11);
	assign w_sys_tmp1226 = 32'sh000000d9;
	assign w_sys_tmp1231 = (w_sys_tmp1232 + r_run_k_11);
	assign w_sys_tmp1232 = 32'sh000000f8;
	assign w_sys_tmp1237 = (w_sys_tmp1238 + r_run_k_11);
	assign w_sys_tmp1238 = 32'sh00000117;
	assign w_sys_tmp1243 = (w_sys_tmp1244 + r_run_k_11);
	assign w_sys_tmp1244 = 32'sh00000136;
	assign w_sys_tmp1249 = (w_sys_tmp1250 + r_run_k_11);
	assign w_sys_tmp1250 = 32'sh00000155;
	assign w_sys_tmp1255 = (w_sys_tmp1256 + r_run_k_11);
	assign w_sys_tmp1256 = 32'sh00000174;
	assign w_sys_tmp1260 = (w_sys_tmp1261 + r_run_k_11);
	assign w_sys_tmp1261 = 32'sh00000193;
	assign w_sys_tmp1265 = (w_sys_tmp1266 + r_run_k_11);
	assign w_sys_tmp1266 = 32'sh000001b2;
	assign w_sys_tmp1270 = (w_sys_tmp1271 + r_run_k_11);
	assign w_sys_tmp1271 = 32'sh000001d1;
	assign w_sys_tmp1275 = (w_sys_tmp1276 + r_run_k_11);
	assign w_sys_tmp1276 = 32'sh000001f0;
	assign w_sys_tmp1280 = (w_sys_tmp1281 + r_run_k_11);
	assign w_sys_tmp1281 = 32'sh0000020f;
	assign w_sys_tmp1285 = (w_sys_tmp1286 + r_run_k_11);
	assign w_sys_tmp1286 = 32'sh0000022e;
	assign w_sys_tmp1290 = (w_sys_tmp1291 + r_run_k_11);
	assign w_sys_tmp1291 = 32'sh0000024d;
	assign w_sys_tmp1295 = (w_sys_tmp1296 + r_run_k_11);
	assign w_sys_tmp1296 = 32'sh0000026c;
	assign w_sys_tmp1300 = (w_sys_tmp1301 + r_run_k_11);
	assign w_sys_tmp1301 = 32'sh0000028b;
	assign w_sys_tmp1305 = (w_sys_tmp1306 + r_run_k_11);
	assign w_sys_tmp1306 = 32'sh000002aa;
	assign w_sys_tmp1315 = (w_sys_tmp1316 + r_run_k_11);
	assign w_sys_tmp1316 = 32'sh000002c9;
	assign w_sys_tmp1320 = (w_sys_tmp1321 + r_run_k_11);
	assign w_sys_tmp1321 = 32'sh000002e8;
	assign w_sys_tmp1325 = (w_sys_tmp1326 + r_run_k_11);
	assign w_sys_tmp1326 = 32'sh00000307;
	assign w_sys_tmp1330 = (w_sys_tmp1331 + r_run_k_11);
	assign w_sys_tmp1331 = 32'sh00000326;
	assign w_sys_tmp1335 = (w_sys_tmp1336 + r_run_k_11);
	assign w_sys_tmp1336 = 32'sh00000345;
	assign w_sys_tmp1340 = (w_sys_tmp1341 + r_run_k_11);
	assign w_sys_tmp1341 = 32'sh00000364;
	assign w_sys_tmp1345 = (w_sys_tmp1346 + r_run_k_11);
	assign w_sys_tmp1346 = 32'sh00000383;
	assign w_sys_tmp1350 = (w_sys_tmp1351 + r_run_k_11);
	assign w_sys_tmp1351 = 32'sh000003a2;
	assign w_sys_tmp1354 = (r_run_k_11 + w_sys_intOne);


	sub08
		sub08_inst(
			.i_fld_result_1_addr_0 (w_sub08_result_addr),
			.i_fld_result_1_datain_0 (w_sub08_result_datain),
			.o_fld_result_1_dataout_0 (w_sub08_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub08_result_r_w),
			.i_fld_u_0_addr_0 (w_sub08_u_addr),
			.i_fld_u_0_datain_0 (w_sub08_u_datain),
			.o_fld_u_0_dataout_0 (w_sub08_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub08_u_r_w),
			.o_run_busy (w_sub08_run_busy),
			.i_run_req (r_sub08_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub03
		sub03_inst(
			.i_fld_result_1_addr_0 (w_sub03_result_addr),
			.i_fld_result_1_datain_0 (w_sub03_result_datain),
			.o_fld_result_1_dataout_0 (w_sub03_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub03_result_r_w),
			.i_fld_u_0_addr_0 (w_sub03_u_addr),
			.i_fld_u_0_datain_0 (w_sub03_u_datain),
			.o_fld_u_0_dataout_0 (w_sub03_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub03_u_r_w),
			.o_run_busy (w_sub03_run_busy),
			.i_run_req (r_sub03_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub02
		sub02_inst(
			.i_fld_result_1_addr_0 (w_sub02_result_addr),
			.i_fld_result_1_datain_0 (w_sub02_result_datain),
			.o_fld_result_1_dataout_0 (w_sub02_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub02_result_r_w),
			.i_fld_u_0_addr_0 (w_sub02_u_addr),
			.i_fld_u_0_datain_0 (w_sub02_u_datain),
			.o_fld_u_0_dataout_0 (w_sub02_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub02_u_r_w),
			.o_run_busy (w_sub02_run_busy),
			.i_run_req (r_sub02_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub01
		sub01_inst(
			.i_fld_result_1_addr_0 (w_sub01_result_addr),
			.i_fld_result_1_datain_0 (w_sub01_result_datain),
			.o_fld_result_1_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub01_result_r_w),
			.i_fld_u_0_addr_0 (w_sub01_u_addr),
			.i_fld_u_0_datain_0 (w_sub01_u_datain),
			.o_fld_u_0_dataout_0 (w_sub01_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub01_u_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub00
		sub00_inst(
			.i_fld_result_1_addr_0 (w_sub00_result_addr),
			.i_fld_result_1_datain_0 (w_sub00_result_datain),
			.o_fld_result_1_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub00_result_r_w),
			.i_fld_u_0_addr_0 (w_sub00_u_addr),
			.i_fld_u_0_datain_0 (w_sub00_u_datain),
			.o_fld_u_0_dataout_0 (w_sub00_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub00_u_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub07
		sub07_inst(
			.i_fld_result_1_addr_0 (w_sub07_result_addr),
			.i_fld_result_1_datain_0 (w_sub07_result_datain),
			.o_fld_result_1_dataout_0 (w_sub07_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub07_result_r_w),
			.i_fld_u_0_addr_0 (w_sub07_u_addr),
			.i_fld_u_0_datain_0 (w_sub07_u_datain),
			.o_fld_u_0_dataout_0 (w_sub07_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub07_u_r_w),
			.o_run_busy (w_sub07_run_busy),
			.i_run_req (r_sub07_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub06
		sub06_inst(
			.i_fld_result_1_addr_0 (w_sub06_result_addr),
			.i_fld_result_1_datain_0 (w_sub06_result_datain),
			.o_fld_result_1_dataout_0 (w_sub06_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub06_result_r_w),
			.i_fld_u_0_addr_0 (w_sub06_u_addr),
			.i_fld_u_0_datain_0 (w_sub06_u_datain),
			.o_fld_u_0_dataout_0 (w_sub06_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub06_u_r_w),
			.o_run_busy (w_sub06_run_busy),
			.i_run_req (r_sub06_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub05
		sub05_inst(
			.i_fld_result_1_addr_0 (w_sub05_result_addr),
			.i_fld_result_1_datain_0 (w_sub05_result_datain),
			.o_fld_result_1_dataout_0 (w_sub05_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub05_result_r_w),
			.i_fld_u_0_addr_0 (w_sub05_u_addr),
			.i_fld_u_0_datain_0 (w_sub05_u_datain),
			.o_fld_u_0_dataout_0 (w_sub05_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub05_u_r_w),
			.o_run_busy (w_sub05_run_busy),
			.i_run_req (r_sub05_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub04
		sub04_inst(
			.i_fld_result_1_addr_0 (w_sub04_result_addr),
			.i_fld_result_1_datain_0 (w_sub04_result_datain),
			.o_fld_result_1_dataout_0 (w_sub04_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub04_result_r_w),
			.i_fld_u_0_addr_0 (w_sub04_u_addr),
			.i_fld_u_0_datain_0 (w_sub04_u_datain),
			.o_fld_u_0_dataout_0 (w_sub04_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub04_u_r_w),
			.o_run_busy (w_sub04_run_busy),
			.i_run_req (r_sub04_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(9), .WORDS(484) )
		dpram_u_0(
			.clk (clock),
			.ce_0 (w_fld_u_0_ce_0),
			.addr_0 (w_fld_u_0_addr_0),
			.datain_0 (w_fld_u_0_datain_0),
			.dataout_0 (w_fld_u_0_dataout_0),
			.r_w_0 (w_fld_u_0_r_w_0),
			.ce_1 (w_fld_u_0_ce_1),
			.addr_1 (r_fld_u_0_addr_1),
			.datain_1 (r_fld_u_0_datain_1),
			.dataout_1 (w_fld_u_0_dataout_1),
			.r_w_1 (r_fld_u_0_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(9), .WORDS(484) )
		dpram_uu_1(
			.clk (clock),
			.ce_0 (w_fld_uu_1_ce_0),
			.addr_0 (w_fld_uu_1_addr_0),
			.datain_0 (w_fld_uu_1_datain_0),
			.dataout_0 (w_fld_uu_1_dataout_0),
			.r_w_0 (w_fld_uu_1_r_w_0),
			.ce_1 (w_fld_uu_1_ce_1),
			.addr_1 (r_fld_uu_1_addr_1),
			.datain_1 (r_fld_uu_1_datain_1),
			.dataout_1 (w_fld_uu_1_dataout_1),
			.r_w_1 (r_fld_uu_1_r_w_1)
		);

	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h35: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 6'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_phase <= 6'h2;
						end

						6'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h4;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4) ? 6'h9 : 6'hf);

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'ha;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7) ? 6'hd : 6'h6);

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_run_phase <= 6'ha;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h10;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp94) ? 6'h14 : 6'h35);

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h10;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h15;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp97) ? 6'h18 : 6'h1a);

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1b)) begin
										r_sys_run_phase <= 6'h15;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h1b;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp254) ? 6'h1e : 6'h20);

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h47)) begin
										r_sys_run_phase <= 6'h1b;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h21;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp680) ? 6'h24 : 6'h25);

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h22)) begin
										r_sys_run_phase <= 6'h21;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_phase <= 6'h27;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								4'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_phase <= 6'h29;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h2a;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp884) ? 6'h2d : 6'h2f);

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3b)) begin
										r_sys_run_phase <= 6'h2a;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h30;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1190) ? 6'h33 : 6'h11);

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1f)) begin
										r_sys_run_phase <= 6'h30;

									end
								end

							endcase
						end

						6'h35: begin
							r_sys_run_phase <= 6'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 4'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1b)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h47)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h22)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3b)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1f)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 7'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h5)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h1a)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h46)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h47)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h21)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h22)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub00_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub01_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub02_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub03_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub04_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub05_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub06_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub07_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub08_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3a)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h3b)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h1e)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						6'h35: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_addr_1 <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp11[8:0] );

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h4) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp101[8:0] );

									end
									else
									if((r_sys_run_step==7'h1) || (r_sys_run_step==7'h5) || (r_sys_run_step==7'h9) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp105[8:0] );

									end
									else
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp114[8:0] );

									end
									else
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp109[8:0] );

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h36)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp583[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp289[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp421[8:0] );

									end
									else
									if((r_sys_run_step==7'h37)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp589[8:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp451[8:0] );

									end
									else
									if((r_sys_run_step==7'h29)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp505[8:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp385[8:0] );

									end
									else
									if((r_sys_run_step==7'h45)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp673[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp415[8:0] );

									end
									else
									if((r_sys_run_step==7'h33)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp565[8:0] );

									end
									else
									if((r_sys_run_step==7'h3d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp625[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp277[8:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp439[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp295[8:0] );

									end
									else
									if((r_sys_run_step==7'h25)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp481[8:0] );

									end
									else
									if((r_sys_run_step==7'h27)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp493[8:0] );

									end
									else
									if((r_sys_run_step==7'h22)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp463[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp265[8:0] );

									end
									else
									if((r_sys_run_step==7'h39) || (r_sys_run_step==7'h3b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp601[8:0] );

									end
									else
									if((r_sys_run_step==7'h32)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp559[8:0] );

									end
									else
									if((r_sys_run_step==7'h3f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp637[8:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp427[8:0] );

									end
									else
									if((r_sys_run_step==7'h2b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp517[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp379[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp313[8:0] );

									end
									else
									if((r_sys_run_step==7'h2e) || (r_sys_run_step==7'h30)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp535[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp361[8:0] );

									end
									else
									if((r_sys_run_step==7'h43)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp661[8:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp433[8:0] );

									end
									else
									if((r_sys_run_step==7'h42)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp655[8:0] );

									end
									else
									if((r_sys_run_step==7'h34)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp571[8:0] );

									end
									else
									if((r_sys_run_step==7'h16) || (r_sys_run_step==7'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp391[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp349[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp271[8:0] );

									end
									else
									if((r_sys_run_step==7'h44)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp667[8:0] );

									end
									else
									if((r_sys_run_step==7'h17) || (r_sys_run_step==7'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp397[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp307[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp373[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp283[8:0] );

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp457[8:0] );

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp577[8:0] );

									end
									else
									if((r_sys_run_step==7'h23)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp469[8:0] );

									end
									else
									if((r_sys_run_step==7'h2d) || (r_sys_run_step==7'h2f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp529[8:0] );

									end
									else
									if((r_sys_run_step==7'h40)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp643[8:0] );

									end
									else
									if((r_sys_run_step==7'h3e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp631[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp355[8:0] );

									end
									else
									if((r_sys_run_step==7'h28)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp499[8:0] );

									end
									else
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp319[8:0] );

									end
									else
									if((r_sys_run_step==7'h2c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp523[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp301[8:0] );

									end
									else
									if((r_sys_run_step==7'h24)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp475[8:0] );

									end
									else
									if((r_sys_run_step==7'h31)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp553[8:0] );

									end
									else
									if((r_sys_run_step==7'hb) || (r_sys_run_step==7'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp325[8:0] );

									end
									else
									if((r_sys_run_step==7'h38)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp595[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp367[8:0] );

									end
									else
									if((r_sys_run_step==7'h41)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp649[8:0] );

									end
									else
									if((r_sys_run_step==7'h26)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp487[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp259[8:0] );

									end
									else
									if((r_sys_run_step==7'h3a) || (r_sys_run_step==7'h3c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp607[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp343[8:0] );

									end
									else
									if((r_sys_run_step==7'h2a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp511[8:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp445[8:0] );

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp775[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp799[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp781[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp847[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp721[8:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp859[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp841[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp805[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp769[8:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp835[8:0] );

									end
									else
									if((r_sys_run_step==7'hb) || (r_sys_run_step==7'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp751[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp703[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp793[8:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp865[8:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp871[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp733[8:0] );

									end
									else
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp745[8:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp811[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp739[8:0] );

									end
									else
									if((r_sys_run_step==7'h16) || (r_sys_run_step==7'h17)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp817[8:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp877[8:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp829[8:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp853[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp709[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp685[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp787[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp727[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp715[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp697[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp691[8:0] );

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h15)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp994[8:0] );

									end
									else
									if((r_sys_run_step==7'h2c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1109[8:0] );

									end
									else
									if((r_sys_run_step==7'h25)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1074[8:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1034[8:0] );

									end
									else
									if((r_sys_run_step==7'h29)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1094[8:0] );

									end
									else
									if((r_sys_run_step==7'h23)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1064[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp984[8:0] );

									end
									else
									if((r_sys_run_step==7'h32)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1139[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp889[8:0] );

									end
									else
									if((r_sys_run_step==7'h37)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1164[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp964[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1019[8:0] );

									end
									else
									if((r_sys_run_step==7'h31)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1134[8:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1049[8:0] );

									end
									else
									if((r_sys_run_step==7'h26)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1079[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp959[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp931[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1024[8:0] );

									end
									else
									if((r_sys_run_step==7'h30)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1129[8:0] );

									end
									else
									if((r_sys_run_step==7'h33)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1144[8:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp954[8:0] );

									end
									else
									if((r_sys_run_step==7'h24)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1069[8:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1044[8:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1014[8:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1029[8:0] );

									end
									else
									if((r_sys_run_step==7'h28)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1089[8:0] );

									end
									else
									if((r_sys_run_step==7'h3a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1179[8:0] );

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1004[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp925[8:0] );

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1154[8:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp943[8:0] );

									end
									else
									if((r_sys_run_step==7'h39)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1174[8:0] );

									end
									else
									if((r_sys_run_step==7'h2e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1119[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp913[8:0] );

									end
									else
									if((r_sys_run_step==7'h34)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1149[8:0] );

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp999[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp895[8:0] );

									end
									else
									if((r_sys_run_step==7'h3b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1184[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp989[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp979[8:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp937[8:0] );

									end
									else
									if((r_sys_run_step==7'h22)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1059[8:0] );

									end
									else
									if((r_sys_run_step==7'h2f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1124[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp901[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp974[8:0] );

									end
									else
									if((r_sys_run_step==7'h2d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1114[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp907[8:0] );

									end
									else
									if((r_sys_run_step==7'h2b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1104[8:0] );

									end
									else
									if((r_sys_run_step==7'h38)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1169[8:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1009[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp919[8:0] );

									end
									else
									if((r_sys_run_step==7'h27)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1084[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp969[8:0] );

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1054[8:0] );

									end
									else
									if((r_sys_run_step==7'h2a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1099[8:0] );

									end
									else
									if((r_sys_run_step==7'h36)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1159[8:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1039[8:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp949[8:0] );

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1265[8:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1350[8:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1249[8:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1340[8:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1255[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1225[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1231[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1270[8:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1315[8:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1300[8:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1260[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1219[8:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1243[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1290[8:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1335[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1280[8:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1345[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1237[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1207[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1330[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1195[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1295[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1201[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1213[8:0] );

									end
									else
									if((r_sys_run_step==7'h16) || (r_sys_run_step==7'h17)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1305[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1285[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1275[8:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1320[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1325[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp14;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1a)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp112;

									end
									else
									if((r_sys_run_step==7'h1) || (r_sys_run_step==7'h3) || (r_sys_run_step==7'h5) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'h9) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h1b)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp107;

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h4) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h18)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp103;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h36)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp30_float;

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp23_float;

									end
									else
									if((r_sys_run_step==7'h2f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp32_float;

									end
									else
									if((r_sys_run_step==7'h30)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==7'h34)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp41_float;

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp37_float;

									end
									else
									if((r_sys_run_step==7'h25)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp38_float;

									end
									else
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'hb)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp891;

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==7'h29)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp44_float;

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp18_float;

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp42_float;

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp45_float;

									end
									else
									if((r_sys_run_step==7'h37)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp26_float;

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==7'h2a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp39_float;

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp33_float;

									end
									else
									if((r_sys_run_step==7'h2c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp31_float;

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp24_float;

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp47_float;

									end
									else
									if((r_sys_run_step==7'h32)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp34_float;

									end
									else
									if((r_sys_run_step==7'h24)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp20_float;

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp19_float;

									end
									else
									if((r_sys_run_step==7'h2e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp22_float;

									end
									else
									if((r_sys_run_step==7'h28)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==7'h3b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==7'h2b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp35_float;

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp36_float;

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp28_float;

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp40_float;

									end
									else
									if((r_sys_run_step==7'h2d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp27_float;

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==7'h27)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==7'h31)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==7'h22)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp29_float;

									end
									else
									if((r_sys_run_step==7'h38)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp21_float;

									end
									else
									if((r_sys_run_step==7'h3a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==7'h26)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==7'h33)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp46_float;

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp43_float;

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==7'h23)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp25_float;

									end
									else
									if((r_sys_run_step==7'h39)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp14_float;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'hc) || (r_sys_run_step==7'h16)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp19_float;

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp2_float;

									end
									else
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'hb)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp1197;

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp14_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h1b)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h45)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h20)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h3b)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h1f)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h35: begin
							r_fld_u_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_uu_1_addr_1 <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_uu_1_addr_1 <= $signed( w_sys_tmp16[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_uu_1_datain_1 <= w_sys_tmp14;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_uu_1_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_uu_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h35: begin
							r_fld_uu_1_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h4: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_11 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_11 <= w_sys_tmp6;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_11 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h47)) begin
										r_run_k_11 <= w_sys_tmp678;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_11 <= w_sys_tmp679;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h22)) begin
										r_run_k_11 <= w_sys_tmp882;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_11 <= w_sys_tmp883;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3b)) begin
										r_run_k_11 <= w_sys_tmp1188;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_11 <= w_sys_tmp1189;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1f)) begin
										r_run_k_11 <= w_sys_tmp1354;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_12 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_12 <= w_sys_tmp21;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_12 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h4) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h18)) begin
										r_run_j_12 <= w_sys_tmp121;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_n_13 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_n_13 <= w_sys_tmp96;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_mx_14 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_my_15 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_nlast_16 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_17 <= r_run_j_12;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_17 <= w_sys_tmp20;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_18 <= r_run_j_12;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h1b)) begin
										r_run_copy0_j_18 <= w_sys_tmp118;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_19 <= r_run_j_12;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1a)) begin
										r_run_copy1_j_19 <= w_sys_tmp119;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy2_j_20 <= r_run_j_12;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1) || (r_sys_run_step==7'h5) || (r_sys_run_step==7'h9) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h19)) begin
										r_run_copy2_j_20 <= w_sys_tmp120;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub08_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub08_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1b)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp835[9:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp847[9:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp859[9:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp817[9:0] );

									end
									else
									if((r_sys_run_step==7'h22)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp877[9:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp829[9:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp853[9:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp865[9:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp841[9:0] );

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp871[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h19<=r_sys_run_step && r_sys_run_step<=7'h22)) begin
										r_sub08_u_datain <= w_sys_tmp687;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h19<=r_sys_run_step && r_sys_run_step<=7'h22)) begin
										r_sub08_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub08_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1350[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1345[9:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1305[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1340[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1320[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1330[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1335[9:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1315[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1325[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub08_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h2: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h29)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp493[9:0] );

									end
									else
									if((r_sys_run_step==7'h27)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp481[9:0] );

									end
									else
									if((r_sys_run_step==7'h25)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp469[9:0] );

									end
									else
									if((r_sys_run_step==7'h26)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp475[9:0] );

									end
									else
									if((r_sys_run_step==7'h2f)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp529[9:0] );

									end
									else
									if((r_sys_run_step==7'h2d)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp517[9:0] );

									end
									else
									if((r_sys_run_step==7'h28)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp487[9:0] );

									end
									else
									if((r_sys_run_step==7'h2b)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp505[9:0] );

									end
									else
									if((r_sys_run_step==7'h30)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp535[9:0] );

									end
									else
									if((r_sys_run_step==7'h2a)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp499[9:0] );

									end
									else
									if((r_sys_run_step==7'h2c)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp511[9:0] );

									end
									else
									if((r_sys_run_step==7'h2e)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp523[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h25<=r_sys_run_step && r_sys_run_step<=7'h30)) begin
										r_sub03_u_datain <= w_sys_tmp261;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h25<=r_sys_run_step && r_sys_run_step<=7'h30)) begin
										r_sub03_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub03_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1064[9:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1049[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1079[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1084[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1059[9:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1044[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1074[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1054[9:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1089[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1069[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h9)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub03_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h23)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp457[9:0] );

									end
									else
									if((r_sys_run_step==7'h24)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp463[9:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp433[9:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp427[9:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp415[9:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp391[9:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp421[9:0] );

									end
									else
									if((r_sys_run_step==7'h22)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp451[9:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp397[9:0] );

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp445[9:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp439[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h1a<=r_sys_run_step && r_sys_run_step<=7'h24)) begin
										r_sub02_u_datain <= w_sys_tmp261;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h1a<=r_sys_run_step && r_sys_run_step<=7'h24)) begin
										r_sub02_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub02_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1009[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1024[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1014[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1029[9:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp999[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1039[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1034[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1019[9:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1004[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub02_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h17)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp385[9:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp367[9:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp391[9:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp355[9:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp349[9:0] );

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp379[9:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp325[9:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp343[9:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp397[9:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp361[9:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp319[9:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp373[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h19)) begin
										r_sub01_u_datain <= w_sys_tmp261;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h19)) begin
										r_sub01_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub01_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp994[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp989[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp979[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp984[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp959[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp969[9:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp954[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp964[9:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp949[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp974[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h9)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h6: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp301[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp295[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp289[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp265[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp271[9:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp325[9:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp313[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp259[9:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp319[9:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp307[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp277[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp283[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub00_u_datain <= w_sys_tmp261;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub00_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub00_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp907[9:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp943[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp919[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp937[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp913[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp931[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp925[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp901[9:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp889[9:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp895[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h9)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h5: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub07_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub07_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h11)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp775[9:0] );

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp805[9:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp799[9:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp781[9:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp745[9:0] );

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp811[9:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp787[9:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp769[9:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp751[9:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp817[9:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp793[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h18)) begin
										r_sub07_u_datain <= w_sys_tmp687;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h18)) begin
										r_sub07_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub07_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1265[9:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1300[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1295[9:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1260[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1280[9:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1305[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1290[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1285[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1275[9:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1255[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1270[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'ha)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub07_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h4: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub06_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub06_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp733[9:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp745[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp685[9:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp739[9:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp727[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp721[9:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp751[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp703[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp715[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp709[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp697[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp691[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub06_u_datain <= w_sys_tmp687;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub06_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub06_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1195[9:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1201[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1219[9:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1249[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1243[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1213[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1237[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1207[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1225[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1231[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h9)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub06_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h3: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub05_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub05_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h41)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp637[9:0] );

									end
									else
									if((r_sys_run_step==7'h44)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp655[9:0] );

									end
									else
									if((r_sys_run_step==7'h47)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp673[9:0] );

									end
									else
									if((r_sys_run_step==7'h43)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp649[9:0] );

									end
									else
									if((r_sys_run_step==7'h42)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp643[9:0] );

									end
									else
									if((r_sys_run_step==7'h40)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp631[9:0] );

									end
									else
									if((r_sys_run_step==7'h3e)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp607[9:0] );

									end
									else
									if((r_sys_run_step==7'h46)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp667[9:0] );

									end
									else
									if((r_sys_run_step==7'h3f)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp625[9:0] );

									end
									else
									if((r_sys_run_step==7'h3d)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp601[9:0] );

									end
									else
									if((r_sys_run_step==7'h45)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp661[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h3d<=r_sys_run_step && r_sys_run_step<=7'h47)) begin
										r_sub05_u_datain <= w_sys_tmp261;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h3d<=r_sys_run_step && r_sys_run_step<=7'h47)) begin
										r_sub05_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub05_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1169[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1174[9:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1149[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1154[9:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1144[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1164[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1159[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1179[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1184[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub05_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h7: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub04_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub04_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h38)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp583[9:0] );

									end
									else
									if((r_sys_run_step==7'h37)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp577[9:0] );

									end
									else
									if((r_sys_run_step==7'h34)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp559[9:0] );

									end
									else
									if((r_sys_run_step==7'h3a)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp595[9:0] );

									end
									else
									if((r_sys_run_step==7'h36)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp571[9:0] );

									end
									else
									if((r_sys_run_step==7'h33)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp553[9:0] );

									end
									else
									if((r_sys_run_step==7'h31)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp529[9:0] );

									end
									else
									if((r_sys_run_step==7'h39)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp589[9:0] );

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp565[9:0] );

									end
									else
									if((r_sys_run_step==7'h3c)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp607[9:0] );

									end
									else
									if((r_sys_run_step==7'h32)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp535[9:0] );

									end
									else
									if((r_sys_run_step==7'h3b)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp601[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h31<=r_sys_run_step && r_sys_run_step<=7'h3c)) begin
										r_sub04_u_datain <= w_sys_tmp261;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h31<=r_sys_run_step && r_sys_run_step<=7'h3c)) begin
										r_sub04_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub04_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1134[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1104[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1119[9:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1139[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1124[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1109[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1129[9:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1099[9:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1094[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1114[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h9)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub04_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'hb)) begin
										r_sys_tmp0_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'hb)) begin
										r_sys_tmp0_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'hb)) begin
										r_sys_tmp1_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sys_tmp1_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'hb)) begin
										r_sys_tmp2_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sys_tmp2_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sys_tmp3_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sys_tmp3_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sys_tmp4_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sys_tmp4_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sys_tmp5_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_tmp5_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sys_tmp6_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_tmp6_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sys_tmp7_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sys_tmp7_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sys_tmp8_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sys_tmp8_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sys_tmp9_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_tmp9_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sys_tmp10_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_tmp10_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sys_tmp11_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp11_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sys_tmp12_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp12_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_tmp13_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp13_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_tmp14_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp14_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_tmp15_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp15_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_tmp16_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp16_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_tmp17_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp17_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sys_tmp18_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sys_tmp19_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'hc)) begin
										r_sys_tmp19_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sys_tmp20_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sys_tmp21_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sys_tmp22_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_tmp23_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_tmp24_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_tmp25_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_tmp26_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_tmp27_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp28_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp29_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp30_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp31_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp32_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp33_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp34_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp35_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp36_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp37_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp38_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp39_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp40_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp41_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp42_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp43_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp44_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp45_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp46_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp47_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
