/*
TimeStamp:	2016/6/17		18:46
*/


module P3_2dim(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy,	
	output signed  [31:0] o_run_return	
);

	reg  signed [31:0] r_ip_DivInt_dividend_0;
	reg  signed [31:0] r_ip_DivInt_divisor_0;
	wire signed [31:0] w_ip_DivInt_quotient_0;
	wire signed [31:0] w_ip_DivInt_fractional_0;
	reg         [31:0] r_ip_AddFloat_portA_0;
	reg         [31:0] r_ip_AddFloat_portB_0;
	wire        [31:0] w_ip_AddFloat_result_0;
	reg         [31:0] r_ip_MultFloat_multiplicand_0;
	reg         [31:0] r_ip_MultFloat_multiplier_0;
	wire        [31:0] w_ip_MultFloat_product_0;
	reg  signed [31:0] r_ip_FixedToFloat_fixed_0;
	wire        [31:0] w_ip_FixedToFloat_floating_0;
	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [31:0] r_sys_run_return;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 6:0] r_sys_run_phase;
	reg         [ 4:0] r_sys_run_stage;
	reg         [ 6:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 4:0] w_sys_run_stage_p1;
	wire        [ 6:0] w_sys_run_step_p1;
	wire signed [ 8:0] w_fld_T_0_addr_0;
	wire        [31:0] w_fld_T_0_datain_0;
	wire        [31:0] w_fld_T_0_dataout_0;
	wire               w_fld_T_0_r_w_0;
	wire               w_fld_T_0_ce_0;
	reg  signed [ 8:0] r_fld_T_0_addr_1;
	reg         [31:0] r_fld_T_0_datain_1;
	wire        [31:0] w_fld_T_0_dataout_1;
	reg                r_fld_T_0_r_w_1;
	wire               w_fld_T_0_ce_1;
	wire signed [ 8:0] w_fld_TT_1_addr_0;
	wire        [31:0] w_fld_TT_1_datain_0;
	wire        [31:0] w_fld_TT_1_dataout_0;
	wire               w_fld_TT_1_r_w_0;
	wire               w_fld_TT_1_ce_0;
	reg  signed [ 8:0] r_fld_TT_1_addr_1;
	reg         [31:0] r_fld_TT_1_datain_1;
	wire        [31:0] w_fld_TT_1_dataout_1;
	reg                r_fld_TT_1_r_w_1;
	wire               w_fld_TT_1_ce_1;
	wire signed [ 8:0] w_fld_U_2_addr_0;
	wire        [31:0] w_fld_U_2_datain_0;
	wire        [31:0] w_fld_U_2_dataout_0;
	wire               w_fld_U_2_r_w_0;
	wire               w_fld_U_2_ce_0;
	reg  signed [ 8:0] r_fld_U_2_addr_1;
	reg         [31:0] r_fld_U_2_datain_1;
	wire        [31:0] w_fld_U_2_dataout_1;
	reg                r_fld_U_2_r_w_1;
	wire               w_fld_U_2_ce_1;
	wire signed [ 8:0] w_fld_V_3_addr_0;
	wire        [31:0] w_fld_V_3_datain_0;
	wire        [31:0] w_fld_V_3_dataout_0;
	wire               w_fld_V_3_r_w_0;
	wire               w_fld_V_3_ce_0;
	reg  signed [ 8:0] r_fld_V_3_addr_1;
	reg         [31:0] r_fld_V_3_datain_1;
	wire        [31:0] w_fld_V_3_dataout_1;
	reg                r_fld_V_3_r_w_1;
	wire               w_fld_V_3_ce_1;
	reg  signed [31:0] r_run_k_29;
	reg  signed [31:0] r_run_j_30;
	reg  signed [31:0] r_run_n_31;
	reg  signed [31:0] r_run_mx_32;
	reg  signed [31:0] r_run_my_33;
	reg         [31:0] r_run_dt_34;
	reg         [31:0] r_run_dx_35;
	reg         [31:0] r_run_dy_36;
	reg         [31:0] r_run_r1_37;
	reg         [31:0] r_run_r2_38;
	reg         [31:0] r_run_r3_39;
	reg         [31:0] r_run_r4_40;
	reg         [31:0] r_run_YY_41;
	reg  signed [31:0] r_run_kx_42;
	reg  signed [31:0] r_run_ky_43;
	reg  signed [31:0] r_run_nlast_44;
	reg  signed [31:0] r_run_copy0_j_45;
	reg  signed [31:0] r_run_copy1_j_46;
	reg  signed [31:0] r_run_copy2_j_47;
	reg  signed [31:0] r_run_copy0_j_48;
	reg                r_sub19_run_req;
	wire               w_sub19_run_busy;
	wire signed [ 8:0] w_sub19_T_addr;
	reg  signed [ 8:0] r_sub19_T_addr;
	wire        [31:0] w_sub19_T_datain;
	reg         [31:0] r_sub19_T_datain;
	wire        [31:0] w_sub19_T_dataout;
	wire               w_sub19_T_r_w;
	reg                r_sub19_T_r_w;
	wire signed [ 8:0] w_sub19_V_addr;
	reg  signed [ 8:0] r_sub19_V_addr;
	wire        [31:0] w_sub19_V_datain;
	reg         [31:0] r_sub19_V_datain;
	wire        [31:0] w_sub19_V_dataout;
	wire               w_sub19_V_r_w;
	reg                r_sub19_V_r_w;
	wire signed [ 8:0] w_sub19_U_addr;
	reg  signed [ 8:0] r_sub19_U_addr;
	wire        [31:0] w_sub19_U_datain;
	reg         [31:0] r_sub19_U_datain;
	wire        [31:0] w_sub19_U_dataout;
	wire               w_sub19_U_r_w;
	reg                r_sub19_U_r_w;
	wire signed [ 8:0] w_sub19_result_addr;
	reg  signed [ 8:0] r_sub19_result_addr;
	wire        [31:0] w_sub19_result_datain;
	reg         [31:0] r_sub19_result_datain;
	wire        [31:0] w_sub19_result_dataout;
	wire               w_sub19_result_r_w;
	reg                r_sub19_result_r_w;
	reg                r_sub09_run_req;
	wire               w_sub09_run_busy;
	wire signed [ 8:0] w_sub09_T_addr;
	reg  signed [ 8:0] r_sub09_T_addr;
	wire        [31:0] w_sub09_T_datain;
	reg         [31:0] r_sub09_T_datain;
	wire        [31:0] w_sub09_T_dataout;
	wire               w_sub09_T_r_w;
	reg                r_sub09_T_r_w;
	wire signed [ 8:0] w_sub09_V_addr;
	reg  signed [ 8:0] r_sub09_V_addr;
	wire        [31:0] w_sub09_V_datain;
	reg         [31:0] r_sub09_V_datain;
	wire        [31:0] w_sub09_V_dataout;
	wire               w_sub09_V_r_w;
	reg                r_sub09_V_r_w;
	wire signed [ 8:0] w_sub09_U_addr;
	reg  signed [ 8:0] r_sub09_U_addr;
	wire        [31:0] w_sub09_U_datain;
	reg         [31:0] r_sub09_U_datain;
	wire        [31:0] w_sub09_U_dataout;
	wire               w_sub09_U_r_w;
	reg                r_sub09_U_r_w;
	wire signed [ 8:0] w_sub09_result_addr;
	reg  signed [ 8:0] r_sub09_result_addr;
	wire        [31:0] w_sub09_result_datain;
	reg         [31:0] r_sub09_result_datain;
	wire        [31:0] w_sub09_result_dataout;
	wire               w_sub09_result_r_w;
	reg                r_sub09_result_r_w;
	reg                r_sub08_run_req;
	wire               w_sub08_run_busy;
	wire signed [ 8:0] w_sub08_T_addr;
	reg  signed [ 8:0] r_sub08_T_addr;
	wire        [31:0] w_sub08_T_datain;
	reg         [31:0] r_sub08_T_datain;
	wire        [31:0] w_sub08_T_dataout;
	wire               w_sub08_T_r_w;
	reg                r_sub08_T_r_w;
	wire signed [ 8:0] w_sub08_V_addr;
	reg  signed [ 8:0] r_sub08_V_addr;
	wire        [31:0] w_sub08_V_datain;
	reg         [31:0] r_sub08_V_datain;
	wire        [31:0] w_sub08_V_dataout;
	wire               w_sub08_V_r_w;
	reg                r_sub08_V_r_w;
	wire signed [ 8:0] w_sub08_U_addr;
	reg  signed [ 8:0] r_sub08_U_addr;
	wire        [31:0] w_sub08_U_datain;
	reg         [31:0] r_sub08_U_datain;
	wire        [31:0] w_sub08_U_dataout;
	wire               w_sub08_U_r_w;
	reg                r_sub08_U_r_w;
	wire signed [ 8:0] w_sub08_result_addr;
	reg  signed [ 8:0] r_sub08_result_addr;
	wire        [31:0] w_sub08_result_datain;
	reg         [31:0] r_sub08_result_datain;
	wire        [31:0] w_sub08_result_dataout;
	wire               w_sub08_result_r_w;
	reg                r_sub08_result_r_w;
	reg                r_sub24_run_req;
	wire               w_sub24_run_busy;
	wire signed [ 8:0] w_sub24_T_addr;
	reg  signed [ 8:0] r_sub24_T_addr;
	wire        [31:0] w_sub24_T_datain;
	reg         [31:0] r_sub24_T_datain;
	wire        [31:0] w_sub24_T_dataout;
	wire               w_sub24_T_r_w;
	reg                r_sub24_T_r_w;
	wire signed [ 8:0] w_sub24_V_addr;
	reg  signed [ 8:0] r_sub24_V_addr;
	wire        [31:0] w_sub24_V_datain;
	reg         [31:0] r_sub24_V_datain;
	wire        [31:0] w_sub24_V_dataout;
	wire               w_sub24_V_r_w;
	reg                r_sub24_V_r_w;
	wire signed [ 8:0] w_sub24_U_addr;
	reg  signed [ 8:0] r_sub24_U_addr;
	wire        [31:0] w_sub24_U_datain;
	reg         [31:0] r_sub24_U_datain;
	wire        [31:0] w_sub24_U_dataout;
	wire               w_sub24_U_r_w;
	reg                r_sub24_U_r_w;
	wire signed [ 8:0] w_sub24_result_addr;
	reg  signed [ 8:0] r_sub24_result_addr;
	wire        [31:0] w_sub24_result_datain;
	reg         [31:0] r_sub24_result_datain;
	wire        [31:0] w_sub24_result_dataout;
	wire               w_sub24_result_r_w;
	reg                r_sub24_result_r_w;
	reg                r_sub22_run_req;
	wire               w_sub22_run_busy;
	wire signed [ 8:0] w_sub22_T_addr;
	reg  signed [ 8:0] r_sub22_T_addr;
	wire        [31:0] w_sub22_T_datain;
	reg         [31:0] r_sub22_T_datain;
	wire        [31:0] w_sub22_T_dataout;
	wire               w_sub22_T_r_w;
	reg                r_sub22_T_r_w;
	wire signed [ 8:0] w_sub22_V_addr;
	reg  signed [ 8:0] r_sub22_V_addr;
	wire        [31:0] w_sub22_V_datain;
	reg         [31:0] r_sub22_V_datain;
	wire        [31:0] w_sub22_V_dataout;
	wire               w_sub22_V_r_w;
	reg                r_sub22_V_r_w;
	wire signed [ 8:0] w_sub22_U_addr;
	reg  signed [ 8:0] r_sub22_U_addr;
	wire        [31:0] w_sub22_U_datain;
	reg         [31:0] r_sub22_U_datain;
	wire        [31:0] w_sub22_U_dataout;
	wire               w_sub22_U_r_w;
	reg                r_sub22_U_r_w;
	wire signed [ 8:0] w_sub22_result_addr;
	reg  signed [ 8:0] r_sub22_result_addr;
	wire        [31:0] w_sub22_result_datain;
	reg         [31:0] r_sub22_result_datain;
	wire        [31:0] w_sub22_result_dataout;
	wire               w_sub22_result_r_w;
	reg                r_sub22_result_r_w;
	reg                r_sub23_run_req;
	wire               w_sub23_run_busy;
	wire signed [ 8:0] w_sub23_T_addr;
	reg  signed [ 8:0] r_sub23_T_addr;
	wire        [31:0] w_sub23_T_datain;
	reg         [31:0] r_sub23_T_datain;
	wire        [31:0] w_sub23_T_dataout;
	wire               w_sub23_T_r_w;
	reg                r_sub23_T_r_w;
	wire signed [ 8:0] w_sub23_V_addr;
	reg  signed [ 8:0] r_sub23_V_addr;
	wire        [31:0] w_sub23_V_datain;
	reg         [31:0] r_sub23_V_datain;
	wire        [31:0] w_sub23_V_dataout;
	wire               w_sub23_V_r_w;
	reg                r_sub23_V_r_w;
	wire signed [ 8:0] w_sub23_U_addr;
	reg  signed [ 8:0] r_sub23_U_addr;
	wire        [31:0] w_sub23_U_datain;
	reg         [31:0] r_sub23_U_datain;
	wire        [31:0] w_sub23_U_dataout;
	wire               w_sub23_U_r_w;
	reg                r_sub23_U_r_w;
	wire signed [ 8:0] w_sub23_result_addr;
	reg  signed [ 8:0] r_sub23_result_addr;
	wire        [31:0] w_sub23_result_datain;
	reg         [31:0] r_sub23_result_datain;
	wire        [31:0] w_sub23_result_dataout;
	wire               w_sub23_result_r_w;
	reg                r_sub23_result_r_w;
	reg                r_sub12_run_req;
	wire               w_sub12_run_busy;
	wire signed [ 8:0] w_sub12_T_addr;
	reg  signed [ 8:0] r_sub12_T_addr;
	wire        [31:0] w_sub12_T_datain;
	reg         [31:0] r_sub12_T_datain;
	wire        [31:0] w_sub12_T_dataout;
	wire               w_sub12_T_r_w;
	reg                r_sub12_T_r_w;
	wire signed [ 8:0] w_sub12_V_addr;
	reg  signed [ 8:0] r_sub12_V_addr;
	wire        [31:0] w_sub12_V_datain;
	reg         [31:0] r_sub12_V_datain;
	wire        [31:0] w_sub12_V_dataout;
	wire               w_sub12_V_r_w;
	reg                r_sub12_V_r_w;
	wire signed [ 8:0] w_sub12_U_addr;
	reg  signed [ 8:0] r_sub12_U_addr;
	wire        [31:0] w_sub12_U_datain;
	reg         [31:0] r_sub12_U_datain;
	wire        [31:0] w_sub12_U_dataout;
	wire               w_sub12_U_r_w;
	reg                r_sub12_U_r_w;
	wire signed [ 8:0] w_sub12_result_addr;
	reg  signed [ 8:0] r_sub12_result_addr;
	wire        [31:0] w_sub12_result_datain;
	reg         [31:0] r_sub12_result_datain;
	wire        [31:0] w_sub12_result_dataout;
	wire               w_sub12_result_r_w;
	reg                r_sub12_result_r_w;
	reg                r_sub03_run_req;
	wire               w_sub03_run_busy;
	wire signed [ 8:0] w_sub03_T_addr;
	reg  signed [ 8:0] r_sub03_T_addr;
	wire        [31:0] w_sub03_T_datain;
	reg         [31:0] r_sub03_T_datain;
	wire        [31:0] w_sub03_T_dataout;
	wire               w_sub03_T_r_w;
	reg                r_sub03_T_r_w;
	wire signed [ 8:0] w_sub03_V_addr;
	reg  signed [ 8:0] r_sub03_V_addr;
	wire        [31:0] w_sub03_V_datain;
	reg         [31:0] r_sub03_V_datain;
	wire        [31:0] w_sub03_V_dataout;
	wire               w_sub03_V_r_w;
	reg                r_sub03_V_r_w;
	wire signed [ 8:0] w_sub03_U_addr;
	reg  signed [ 8:0] r_sub03_U_addr;
	wire        [31:0] w_sub03_U_datain;
	reg         [31:0] r_sub03_U_datain;
	wire        [31:0] w_sub03_U_dataout;
	wire               w_sub03_U_r_w;
	reg                r_sub03_U_r_w;
	wire signed [ 8:0] w_sub03_result_addr;
	reg  signed [ 8:0] r_sub03_result_addr;
	wire        [31:0] w_sub03_result_datain;
	reg         [31:0] r_sub03_result_datain;
	wire        [31:0] w_sub03_result_dataout;
	wire               w_sub03_result_r_w;
	reg                r_sub03_result_r_w;
	reg                r_sub02_run_req;
	wire               w_sub02_run_busy;
	wire signed [ 8:0] w_sub02_T_addr;
	reg  signed [ 8:0] r_sub02_T_addr;
	wire        [31:0] w_sub02_T_datain;
	reg         [31:0] r_sub02_T_datain;
	wire        [31:0] w_sub02_T_dataout;
	wire               w_sub02_T_r_w;
	reg                r_sub02_T_r_w;
	wire signed [ 8:0] w_sub02_V_addr;
	reg  signed [ 8:0] r_sub02_V_addr;
	wire        [31:0] w_sub02_V_datain;
	reg         [31:0] r_sub02_V_datain;
	wire        [31:0] w_sub02_V_dataout;
	wire               w_sub02_V_r_w;
	reg                r_sub02_V_r_w;
	wire signed [ 8:0] w_sub02_U_addr;
	reg  signed [ 8:0] r_sub02_U_addr;
	wire        [31:0] w_sub02_U_datain;
	reg         [31:0] r_sub02_U_datain;
	wire        [31:0] w_sub02_U_dataout;
	wire               w_sub02_U_r_w;
	reg                r_sub02_U_r_w;
	wire signed [ 8:0] w_sub02_result_addr;
	reg  signed [ 8:0] r_sub02_result_addr;
	wire        [31:0] w_sub02_result_datain;
	reg         [31:0] r_sub02_result_datain;
	wire        [31:0] w_sub02_result_dataout;
	wire               w_sub02_result_r_w;
	reg                r_sub02_result_r_w;
	reg                r_sub11_run_req;
	wire               w_sub11_run_busy;
	wire signed [ 8:0] w_sub11_T_addr;
	reg  signed [ 8:0] r_sub11_T_addr;
	wire        [31:0] w_sub11_T_datain;
	reg         [31:0] r_sub11_T_datain;
	wire        [31:0] w_sub11_T_dataout;
	wire               w_sub11_T_r_w;
	reg                r_sub11_T_r_w;
	wire signed [ 8:0] w_sub11_V_addr;
	reg  signed [ 8:0] r_sub11_V_addr;
	wire        [31:0] w_sub11_V_datain;
	reg         [31:0] r_sub11_V_datain;
	wire        [31:0] w_sub11_V_dataout;
	wire               w_sub11_V_r_w;
	reg                r_sub11_V_r_w;
	wire signed [ 8:0] w_sub11_U_addr;
	reg  signed [ 8:0] r_sub11_U_addr;
	wire        [31:0] w_sub11_U_datain;
	reg         [31:0] r_sub11_U_datain;
	wire        [31:0] w_sub11_U_dataout;
	wire               w_sub11_U_r_w;
	reg                r_sub11_U_r_w;
	wire signed [ 8:0] w_sub11_result_addr;
	reg  signed [ 8:0] r_sub11_result_addr;
	wire        [31:0] w_sub11_result_datain;
	reg         [31:0] r_sub11_result_datain;
	wire        [31:0] w_sub11_result_dataout;
	wire               w_sub11_result_r_w;
	reg                r_sub11_result_r_w;
	reg                r_sub14_run_req;
	wire               w_sub14_run_busy;
	wire signed [ 8:0] w_sub14_T_addr;
	reg  signed [ 8:0] r_sub14_T_addr;
	wire        [31:0] w_sub14_T_datain;
	reg         [31:0] r_sub14_T_datain;
	wire        [31:0] w_sub14_T_dataout;
	wire               w_sub14_T_r_w;
	reg                r_sub14_T_r_w;
	wire signed [ 8:0] w_sub14_V_addr;
	reg  signed [ 8:0] r_sub14_V_addr;
	wire        [31:0] w_sub14_V_datain;
	reg         [31:0] r_sub14_V_datain;
	wire        [31:0] w_sub14_V_dataout;
	wire               w_sub14_V_r_w;
	reg                r_sub14_V_r_w;
	wire signed [ 8:0] w_sub14_U_addr;
	reg  signed [ 8:0] r_sub14_U_addr;
	wire        [31:0] w_sub14_U_datain;
	reg         [31:0] r_sub14_U_datain;
	wire        [31:0] w_sub14_U_dataout;
	wire               w_sub14_U_r_w;
	reg                r_sub14_U_r_w;
	wire signed [ 8:0] w_sub14_result_addr;
	reg  signed [ 8:0] r_sub14_result_addr;
	wire        [31:0] w_sub14_result_datain;
	reg         [31:0] r_sub14_result_datain;
	wire        [31:0] w_sub14_result_dataout;
	wire               w_sub14_result_r_w;
	reg                r_sub14_result_r_w;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [ 8:0] w_sub01_T_addr;
	reg  signed [ 8:0] r_sub01_T_addr;
	wire        [31:0] w_sub01_T_datain;
	reg         [31:0] r_sub01_T_datain;
	wire        [31:0] w_sub01_T_dataout;
	wire               w_sub01_T_r_w;
	reg                r_sub01_T_r_w;
	wire signed [ 8:0] w_sub01_V_addr;
	reg  signed [ 8:0] r_sub01_V_addr;
	wire        [31:0] w_sub01_V_datain;
	reg         [31:0] r_sub01_V_datain;
	wire        [31:0] w_sub01_V_dataout;
	wire               w_sub01_V_r_w;
	reg                r_sub01_V_r_w;
	wire signed [ 8:0] w_sub01_U_addr;
	reg  signed [ 8:0] r_sub01_U_addr;
	wire        [31:0] w_sub01_U_datain;
	reg         [31:0] r_sub01_U_datain;
	wire        [31:0] w_sub01_U_dataout;
	wire               w_sub01_U_r_w;
	reg                r_sub01_U_r_w;
	wire signed [ 8:0] w_sub01_result_addr;
	reg  signed [ 8:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [ 8:0] w_sub00_T_addr;
	reg  signed [ 8:0] r_sub00_T_addr;
	wire        [31:0] w_sub00_T_datain;
	reg         [31:0] r_sub00_T_datain;
	wire        [31:0] w_sub00_T_dataout;
	wire               w_sub00_T_r_w;
	reg                r_sub00_T_r_w;
	wire signed [ 8:0] w_sub00_V_addr;
	reg  signed [ 8:0] r_sub00_V_addr;
	wire        [31:0] w_sub00_V_datain;
	reg         [31:0] r_sub00_V_datain;
	wire        [31:0] w_sub00_V_dataout;
	wire               w_sub00_V_r_w;
	reg                r_sub00_V_r_w;
	wire signed [ 8:0] w_sub00_U_addr;
	reg  signed [ 8:0] r_sub00_U_addr;
	wire        [31:0] w_sub00_U_datain;
	reg         [31:0] r_sub00_U_datain;
	wire        [31:0] w_sub00_U_dataout;
	wire               w_sub00_U_r_w;
	reg                r_sub00_U_r_w;
	wire signed [ 8:0] w_sub00_result_addr;
	reg  signed [ 8:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	reg                r_sub13_run_req;
	wire               w_sub13_run_busy;
	wire signed [ 8:0] w_sub13_T_addr;
	reg  signed [ 8:0] r_sub13_T_addr;
	wire        [31:0] w_sub13_T_datain;
	reg         [31:0] r_sub13_T_datain;
	wire        [31:0] w_sub13_T_dataout;
	wire               w_sub13_T_r_w;
	reg                r_sub13_T_r_w;
	wire signed [ 8:0] w_sub13_V_addr;
	reg  signed [ 8:0] r_sub13_V_addr;
	wire        [31:0] w_sub13_V_datain;
	reg         [31:0] r_sub13_V_datain;
	wire        [31:0] w_sub13_V_dataout;
	wire               w_sub13_V_r_w;
	reg                r_sub13_V_r_w;
	wire signed [ 8:0] w_sub13_U_addr;
	reg  signed [ 8:0] r_sub13_U_addr;
	wire        [31:0] w_sub13_U_datain;
	reg         [31:0] r_sub13_U_datain;
	wire        [31:0] w_sub13_U_dataout;
	wire               w_sub13_U_r_w;
	reg                r_sub13_U_r_w;
	wire signed [ 8:0] w_sub13_result_addr;
	reg  signed [ 8:0] r_sub13_result_addr;
	wire        [31:0] w_sub13_result_datain;
	reg         [31:0] r_sub13_result_datain;
	wire        [31:0] w_sub13_result_dataout;
	wire               w_sub13_result_r_w;
	reg                r_sub13_result_r_w;
	reg                r_sub07_run_req;
	wire               w_sub07_run_busy;
	wire signed [ 8:0] w_sub07_T_addr;
	reg  signed [ 8:0] r_sub07_T_addr;
	wire        [31:0] w_sub07_T_datain;
	reg         [31:0] r_sub07_T_datain;
	wire        [31:0] w_sub07_T_dataout;
	wire               w_sub07_T_r_w;
	reg                r_sub07_T_r_w;
	wire signed [ 8:0] w_sub07_V_addr;
	reg  signed [ 8:0] r_sub07_V_addr;
	wire        [31:0] w_sub07_V_datain;
	reg         [31:0] r_sub07_V_datain;
	wire        [31:0] w_sub07_V_dataout;
	wire               w_sub07_V_r_w;
	reg                r_sub07_V_r_w;
	wire signed [ 8:0] w_sub07_U_addr;
	reg  signed [ 8:0] r_sub07_U_addr;
	wire        [31:0] w_sub07_U_datain;
	reg         [31:0] r_sub07_U_datain;
	wire        [31:0] w_sub07_U_dataout;
	wire               w_sub07_U_r_w;
	reg                r_sub07_U_r_w;
	wire signed [ 8:0] w_sub07_result_addr;
	reg  signed [ 8:0] r_sub07_result_addr;
	wire        [31:0] w_sub07_result_datain;
	reg         [31:0] r_sub07_result_datain;
	wire        [31:0] w_sub07_result_dataout;
	wire               w_sub07_result_r_w;
	reg                r_sub07_result_r_w;
	reg                r_sub16_run_req;
	wire               w_sub16_run_busy;
	wire signed [ 8:0] w_sub16_T_addr;
	reg  signed [ 8:0] r_sub16_T_addr;
	wire        [31:0] w_sub16_T_datain;
	reg         [31:0] r_sub16_T_datain;
	wire        [31:0] w_sub16_T_dataout;
	wire               w_sub16_T_r_w;
	reg                r_sub16_T_r_w;
	wire signed [ 8:0] w_sub16_V_addr;
	reg  signed [ 8:0] r_sub16_V_addr;
	wire        [31:0] w_sub16_V_datain;
	reg         [31:0] r_sub16_V_datain;
	wire        [31:0] w_sub16_V_dataout;
	wire               w_sub16_V_r_w;
	reg                r_sub16_V_r_w;
	wire signed [ 8:0] w_sub16_U_addr;
	reg  signed [ 8:0] r_sub16_U_addr;
	wire        [31:0] w_sub16_U_datain;
	reg         [31:0] r_sub16_U_datain;
	wire        [31:0] w_sub16_U_dataout;
	wire               w_sub16_U_r_w;
	reg                r_sub16_U_r_w;
	wire signed [ 8:0] w_sub16_result_addr;
	reg  signed [ 8:0] r_sub16_result_addr;
	wire        [31:0] w_sub16_result_datain;
	reg         [31:0] r_sub16_result_datain;
	wire        [31:0] w_sub16_result_dataout;
	wire               w_sub16_result_r_w;
	reg                r_sub16_result_r_w;
	reg                r_sub06_run_req;
	wire               w_sub06_run_busy;
	wire signed [ 8:0] w_sub06_T_addr;
	reg  signed [ 8:0] r_sub06_T_addr;
	wire        [31:0] w_sub06_T_datain;
	reg         [31:0] r_sub06_T_datain;
	wire        [31:0] w_sub06_T_dataout;
	wire               w_sub06_T_r_w;
	reg                r_sub06_T_r_w;
	wire signed [ 8:0] w_sub06_V_addr;
	reg  signed [ 8:0] r_sub06_V_addr;
	wire        [31:0] w_sub06_V_datain;
	reg         [31:0] r_sub06_V_datain;
	wire        [31:0] w_sub06_V_dataout;
	wire               w_sub06_V_r_w;
	reg                r_sub06_V_r_w;
	wire signed [ 8:0] w_sub06_U_addr;
	reg  signed [ 8:0] r_sub06_U_addr;
	wire        [31:0] w_sub06_U_datain;
	reg         [31:0] r_sub06_U_datain;
	wire        [31:0] w_sub06_U_dataout;
	wire               w_sub06_U_r_w;
	reg                r_sub06_U_r_w;
	wire signed [ 8:0] w_sub06_result_addr;
	reg  signed [ 8:0] r_sub06_result_addr;
	wire        [31:0] w_sub06_result_datain;
	reg         [31:0] r_sub06_result_datain;
	wire        [31:0] w_sub06_result_dataout;
	wire               w_sub06_result_r_w;
	reg                r_sub06_result_r_w;
	reg                r_sub15_run_req;
	wire               w_sub15_run_busy;
	wire signed [ 8:0] w_sub15_T_addr;
	reg  signed [ 8:0] r_sub15_T_addr;
	wire        [31:0] w_sub15_T_datain;
	reg         [31:0] r_sub15_T_datain;
	wire        [31:0] w_sub15_T_dataout;
	wire               w_sub15_T_r_w;
	reg                r_sub15_T_r_w;
	wire signed [ 8:0] w_sub15_V_addr;
	reg  signed [ 8:0] r_sub15_V_addr;
	wire        [31:0] w_sub15_V_datain;
	reg         [31:0] r_sub15_V_datain;
	wire        [31:0] w_sub15_V_dataout;
	wire               w_sub15_V_r_w;
	reg                r_sub15_V_r_w;
	wire signed [ 8:0] w_sub15_U_addr;
	reg  signed [ 8:0] r_sub15_U_addr;
	wire        [31:0] w_sub15_U_datain;
	reg         [31:0] r_sub15_U_datain;
	wire        [31:0] w_sub15_U_dataout;
	wire               w_sub15_U_r_w;
	reg                r_sub15_U_r_w;
	wire signed [ 8:0] w_sub15_result_addr;
	reg  signed [ 8:0] r_sub15_result_addr;
	wire        [31:0] w_sub15_result_datain;
	reg         [31:0] r_sub15_result_datain;
	wire        [31:0] w_sub15_result_dataout;
	wire               w_sub15_result_r_w;
	reg                r_sub15_result_r_w;
	reg                r_sub05_run_req;
	wire               w_sub05_run_busy;
	wire signed [ 8:0] w_sub05_T_addr;
	reg  signed [ 8:0] r_sub05_T_addr;
	wire        [31:0] w_sub05_T_datain;
	reg         [31:0] r_sub05_T_datain;
	wire        [31:0] w_sub05_T_dataout;
	wire               w_sub05_T_r_w;
	reg                r_sub05_T_r_w;
	wire signed [ 8:0] w_sub05_V_addr;
	reg  signed [ 8:0] r_sub05_V_addr;
	wire        [31:0] w_sub05_V_datain;
	reg         [31:0] r_sub05_V_datain;
	wire        [31:0] w_sub05_V_dataout;
	wire               w_sub05_V_r_w;
	reg                r_sub05_V_r_w;
	wire signed [ 8:0] w_sub05_U_addr;
	reg  signed [ 8:0] r_sub05_U_addr;
	wire        [31:0] w_sub05_U_datain;
	reg         [31:0] r_sub05_U_datain;
	wire        [31:0] w_sub05_U_dataout;
	wire               w_sub05_U_r_w;
	reg                r_sub05_U_r_w;
	wire signed [ 8:0] w_sub05_result_addr;
	reg  signed [ 8:0] r_sub05_result_addr;
	wire        [31:0] w_sub05_result_datain;
	reg         [31:0] r_sub05_result_datain;
	wire        [31:0] w_sub05_result_dataout;
	wire               w_sub05_result_r_w;
	reg                r_sub05_result_r_w;
	reg                r_sub18_run_req;
	wire               w_sub18_run_busy;
	wire signed [ 8:0] w_sub18_T_addr;
	reg  signed [ 8:0] r_sub18_T_addr;
	wire        [31:0] w_sub18_T_datain;
	reg         [31:0] r_sub18_T_datain;
	wire        [31:0] w_sub18_T_dataout;
	wire               w_sub18_T_r_w;
	reg                r_sub18_T_r_w;
	wire signed [ 8:0] w_sub18_V_addr;
	reg  signed [ 8:0] r_sub18_V_addr;
	wire        [31:0] w_sub18_V_datain;
	reg         [31:0] r_sub18_V_datain;
	wire        [31:0] w_sub18_V_dataout;
	wire               w_sub18_V_r_w;
	reg                r_sub18_V_r_w;
	wire signed [ 8:0] w_sub18_U_addr;
	reg  signed [ 8:0] r_sub18_U_addr;
	wire        [31:0] w_sub18_U_datain;
	reg         [31:0] r_sub18_U_datain;
	wire        [31:0] w_sub18_U_dataout;
	wire               w_sub18_U_r_w;
	reg                r_sub18_U_r_w;
	wire signed [ 8:0] w_sub18_result_addr;
	reg  signed [ 8:0] r_sub18_result_addr;
	wire        [31:0] w_sub18_result_datain;
	reg         [31:0] r_sub18_result_datain;
	wire        [31:0] w_sub18_result_dataout;
	wire               w_sub18_result_r_w;
	reg                r_sub18_result_r_w;
	reg                r_sub04_run_req;
	wire               w_sub04_run_busy;
	wire signed [ 8:0] w_sub04_T_addr;
	reg  signed [ 8:0] r_sub04_T_addr;
	wire        [31:0] w_sub04_T_datain;
	reg         [31:0] r_sub04_T_datain;
	wire        [31:0] w_sub04_T_dataout;
	wire               w_sub04_T_r_w;
	reg                r_sub04_T_r_w;
	wire signed [ 8:0] w_sub04_V_addr;
	reg  signed [ 8:0] r_sub04_V_addr;
	wire        [31:0] w_sub04_V_datain;
	reg         [31:0] r_sub04_V_datain;
	wire        [31:0] w_sub04_V_dataout;
	wire               w_sub04_V_r_w;
	reg                r_sub04_V_r_w;
	wire signed [ 8:0] w_sub04_U_addr;
	reg  signed [ 8:0] r_sub04_U_addr;
	wire        [31:0] w_sub04_U_datain;
	reg         [31:0] r_sub04_U_datain;
	wire        [31:0] w_sub04_U_dataout;
	wire               w_sub04_U_r_w;
	reg                r_sub04_U_r_w;
	wire signed [ 8:0] w_sub04_result_addr;
	reg  signed [ 8:0] r_sub04_result_addr;
	wire        [31:0] w_sub04_result_datain;
	reg         [31:0] r_sub04_result_datain;
	wire        [31:0] w_sub04_result_dataout;
	wire               w_sub04_result_r_w;
	reg                r_sub04_result_r_w;
	reg                r_sub17_run_req;
	wire               w_sub17_run_busy;
	wire signed [ 8:0] w_sub17_T_addr;
	reg  signed [ 8:0] r_sub17_T_addr;
	wire        [31:0] w_sub17_T_datain;
	reg         [31:0] r_sub17_T_datain;
	wire        [31:0] w_sub17_T_dataout;
	wire               w_sub17_T_r_w;
	reg                r_sub17_T_r_w;
	wire signed [ 8:0] w_sub17_V_addr;
	reg  signed [ 8:0] r_sub17_V_addr;
	wire        [31:0] w_sub17_V_datain;
	reg         [31:0] r_sub17_V_datain;
	wire        [31:0] w_sub17_V_dataout;
	wire               w_sub17_V_r_w;
	reg                r_sub17_V_r_w;
	wire signed [ 8:0] w_sub17_U_addr;
	reg  signed [ 8:0] r_sub17_U_addr;
	wire        [31:0] w_sub17_U_datain;
	reg         [31:0] r_sub17_U_datain;
	wire        [31:0] w_sub17_U_dataout;
	wire               w_sub17_U_r_w;
	reg                r_sub17_U_r_w;
	wire signed [ 8:0] w_sub17_result_addr;
	reg  signed [ 8:0] r_sub17_result_addr;
	wire        [31:0] w_sub17_result_datain;
	reg         [31:0] r_sub17_result_datain;
	wire        [31:0] w_sub17_result_dataout;
	wire               w_sub17_result_r_w;
	reg                r_sub17_result_r_w;
	reg                r_sub10_run_req;
	wire               w_sub10_run_busy;
	wire signed [ 8:0] w_sub10_T_addr;
	reg  signed [ 8:0] r_sub10_T_addr;
	wire        [31:0] w_sub10_T_datain;
	reg         [31:0] r_sub10_T_datain;
	wire        [31:0] w_sub10_T_dataout;
	wire               w_sub10_T_r_w;
	reg                r_sub10_T_r_w;
	wire signed [ 8:0] w_sub10_V_addr;
	reg  signed [ 8:0] r_sub10_V_addr;
	wire        [31:0] w_sub10_V_datain;
	reg         [31:0] r_sub10_V_datain;
	wire        [31:0] w_sub10_V_dataout;
	wire               w_sub10_V_r_w;
	reg                r_sub10_V_r_w;
	wire signed [ 8:0] w_sub10_U_addr;
	reg  signed [ 8:0] r_sub10_U_addr;
	wire        [31:0] w_sub10_U_datain;
	reg         [31:0] r_sub10_U_datain;
	wire        [31:0] w_sub10_U_dataout;
	wire               w_sub10_U_r_w;
	reg                r_sub10_U_r_w;
	wire signed [ 8:0] w_sub10_result_addr;
	reg  signed [ 8:0] r_sub10_result_addr;
	wire        [31:0] w_sub10_result_datain;
	reg         [31:0] r_sub10_result_datain;
	wire        [31:0] w_sub10_result_dataout;
	wire               w_sub10_result_r_w;
	reg                r_sub10_result_r_w;
	reg                r_sub20_run_req;
	wire               w_sub20_run_busy;
	wire signed [ 8:0] w_sub20_T_addr;
	reg  signed [ 8:0] r_sub20_T_addr;
	wire        [31:0] w_sub20_T_datain;
	reg         [31:0] r_sub20_T_datain;
	wire        [31:0] w_sub20_T_dataout;
	wire               w_sub20_T_r_w;
	reg                r_sub20_T_r_w;
	wire signed [ 8:0] w_sub20_V_addr;
	reg  signed [ 8:0] r_sub20_V_addr;
	wire        [31:0] w_sub20_V_datain;
	reg         [31:0] r_sub20_V_datain;
	wire        [31:0] w_sub20_V_dataout;
	wire               w_sub20_V_r_w;
	reg                r_sub20_V_r_w;
	wire signed [ 8:0] w_sub20_U_addr;
	reg  signed [ 8:0] r_sub20_U_addr;
	wire        [31:0] w_sub20_U_datain;
	reg         [31:0] r_sub20_U_datain;
	wire        [31:0] w_sub20_U_dataout;
	wire               w_sub20_U_r_w;
	reg                r_sub20_U_r_w;
	wire signed [ 8:0] w_sub20_result_addr;
	reg  signed [ 8:0] r_sub20_result_addr;
	wire        [31:0] w_sub20_result_datain;
	reg         [31:0] r_sub20_result_datain;
	wire        [31:0] w_sub20_result_dataout;
	wire               w_sub20_result_r_w;
	reg                r_sub20_result_r_w;
	reg                r_sub21_run_req;
	wire               w_sub21_run_busy;
	wire signed [ 8:0] w_sub21_T_addr;
	reg  signed [ 8:0] r_sub21_T_addr;
	wire        [31:0] w_sub21_T_datain;
	reg         [31:0] r_sub21_T_datain;
	wire        [31:0] w_sub21_T_dataout;
	wire               w_sub21_T_r_w;
	reg                r_sub21_T_r_w;
	wire signed [ 8:0] w_sub21_V_addr;
	reg  signed [ 8:0] r_sub21_V_addr;
	wire        [31:0] w_sub21_V_datain;
	reg         [31:0] r_sub21_V_datain;
	wire        [31:0] w_sub21_V_dataout;
	wire               w_sub21_V_r_w;
	reg                r_sub21_V_r_w;
	wire signed [ 8:0] w_sub21_U_addr;
	reg  signed [ 8:0] r_sub21_U_addr;
	wire        [31:0] w_sub21_U_datain;
	reg         [31:0] r_sub21_U_datain;
	wire        [31:0] w_sub21_U_dataout;
	wire               w_sub21_U_r_w;
	reg                r_sub21_U_r_w;
	wire signed [ 8:0] w_sub21_result_addr;
	reg  signed [ 8:0] r_sub21_result_addr;
	wire        [31:0] w_sub21_result_datain;
	reg         [31:0] r_sub21_result_datain;
	wire        [31:0] w_sub21_result_dataout;
	wire               w_sub21_result_r_w;
	reg                r_sub21_result_r_w;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg         [31:0] r_sys_tmp4_float;
	reg         [31:0] r_sys_tmp5_float;
	reg         [31:0] r_sys_tmp6_float;
	reg         [31:0] r_sys_tmp7_float;
	reg         [31:0] r_sys_tmp8_float;
	reg         [31:0] r_sys_tmp9_float;
	reg         [31:0] r_sys_tmp10_float;
	reg         [31:0] r_sys_tmp11_float;
	reg         [31:0] r_sys_tmp12_float;
	reg         [31:0] r_sys_tmp13_float;
	reg         [31:0] r_sys_tmp14_float;
	reg         [31:0] r_sys_tmp15_float;
	reg         [31:0] r_sys_tmp16_float;
	reg         [31:0] r_sys_tmp17_float;
	reg         [31:0] r_sys_tmp18_float;
	reg         [31:0] r_sys_tmp19_float;
	reg         [31:0] r_sys_tmp20_float;
	reg         [31:0] r_sys_tmp21_float;
	reg         [31:0] r_sys_tmp22_float;
	reg         [31:0] r_sys_tmp23_float;
	reg         [31:0] r_sys_tmp24_float;
	reg         [31:0] r_sys_tmp25_float;
	reg         [31:0] r_sys_tmp26_float;
	reg         [31:0] r_sys_tmp27_float;
	reg         [31:0] r_sys_tmp28_float;
	reg         [31:0] r_sys_tmp29_float;
	reg         [31:0] r_sys_tmp30_float;
	reg         [31:0] r_sys_tmp31_float;
	reg         [31:0] r_sys_tmp32_float;
	reg         [31:0] r_sys_tmp33_float;
	reg         [31:0] r_sys_tmp34_float;
	reg         [31:0] r_sys_tmp35_float;
	reg         [31:0] r_sys_tmp36_float;
	reg         [31:0] r_sys_tmp37_float;
	reg         [31:0] r_sys_tmp38_float;
	reg         [31:0] r_sys_tmp39_float;
	reg         [31:0] r_sys_tmp40_float;
	reg         [31:0] r_sys_tmp41_float;
	reg         [31:0] r_sys_tmp42_float;
	reg         [31:0] r_sys_tmp43_float;
	reg         [31:0] r_sys_tmp44_float;
	reg         [31:0] r_sys_tmp45_float;
	reg         [31:0] r_sys_tmp46_float;
	reg         [31:0] r_sys_tmp47_float;
	reg         [31:0] r_sys_tmp48_float;
	reg         [31:0] r_sys_tmp49_float;
	reg         [31:0] r_sys_tmp50_float;
	reg         [31:0] r_sys_tmp51_float;
	reg         [31:0] r_sys_tmp52_float;
	reg         [31:0] r_sys_tmp53_float;
	reg         [31:0] r_sys_tmp54_float;
	reg         [31:0] r_sys_tmp55_float;
	reg         [31:0] r_sys_tmp56_float;
	reg         [31:0] r_sys_tmp57_float;
	reg         [31:0] r_sys_tmp58_float;
	reg         [31:0] r_sys_tmp59_float;
	reg         [31:0] r_sys_tmp60_float;
	reg         [31:0] r_sys_tmp61_float;
	reg         [31:0] r_sys_tmp62_float;
	reg         [31:0] r_sys_tmp63_float;
	reg         [31:0] r_sys_tmp64_float;
	reg         [31:0] r_sys_tmp65_float;
	reg         [31:0] r_sys_tmp66_float;
	reg         [31:0] r_sys_tmp67_float;
	reg         [31:0] r_sys_tmp68_float;
	reg         [31:0] r_sys_tmp69_float;
	reg         [31:0] r_sys_tmp70_float;
	wire signed [31:0] w_sys_tmp1;
	wire signed [31:0] w_sys_tmp3;
	wire        [31:0] w_sys_tmp5;
	wire signed [31:0] w_sys_tmp6;
	wire        [31:0] w_sys_tmp7;
	wire        [31:0] w_sys_tmp8;
	wire        [31:0] w_sys_tmp9;
	wire        [31:0] w_sys_tmp10;
	wire        [31:0] w_sys_tmp11;
	wire        [31:0] w_sys_tmp12;
	wire               w_sys_tmp13;
	wire               w_sys_tmp14;
	wire signed [31:0] w_sys_tmp15;
	wire               w_sys_tmp16;
	wire               w_sys_tmp17;
	wire        [31:0] w_sys_tmp19;
	wire        [31:0] w_sys_tmp20;
	wire signed [31:0] w_sys_tmp21;
	wire signed [31:0] w_sys_tmp23;
	wire signed [31:0] w_sys_tmp24;
	wire signed [31:0] w_sys_tmp25;
	wire        [31:0] w_sys_tmp26;
	wire signed [31:0] w_sys_tmp28;
	wire signed [31:0] w_sys_tmp29;
	wire signed [31:0] w_sys_tmp33;
	wire signed [31:0] w_sys_tmp34;
	wire        [31:0] w_sys_tmp37;
	wire        [31:0] w_sys_tmp38;
	wire        [31:0] w_sys_tmp39;
	wire signed [31:0] w_sys_tmp42;
	wire signed [31:0] w_sys_tmp43;
	wire signed [31:0] w_sys_tmp46;
	wire signed [31:0] w_sys_tmp47;
	wire signed [31:0] w_sys_tmp48;
	wire signed [31:0] w_sys_tmp49;
	wire        [31:0] w_sys_tmp129;
	wire               w_sys_tmp227;
	wire               w_sys_tmp228;
	wire signed [31:0] w_sys_tmp229;
	wire signed [31:0] w_sys_tmp232;
	wire signed [31:0] w_sys_tmp233;
	wire        [31:0] w_sys_tmp234;
	wire signed [31:0] w_sys_tmp238;
	wire signed [31:0] w_sys_tmp239;
	wire signed [31:0] w_sys_tmp244;
	wire signed [31:0] w_sys_tmp245;
	wire signed [31:0] w_sys_tmp250;
	wire signed [31:0] w_sys_tmp251;
	wire signed [31:0] w_sys_tmp256;
	wire signed [31:0] w_sys_tmp257;
	wire signed [31:0] w_sys_tmp262;
	wire signed [31:0] w_sys_tmp263;
	wire signed [31:0] w_sys_tmp280;
	wire signed [31:0] w_sys_tmp281;
	wire signed [31:0] w_sys_tmp286;
	wire signed [31:0] w_sys_tmp287;
	wire signed [31:0] w_sys_tmp292;
	wire signed [31:0] w_sys_tmp293;
	wire signed [31:0] w_sys_tmp298;
	wire signed [31:0] w_sys_tmp299;
	wire signed [31:0] w_sys_tmp316;
	wire signed [31:0] w_sys_tmp317;
	wire signed [31:0] w_sys_tmp322;
	wire signed [31:0] w_sys_tmp323;
	wire signed [31:0] w_sys_tmp328;
	wire signed [31:0] w_sys_tmp329;
	wire signed [31:0] w_sys_tmp334;
	wire signed [31:0] w_sys_tmp335;
	wire signed [31:0] w_sys_tmp352;
	wire signed [31:0] w_sys_tmp353;
	wire signed [31:0] w_sys_tmp358;
	wire signed [31:0] w_sys_tmp359;
	wire signed [31:0] w_sys_tmp364;
	wire signed [31:0] w_sys_tmp365;
	wire signed [31:0] w_sys_tmp376;
	wire signed [31:0] w_sys_tmp377;
	wire signed [31:0] w_sys_tmp382;
	wire signed [31:0] w_sys_tmp383;
	wire signed [31:0] w_sys_tmp388;
	wire signed [31:0] w_sys_tmp389;
	wire        [31:0] w_sys_tmp396;
	wire signed [31:0] w_sys_tmp556;
	wire signed [31:0] w_sys_tmp557;
	wire signed [31:0] w_sys_tmp562;
	wire signed [31:0] w_sys_tmp563;
	wire signed [31:0] w_sys_tmp568;
	wire signed [31:0] w_sys_tmp569;
	wire signed [31:0] w_sys_tmp574;
	wire signed [31:0] w_sys_tmp575;
	wire signed [31:0] w_sys_tmp580;
	wire signed [31:0] w_sys_tmp581;
	wire signed [31:0] w_sys_tmp586;
	wire signed [31:0] w_sys_tmp587;
	wire signed [31:0] w_sys_tmp604;
	wire signed [31:0] w_sys_tmp605;
	wire signed [31:0] w_sys_tmp610;
	wire signed [31:0] w_sys_tmp611;
	wire signed [31:0] w_sys_tmp616;
	wire signed [31:0] w_sys_tmp617;
	wire signed [31:0] w_sys_tmp622;
	wire signed [31:0] w_sys_tmp623;
	wire signed [31:0] w_sys_tmp640;
	wire signed [31:0] w_sys_tmp641;
	wire signed [31:0] w_sys_tmp646;
	wire signed [31:0] w_sys_tmp647;
	wire signed [31:0] w_sys_tmp652;
	wire signed [31:0] w_sys_tmp653;
	wire signed [31:0] w_sys_tmp658;
	wire signed [31:0] w_sys_tmp659;
	wire signed [31:0] w_sys_tmp676;
	wire signed [31:0] w_sys_tmp677;
	wire signed [31:0] w_sys_tmp682;
	wire signed [31:0] w_sys_tmp683;
	wire signed [31:0] w_sys_tmp688;
	wire signed [31:0] w_sys_tmp689;
	wire signed [31:0] w_sys_tmp700;
	wire signed [31:0] w_sys_tmp701;
	wire signed [31:0] w_sys_tmp706;
	wire signed [31:0] w_sys_tmp707;
	wire signed [31:0] w_sys_tmp712;
	wire signed [31:0] w_sys_tmp713;
	wire signed [31:0] w_sys_tmp880;
	wire signed [31:0] w_sys_tmp881;
	wire signed [31:0] w_sys_tmp886;
	wire signed [31:0] w_sys_tmp887;
	wire signed [31:0] w_sys_tmp892;
	wire signed [31:0] w_sys_tmp893;
	wire signed [31:0] w_sys_tmp898;
	wire signed [31:0] w_sys_tmp899;
	wire signed [31:0] w_sys_tmp904;
	wire signed [31:0] w_sys_tmp905;
	wire signed [31:0] w_sys_tmp910;
	wire signed [31:0] w_sys_tmp911;
	wire signed [31:0] w_sys_tmp928;
	wire signed [31:0] w_sys_tmp929;
	wire signed [31:0] w_sys_tmp934;
	wire signed [31:0] w_sys_tmp935;
	wire signed [31:0] w_sys_tmp940;
	wire signed [31:0] w_sys_tmp941;
	wire signed [31:0] w_sys_tmp946;
	wire signed [31:0] w_sys_tmp947;
	wire signed [31:0] w_sys_tmp964;
	wire signed [31:0] w_sys_tmp965;
	wire signed [31:0] w_sys_tmp970;
	wire signed [31:0] w_sys_tmp971;
	wire signed [31:0] w_sys_tmp976;
	wire signed [31:0] w_sys_tmp977;
	wire signed [31:0] w_sys_tmp982;
	wire signed [31:0] w_sys_tmp983;
	wire signed [31:0] w_sys_tmp1000;
	wire signed [31:0] w_sys_tmp1001;
	wire signed [31:0] w_sys_tmp1006;
	wire signed [31:0] w_sys_tmp1007;
	wire signed [31:0] w_sys_tmp1012;
	wire signed [31:0] w_sys_tmp1013;
	wire signed [31:0] w_sys_tmp1024;
	wire signed [31:0] w_sys_tmp1025;
	wire signed [31:0] w_sys_tmp1030;
	wire signed [31:0] w_sys_tmp1031;
	wire signed [31:0] w_sys_tmp1036;
	wire signed [31:0] w_sys_tmp1037;
	wire signed [31:0] w_sys_tmp1204;
	wire signed [31:0] w_sys_tmp1205;
	wire signed [31:0] w_sys_tmp1210;
	wire signed [31:0] w_sys_tmp1211;
	wire signed [31:0] w_sys_tmp1216;
	wire signed [31:0] w_sys_tmp1217;
	wire signed [31:0] w_sys_tmp1222;
	wire signed [31:0] w_sys_tmp1223;
	wire signed [31:0] w_sys_tmp1228;
	wire signed [31:0] w_sys_tmp1229;
	wire signed [31:0] w_sys_tmp1234;
	wire signed [31:0] w_sys_tmp1235;
	wire signed [31:0] w_sys_tmp1252;
	wire signed [31:0] w_sys_tmp1253;
	wire signed [31:0] w_sys_tmp1258;
	wire signed [31:0] w_sys_tmp1259;
	wire signed [31:0] w_sys_tmp1264;
	wire signed [31:0] w_sys_tmp1265;
	wire signed [31:0] w_sys_tmp1270;
	wire signed [31:0] w_sys_tmp1271;
	wire signed [31:0] w_sys_tmp1288;
	wire signed [31:0] w_sys_tmp1289;
	wire signed [31:0] w_sys_tmp1294;
	wire signed [31:0] w_sys_tmp1295;
	wire signed [31:0] w_sys_tmp1300;
	wire signed [31:0] w_sys_tmp1301;
	wire signed [31:0] w_sys_tmp1306;
	wire signed [31:0] w_sys_tmp1307;
	wire signed [31:0] w_sys_tmp1324;
	wire signed [31:0] w_sys_tmp1325;
	wire signed [31:0] w_sys_tmp1330;
	wire signed [31:0] w_sys_tmp1331;
	wire signed [31:0] w_sys_tmp1336;
	wire signed [31:0] w_sys_tmp1337;
	wire signed [31:0] w_sys_tmp1348;
	wire signed [31:0] w_sys_tmp1349;
	wire signed [31:0] w_sys_tmp1354;
	wire signed [31:0] w_sys_tmp1355;
	wire signed [31:0] w_sys_tmp1360;
	wire signed [31:0] w_sys_tmp1361;
	wire signed [31:0] w_sys_tmp1527;
	wire signed [31:0] w_sys_tmp1528;
	wire               w_sys_tmp1529;
	wire               w_sys_tmp1530;
	wire signed [31:0] w_sys_tmp1531;
	wire signed [31:0] w_sys_tmp1534;
	wire signed [31:0] w_sys_tmp1535;
	wire        [31:0] w_sys_tmp1536;
	wire signed [31:0] w_sys_tmp1540;
	wire signed [31:0] w_sys_tmp1541;
	wire signed [31:0] w_sys_tmp1546;
	wire signed [31:0] w_sys_tmp1547;
	wire signed [31:0] w_sys_tmp1552;
	wire signed [31:0] w_sys_tmp1553;
	wire signed [31:0] w_sys_tmp1558;
	wire signed [31:0] w_sys_tmp1559;
	wire signed [31:0] w_sys_tmp1564;
	wire signed [31:0] w_sys_tmp1565;
	wire signed [31:0] w_sys_tmp1582;
	wire signed [31:0] w_sys_tmp1583;
	wire signed [31:0] w_sys_tmp1588;
	wire signed [31:0] w_sys_tmp1589;
	wire signed [31:0] w_sys_tmp1594;
	wire signed [31:0] w_sys_tmp1595;
	wire signed [31:0] w_sys_tmp1600;
	wire signed [31:0] w_sys_tmp1601;
	wire signed [31:0] w_sys_tmp1618;
	wire signed [31:0] w_sys_tmp1619;
	wire signed [31:0] w_sys_tmp1624;
	wire signed [31:0] w_sys_tmp1625;
	wire signed [31:0] w_sys_tmp1630;
	wire signed [31:0] w_sys_tmp1631;
	wire signed [31:0] w_sys_tmp1636;
	wire signed [31:0] w_sys_tmp1637;
	wire signed [31:0] w_sys_tmp1654;
	wire signed [31:0] w_sys_tmp1655;
	wire signed [31:0] w_sys_tmp1660;
	wire signed [31:0] w_sys_tmp1661;
	wire signed [31:0] w_sys_tmp1666;
	wire signed [31:0] w_sys_tmp1667;
	wire signed [31:0] w_sys_tmp1678;
	wire signed [31:0] w_sys_tmp1679;
	wire signed [31:0] w_sys_tmp1684;
	wire signed [31:0] w_sys_tmp1685;
	wire signed [31:0] w_sys_tmp1690;
	wire signed [31:0] w_sys_tmp1691;
	wire        [31:0] w_sys_tmp1698;
	wire signed [31:0] w_sys_tmp1857;
	wire               w_sys_tmp1858;
	wire               w_sys_tmp1859;
	wire signed [31:0] w_sys_tmp1860;
	wire               w_sys_tmp1861;
	wire               w_sys_tmp1862;
	wire signed [31:0] w_sys_tmp1865;
	wire signed [31:0] w_sys_tmp1866;
	wire        [31:0] w_sys_tmp1867;
	wire signed [31:0] w_sys_tmp1869;
	wire signed [31:0] w_sys_tmp1870;
	wire        [31:0] w_sys_tmp1872;
	wire signed [31:0] w_sys_tmp1873;
	wire signed [31:0] w_sys_tmp1874;
	wire signed [31:0] w_sys_tmp1875;
	wire signed [31:0] w_sys_tmp1877;
	wire               w_sys_tmp1878;
	wire               w_sys_tmp1879;
	wire signed [31:0] w_sys_tmp1882;
	wire signed [31:0] w_sys_tmp1883;
	wire signed [31:0] w_sys_tmp1884;
	wire        [31:0] w_sys_tmp1885;
	wire signed [31:0] w_sys_tmp1887;
	wire signed [31:0] w_sys_tmp1888;
	wire signed [31:0] w_sys_tmp1891;
	wire signed [31:0] w_sys_tmp1892;
	wire signed [31:0] w_sys_tmp1965;
	wire signed [31:0] w_sys_tmp1966;
	wire               w_sys_tmp1967;
	wire               w_sys_tmp1968;
	wire signed [31:0] w_sys_tmp1969;
	wire signed [31:0] w_sys_tmp1970;
	wire signed [31:0] w_sys_tmp1973;
	wire signed [31:0] w_sys_tmp1974;
	wire signed [31:0] w_sys_tmp1975;
	wire        [31:0] w_sys_tmp1976;
	wire signed [31:0] w_sys_tmp1977;
	wire               w_sys_tmp2014;
	wire               w_sys_tmp2015;
	wire signed [31:0] w_sys_tmp2016;
	wire signed [31:0] w_sys_tmp2019;
	wire signed [31:0] w_sys_tmp2020;
	wire        [31:0] w_sys_tmp2021;
	wire signed [31:0] w_sys_tmp2025;
	wire signed [31:0] w_sys_tmp2026;
	wire signed [31:0] w_sys_tmp2031;
	wire signed [31:0] w_sys_tmp2032;
	wire signed [31:0] w_sys_tmp2037;
	wire signed [31:0] w_sys_tmp2038;
	wire signed [31:0] w_sys_tmp2043;
	wire signed [31:0] w_sys_tmp2044;
	wire signed [31:0] w_sys_tmp2049;
	wire signed [31:0] w_sys_tmp2050;
	wire signed [31:0] w_sys_tmp2067;
	wire signed [31:0] w_sys_tmp2068;
	wire signed [31:0] w_sys_tmp2073;
	wire signed [31:0] w_sys_tmp2074;
	wire signed [31:0] w_sys_tmp2079;
	wire signed [31:0] w_sys_tmp2080;
	wire signed [31:0] w_sys_tmp2085;
	wire signed [31:0] w_sys_tmp2086;
	wire signed [31:0] w_sys_tmp2103;
	wire signed [31:0] w_sys_tmp2104;
	wire signed [31:0] w_sys_tmp2109;
	wire signed [31:0] w_sys_tmp2110;
	wire signed [31:0] w_sys_tmp2115;
	wire signed [31:0] w_sys_tmp2116;
	wire signed [31:0] w_sys_tmp2121;
	wire signed [31:0] w_sys_tmp2122;
	wire signed [31:0] w_sys_tmp2139;
	wire signed [31:0] w_sys_tmp2140;
	wire signed [31:0] w_sys_tmp2145;
	wire signed [31:0] w_sys_tmp2146;
	wire signed [31:0] w_sys_tmp2151;
	wire signed [31:0] w_sys_tmp2152;
	wire signed [31:0] w_sys_tmp2163;
	wire signed [31:0] w_sys_tmp2164;
	wire signed [31:0] w_sys_tmp2169;
	wire signed [31:0] w_sys_tmp2170;
	wire signed [31:0] w_sys_tmp2175;
	wire signed [31:0] w_sys_tmp2176;
	wire signed [31:0] w_sys_tmp2181;
	wire signed [31:0] w_sys_tmp2182;
	wire signed [31:0] w_sys_tmp2187;
	wire signed [31:0] w_sys_tmp2188;
	wire signed [31:0] w_sys_tmp2193;
	wire signed [31:0] w_sys_tmp2194;
	wire signed [31:0] w_sys_tmp2199;
	wire signed [31:0] w_sys_tmp2200;
	wire signed [31:0] w_sys_tmp2205;
	wire signed [31:0] w_sys_tmp2206;
	wire signed [31:0] w_sys_tmp2211;
	wire signed [31:0] w_sys_tmp2212;
	wire signed [31:0] w_sys_tmp2229;
	wire signed [31:0] w_sys_tmp2230;
	wire signed [31:0] w_sys_tmp2235;
	wire signed [31:0] w_sys_tmp2236;
	wire signed [31:0] w_sys_tmp2241;
	wire signed [31:0] w_sys_tmp2242;
	wire signed [31:0] w_sys_tmp2247;
	wire signed [31:0] w_sys_tmp2248;
	wire signed [31:0] w_sys_tmp2265;
	wire signed [31:0] w_sys_tmp2266;
	wire signed [31:0] w_sys_tmp2271;
	wire signed [31:0] w_sys_tmp2272;
	wire signed [31:0] w_sys_tmp2277;
	wire signed [31:0] w_sys_tmp2278;
	wire signed [31:0] w_sys_tmp2283;
	wire signed [31:0] w_sys_tmp2284;
	wire signed [31:0] w_sys_tmp2301;
	wire signed [31:0] w_sys_tmp2302;
	wire signed [31:0] w_sys_tmp2307;
	wire signed [31:0] w_sys_tmp2308;
	wire signed [31:0] w_sys_tmp2313;
	wire signed [31:0] w_sys_tmp2314;
	wire signed [31:0] w_sys_tmp2325;
	wire signed [31:0] w_sys_tmp2326;
	wire signed [31:0] w_sys_tmp2331;
	wire signed [31:0] w_sys_tmp2332;
	wire signed [31:0] w_sys_tmp2337;
	wire signed [31:0] w_sys_tmp2338;
	wire signed [31:0] w_sys_tmp2343;
	wire signed [31:0] w_sys_tmp2344;
	wire signed [31:0] w_sys_tmp2349;
	wire signed [31:0] w_sys_tmp2350;
	wire signed [31:0] w_sys_tmp2355;
	wire signed [31:0] w_sys_tmp2356;
	wire signed [31:0] w_sys_tmp2361;
	wire signed [31:0] w_sys_tmp2362;
	wire signed [31:0] w_sys_tmp2367;
	wire signed [31:0] w_sys_tmp2368;
	wire signed [31:0] w_sys_tmp2373;
	wire signed [31:0] w_sys_tmp2374;
	wire signed [31:0] w_sys_tmp2391;
	wire signed [31:0] w_sys_tmp2392;
	wire signed [31:0] w_sys_tmp2397;
	wire signed [31:0] w_sys_tmp2398;
	wire signed [31:0] w_sys_tmp2403;
	wire signed [31:0] w_sys_tmp2404;
	wire signed [31:0] w_sys_tmp2409;
	wire signed [31:0] w_sys_tmp2410;
	wire signed [31:0] w_sys_tmp2427;
	wire signed [31:0] w_sys_tmp2428;
	wire signed [31:0] w_sys_tmp2433;
	wire signed [31:0] w_sys_tmp2434;
	wire signed [31:0] w_sys_tmp2439;
	wire signed [31:0] w_sys_tmp2440;
	wire signed [31:0] w_sys_tmp2445;
	wire signed [31:0] w_sys_tmp2446;
	wire signed [31:0] w_sys_tmp2463;
	wire signed [31:0] w_sys_tmp2464;
	wire signed [31:0] w_sys_tmp2469;
	wire signed [31:0] w_sys_tmp2470;
	wire signed [31:0] w_sys_tmp2475;
	wire signed [31:0] w_sys_tmp2476;
	wire signed [31:0] w_sys_tmp2487;
	wire signed [31:0] w_sys_tmp2488;
	wire signed [31:0] w_sys_tmp2493;
	wire signed [31:0] w_sys_tmp2494;
	wire signed [31:0] w_sys_tmp2499;
	wire signed [31:0] w_sys_tmp2500;
	wire signed [31:0] w_sys_tmp2505;
	wire signed [31:0] w_sys_tmp2506;
	wire signed [31:0] w_sys_tmp2511;
	wire signed [31:0] w_sys_tmp2512;
	wire signed [31:0] w_sys_tmp2517;
	wire signed [31:0] w_sys_tmp2518;
	wire signed [31:0] w_sys_tmp2523;
	wire signed [31:0] w_sys_tmp2524;
	wire signed [31:0] w_sys_tmp2529;
	wire signed [31:0] w_sys_tmp2530;
	wire signed [31:0] w_sys_tmp2535;
	wire signed [31:0] w_sys_tmp2536;
	wire signed [31:0] w_sys_tmp2553;
	wire signed [31:0] w_sys_tmp2554;
	wire signed [31:0] w_sys_tmp2559;
	wire signed [31:0] w_sys_tmp2560;
	wire signed [31:0] w_sys_tmp2565;
	wire signed [31:0] w_sys_tmp2566;
	wire signed [31:0] w_sys_tmp2571;
	wire signed [31:0] w_sys_tmp2572;
	wire signed [31:0] w_sys_tmp2589;
	wire signed [31:0] w_sys_tmp2590;
	wire signed [31:0] w_sys_tmp2595;
	wire signed [31:0] w_sys_tmp2596;
	wire signed [31:0] w_sys_tmp2601;
	wire signed [31:0] w_sys_tmp2602;
	wire signed [31:0] w_sys_tmp2607;
	wire signed [31:0] w_sys_tmp2608;
	wire signed [31:0] w_sys_tmp2625;
	wire signed [31:0] w_sys_tmp2626;
	wire signed [31:0] w_sys_tmp2631;
	wire signed [31:0] w_sys_tmp2632;
	wire signed [31:0] w_sys_tmp2637;
	wire signed [31:0] w_sys_tmp2638;
	wire signed [31:0] w_sys_tmp2649;
	wire signed [31:0] w_sys_tmp2650;
	wire signed [31:0] w_sys_tmp2655;
	wire signed [31:0] w_sys_tmp2656;
	wire signed [31:0] w_sys_tmp2661;
	wire signed [31:0] w_sys_tmp2662;
	wire signed [31:0] w_sys_tmp2666;
	wire signed [31:0] w_sys_tmp2667;
	wire               w_sys_tmp2668;
	wire               w_sys_tmp2669;
	wire signed [31:0] w_sys_tmp2670;
	wire signed [31:0] w_sys_tmp2673;
	wire signed [31:0] w_sys_tmp2674;
	wire        [31:0] w_sys_tmp2675;
	wire signed [31:0] w_sys_tmp2679;
	wire signed [31:0] w_sys_tmp2680;
	wire signed [31:0] w_sys_tmp2685;
	wire signed [31:0] w_sys_tmp2686;
	wire signed [31:0] w_sys_tmp2691;
	wire signed [31:0] w_sys_tmp2692;
	wire signed [31:0] w_sys_tmp2697;
	wire signed [31:0] w_sys_tmp2698;
	wire signed [31:0] w_sys_tmp2703;
	wire signed [31:0] w_sys_tmp2704;
	wire signed [31:0] w_sys_tmp2721;
	wire signed [31:0] w_sys_tmp2722;
	wire signed [31:0] w_sys_tmp2727;
	wire signed [31:0] w_sys_tmp2728;
	wire signed [31:0] w_sys_tmp2733;
	wire signed [31:0] w_sys_tmp2734;
	wire signed [31:0] w_sys_tmp2739;
	wire signed [31:0] w_sys_tmp2740;
	wire signed [31:0] w_sys_tmp2757;
	wire signed [31:0] w_sys_tmp2758;
	wire signed [31:0] w_sys_tmp2763;
	wire signed [31:0] w_sys_tmp2764;
	wire signed [31:0] w_sys_tmp2769;
	wire signed [31:0] w_sys_tmp2770;
	wire signed [31:0] w_sys_tmp2775;
	wire signed [31:0] w_sys_tmp2776;
	wire signed [31:0] w_sys_tmp2793;
	wire signed [31:0] w_sys_tmp2794;
	wire signed [31:0] w_sys_tmp2799;
	wire signed [31:0] w_sys_tmp2800;
	wire signed [31:0] w_sys_tmp2805;
	wire signed [31:0] w_sys_tmp2806;
	wire signed [31:0] w_sys_tmp2817;
	wire signed [31:0] w_sys_tmp2818;
	wire signed [31:0] w_sys_tmp2823;
	wire signed [31:0] w_sys_tmp2824;
	wire signed [31:0] w_sys_tmp2829;
	wire signed [31:0] w_sys_tmp2830;
	wire signed [31:0] w_sys_tmp2834;
	wire signed [31:0] w_sys_tmp2835;
	wire               w_sys_tmp2836;
	wire               w_sys_tmp2837;
	wire signed [31:0] w_sys_tmp2838;
	wire signed [31:0] w_sys_tmp2841;
	wire signed [31:0] w_sys_tmp2842;
	wire        [31:0] w_sys_tmp2843;
	wire signed [31:0] w_sys_tmp2847;
	wire signed [31:0] w_sys_tmp2848;
	wire signed [31:0] w_sys_tmp2853;
	wire signed [31:0] w_sys_tmp2854;
	wire signed [31:0] w_sys_tmp2859;
	wire signed [31:0] w_sys_tmp2860;
	wire signed [31:0] w_sys_tmp2865;
	wire signed [31:0] w_sys_tmp2866;
	wire signed [31:0] w_sys_tmp2870;
	wire signed [31:0] w_sys_tmp2871;
	wire signed [31:0] w_sys_tmp2875;
	wire signed [31:0] w_sys_tmp2876;
	wire signed [31:0] w_sys_tmp2880;
	wire signed [31:0] w_sys_tmp2881;
	wire signed [31:0] w_sys_tmp2885;
	wire signed [31:0] w_sys_tmp2886;
	wire signed [31:0] w_sys_tmp2890;
	wire signed [31:0] w_sys_tmp2891;
	wire signed [31:0] w_sys_tmp2895;
	wire signed [31:0] w_sys_tmp2896;
	wire signed [31:0] w_sys_tmp2900;
	wire signed [31:0] w_sys_tmp2901;
	wire signed [31:0] w_sys_tmp2905;
	wire signed [31:0] w_sys_tmp2906;
	wire signed [31:0] w_sys_tmp2910;
	wire signed [31:0] w_sys_tmp2911;
	wire signed [31:0] w_sys_tmp2915;
	wire signed [31:0] w_sys_tmp2916;
	wire signed [31:0] w_sys_tmp2920;
	wire signed [31:0] w_sys_tmp2921;
	wire signed [31:0] w_sys_tmp2925;
	wire signed [31:0] w_sys_tmp2926;
	wire signed [31:0] w_sys_tmp2930;
	wire signed [31:0] w_sys_tmp2931;
	wire signed [31:0] w_sys_tmp2935;
	wire signed [31:0] w_sys_tmp2936;
	wire signed [31:0] w_sys_tmp2940;
	wire signed [31:0] w_sys_tmp2941;
	wire signed [31:0] w_sys_tmp2945;
	wire signed [31:0] w_sys_tmp2946;
	wire signed [31:0] w_sys_tmp2950;
	wire signed [31:0] w_sys_tmp2951;
	wire signed [31:0] w_sys_tmp2955;
	wire signed [31:0] w_sys_tmp2956;
	wire signed [31:0] w_sys_tmp2960;
	wire signed [31:0] w_sys_tmp2961;
	wire signed [31:0] w_sys_tmp2965;
	wire signed [31:0] w_sys_tmp2966;
	wire signed [31:0] w_sys_tmp2970;
	wire signed [31:0] w_sys_tmp2971;
	wire signed [31:0] w_sys_tmp2975;
	wire signed [31:0] w_sys_tmp2976;
	wire signed [31:0] w_sys_tmp2980;
	wire signed [31:0] w_sys_tmp2981;
	wire signed [31:0] w_sys_tmp2985;
	wire signed [31:0] w_sys_tmp2986;
	wire signed [31:0] w_sys_tmp2990;
	wire signed [31:0] w_sys_tmp2991;
	wire signed [31:0] w_sys_tmp2995;
	wire signed [31:0] w_sys_tmp2996;
	wire signed [31:0] w_sys_tmp3000;
	wire signed [31:0] w_sys_tmp3001;
	wire signed [31:0] w_sys_tmp3005;
	wire signed [31:0] w_sys_tmp3006;
	wire signed [31:0] w_sys_tmp3010;
	wire signed [31:0] w_sys_tmp3011;
	wire signed [31:0] w_sys_tmp3015;
	wire signed [31:0] w_sys_tmp3016;
	wire signed [31:0] w_sys_tmp3020;
	wire signed [31:0] w_sys_tmp3021;
	wire signed [31:0] w_sys_tmp3025;
	wire signed [31:0] w_sys_tmp3026;
	wire signed [31:0] w_sys_tmp3030;
	wire signed [31:0] w_sys_tmp3031;
	wire signed [31:0] w_sys_tmp3035;
	wire signed [31:0] w_sys_tmp3036;
	wire signed [31:0] w_sys_tmp3040;
	wire signed [31:0] w_sys_tmp3041;
	wire signed [31:0] w_sys_tmp3045;
	wire signed [31:0] w_sys_tmp3046;
	wire signed [31:0] w_sys_tmp3050;
	wire signed [31:0] w_sys_tmp3051;
	wire signed [31:0] w_sys_tmp3055;
	wire signed [31:0] w_sys_tmp3056;
	wire signed [31:0] w_sys_tmp3060;
	wire signed [31:0] w_sys_tmp3061;
	wire signed [31:0] w_sys_tmp3065;
	wire signed [31:0] w_sys_tmp3066;
	wire signed [31:0] w_sys_tmp3070;
	wire signed [31:0] w_sys_tmp3071;
	wire signed [31:0] w_sys_tmp3075;
	wire signed [31:0] w_sys_tmp3076;
	wire signed [31:0] w_sys_tmp3080;
	wire signed [31:0] w_sys_tmp3081;
	wire signed [31:0] w_sys_tmp3085;
	wire signed [31:0] w_sys_tmp3086;
	wire signed [31:0] w_sys_tmp3090;
	wire signed [31:0] w_sys_tmp3091;
	wire signed [31:0] w_sys_tmp3095;
	wire signed [31:0] w_sys_tmp3096;
	wire signed [31:0] w_sys_tmp3100;
	wire signed [31:0] w_sys_tmp3101;
	wire signed [31:0] w_sys_tmp3105;
	wire signed [31:0] w_sys_tmp3106;
	wire signed [31:0] w_sys_tmp3110;
	wire signed [31:0] w_sys_tmp3111;
	wire signed [31:0] w_sys_tmp3115;
	wire signed [31:0] w_sys_tmp3116;
	wire signed [31:0] w_sys_tmp3120;
	wire signed [31:0] w_sys_tmp3121;
	wire signed [31:0] w_sys_tmp3125;
	wire signed [31:0] w_sys_tmp3126;
	wire signed [31:0] w_sys_tmp3130;
	wire signed [31:0] w_sys_tmp3131;
	wire signed [31:0] w_sys_tmp3135;
	wire signed [31:0] w_sys_tmp3136;
	wire signed [31:0] w_sys_tmp3140;
	wire signed [31:0] w_sys_tmp3141;
	wire signed [31:0] w_sys_tmp3145;
	wire signed [31:0] w_sys_tmp3146;
	wire signed [31:0] w_sys_tmp3150;
	wire signed [31:0] w_sys_tmp3151;
	wire signed [31:0] w_sys_tmp3155;
	wire signed [31:0] w_sys_tmp3156;
	wire signed [31:0] w_sys_tmp3160;
	wire signed [31:0] w_sys_tmp3161;
	wire signed [31:0] w_sys_tmp3165;
	wire signed [31:0] w_sys_tmp3166;
	wire signed [31:0] w_sys_tmp3170;
	wire signed [31:0] w_sys_tmp3171;
	wire signed [31:0] w_sys_tmp3175;
	wire signed [31:0] w_sys_tmp3176;
	wire signed [31:0] w_sys_tmp3180;
	wire signed [31:0] w_sys_tmp3181;
	wire signed [31:0] w_sys_tmp3185;
	wire signed [31:0] w_sys_tmp3186;
	wire signed [31:0] w_sys_tmp3190;
	wire signed [31:0] w_sys_tmp3191;
	wire signed [31:0] w_sys_tmp3195;
	wire signed [31:0] w_sys_tmp3196;
	wire signed [31:0] w_sys_tmp3200;
	wire signed [31:0] w_sys_tmp3201;
	wire signed [31:0] w_sys_tmp3205;
	wire signed [31:0] w_sys_tmp3206;
	wire signed [31:0] w_sys_tmp3210;
	wire signed [31:0] w_sys_tmp3211;
	wire signed [31:0] w_sys_tmp3215;
	wire signed [31:0] w_sys_tmp3216;
	wire signed [31:0] w_sys_tmp3220;
	wire signed [31:0] w_sys_tmp3221;
	wire signed [31:0] w_sys_tmp3224;
	wire signed [31:0] w_sys_tmp3225;
	wire               w_sys_tmp3226;
	wire               w_sys_tmp3227;
	wire signed [31:0] w_sys_tmp3228;
	wire signed [31:0] w_sys_tmp3231;
	wire signed [31:0] w_sys_tmp3232;
	wire        [31:0] w_sys_tmp3233;
	wire signed [31:0] w_sys_tmp3237;
	wire signed [31:0] w_sys_tmp3238;
	wire signed [31:0] w_sys_tmp3243;
	wire signed [31:0] w_sys_tmp3244;
	wire signed [31:0] w_sys_tmp3249;
	wire signed [31:0] w_sys_tmp3250;
	wire signed [31:0] w_sys_tmp3255;
	wire signed [31:0] w_sys_tmp3256;
	wire signed [31:0] w_sys_tmp3260;
	wire signed [31:0] w_sys_tmp3261;
	wire signed [31:0] w_sys_tmp3265;
	wire signed [31:0] w_sys_tmp3266;
	wire signed [31:0] w_sys_tmp3270;
	wire signed [31:0] w_sys_tmp3271;
	wire signed [31:0] w_sys_tmp3275;
	wire signed [31:0] w_sys_tmp3276;
	wire signed [31:0] w_sys_tmp3280;
	wire signed [31:0] w_sys_tmp3281;
	wire signed [31:0] w_sys_tmp3285;
	wire signed [31:0] w_sys_tmp3286;
	wire signed [31:0] w_sys_tmp3290;
	wire signed [31:0] w_sys_tmp3291;
	wire signed [31:0] w_sys_tmp3295;
	wire signed [31:0] w_sys_tmp3296;
	wire signed [31:0] w_sys_tmp3300;
	wire signed [31:0] w_sys_tmp3301;
	wire signed [31:0] w_sys_tmp3305;
	wire signed [31:0] w_sys_tmp3306;
	wire signed [31:0] w_sys_tmp3310;
	wire signed [31:0] w_sys_tmp3311;
	wire signed [31:0] w_sys_tmp3315;
	wire signed [31:0] w_sys_tmp3316;
	wire signed [31:0] w_sys_tmp3320;
	wire signed [31:0] w_sys_tmp3321;
	wire signed [31:0] w_sys_tmp3325;
	wire signed [31:0] w_sys_tmp3326;
	wire signed [31:0] w_sys_tmp3329;
	wire        [31:0] w_sys_tmp3330;
	wire signed [31:0] w_sys_tmp3331;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign o_run_return = r_sys_run_return;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 5'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 7'h1);
	assign w_fld_T_0_addr_0 = 9'sh0;
	assign w_fld_T_0_datain_0 = 32'h0;
	assign w_fld_T_0_r_w_0 = 1'h0;
	assign w_fld_T_0_ce_0 = w_sys_ce;
	assign w_fld_T_0_ce_1 = w_sys_ce;
	assign w_fld_TT_1_addr_0 = 9'sh0;
	assign w_fld_TT_1_datain_0 = 32'h0;
	assign w_fld_TT_1_r_w_0 = 1'h0;
	assign w_fld_TT_1_ce_0 = w_sys_ce;
	assign w_fld_TT_1_ce_1 = w_sys_ce;
	assign w_fld_U_2_addr_0 = 9'sh0;
	assign w_fld_U_2_datain_0 = 32'h0;
	assign w_fld_U_2_r_w_0 = 1'h0;
	assign w_fld_U_2_ce_0 = w_sys_ce;
	assign w_fld_U_2_ce_1 = w_sys_ce;
	assign w_fld_V_3_addr_0 = 9'sh0;
	assign w_fld_V_3_datain_0 = 32'h0;
	assign w_fld_V_3_r_w_0 = 1'h0;
	assign w_fld_V_3_ce_0 = w_sys_ce;
	assign w_fld_V_3_ce_1 = w_sys_ce;
	assign w_sub19_T_addr = ( (|r_sys_processing_methodID) ? r_sub19_T_addr : 9'sh0 ) ;
	assign w_sub19_T_datain = ( (|r_sys_processing_methodID) ? r_sub19_T_datain : 32'h0 ) ;
	assign w_sub19_T_r_w = ( (|r_sys_processing_methodID) ? r_sub19_T_r_w : 1'h0 ) ;
	assign w_sub19_V_addr = ( (|r_sys_processing_methodID) ? r_sub19_V_addr : 9'sh0 ) ;
	assign w_sub19_V_datain = ( (|r_sys_processing_methodID) ? r_sub19_V_datain : 32'h0 ) ;
	assign w_sub19_V_r_w = ( (|r_sys_processing_methodID) ? r_sub19_V_r_w : 1'h0 ) ;
	assign w_sub19_U_addr = ( (|r_sys_processing_methodID) ? r_sub19_U_addr : 9'sh0 ) ;
	assign w_sub19_U_datain = ( (|r_sys_processing_methodID) ? r_sub19_U_datain : 32'h0 ) ;
	assign w_sub19_U_r_w = ( (|r_sys_processing_methodID) ? r_sub19_U_r_w : 1'h0 ) ;
	assign w_sub19_result_addr = ( (|r_sys_processing_methodID) ? r_sub19_result_addr : 9'sh0 ) ;
	assign w_sub19_result_datain = ( (|r_sys_processing_methodID) ? r_sub19_result_datain : 32'h0 ) ;
	assign w_sub19_result_r_w = ( (|r_sys_processing_methodID) ? r_sub19_result_r_w : 1'h0 ) ;
	assign w_sub09_T_addr = ( (|r_sys_processing_methodID) ? r_sub09_T_addr : 9'sh0 ) ;
	assign w_sub09_T_datain = ( (|r_sys_processing_methodID) ? r_sub09_T_datain : 32'h0 ) ;
	assign w_sub09_T_r_w = ( (|r_sys_processing_methodID) ? r_sub09_T_r_w : 1'h0 ) ;
	assign w_sub09_V_addr = ( (|r_sys_processing_methodID) ? r_sub09_V_addr : 9'sh0 ) ;
	assign w_sub09_V_datain = ( (|r_sys_processing_methodID) ? r_sub09_V_datain : 32'h0 ) ;
	assign w_sub09_V_r_w = ( (|r_sys_processing_methodID) ? r_sub09_V_r_w : 1'h0 ) ;
	assign w_sub09_U_addr = ( (|r_sys_processing_methodID) ? r_sub09_U_addr : 9'sh0 ) ;
	assign w_sub09_U_datain = ( (|r_sys_processing_methodID) ? r_sub09_U_datain : 32'h0 ) ;
	assign w_sub09_U_r_w = ( (|r_sys_processing_methodID) ? r_sub09_U_r_w : 1'h0 ) ;
	assign w_sub09_result_addr = ( (|r_sys_processing_methodID) ? r_sub09_result_addr : 9'sh0 ) ;
	assign w_sub09_result_datain = ( (|r_sys_processing_methodID) ? r_sub09_result_datain : 32'h0 ) ;
	assign w_sub09_result_r_w = ( (|r_sys_processing_methodID) ? r_sub09_result_r_w : 1'h0 ) ;
	assign w_sub08_T_addr = ( (|r_sys_processing_methodID) ? r_sub08_T_addr : 9'sh0 ) ;
	assign w_sub08_T_datain = ( (|r_sys_processing_methodID) ? r_sub08_T_datain : 32'h0 ) ;
	assign w_sub08_T_r_w = ( (|r_sys_processing_methodID) ? r_sub08_T_r_w : 1'h0 ) ;
	assign w_sub08_V_addr = ( (|r_sys_processing_methodID) ? r_sub08_V_addr : 9'sh0 ) ;
	assign w_sub08_V_datain = ( (|r_sys_processing_methodID) ? r_sub08_V_datain : 32'h0 ) ;
	assign w_sub08_V_r_w = ( (|r_sys_processing_methodID) ? r_sub08_V_r_w : 1'h0 ) ;
	assign w_sub08_U_addr = ( (|r_sys_processing_methodID) ? r_sub08_U_addr : 9'sh0 ) ;
	assign w_sub08_U_datain = ( (|r_sys_processing_methodID) ? r_sub08_U_datain : 32'h0 ) ;
	assign w_sub08_U_r_w = ( (|r_sys_processing_methodID) ? r_sub08_U_r_w : 1'h0 ) ;
	assign w_sub08_result_addr = ( (|r_sys_processing_methodID) ? r_sub08_result_addr : 9'sh0 ) ;
	assign w_sub08_result_datain = ( (|r_sys_processing_methodID) ? r_sub08_result_datain : 32'h0 ) ;
	assign w_sub08_result_r_w = ( (|r_sys_processing_methodID) ? r_sub08_result_r_w : 1'h0 ) ;
	assign w_sub24_T_addr = ( (|r_sys_processing_methodID) ? r_sub24_T_addr : 9'sh0 ) ;
	assign w_sub24_T_datain = ( (|r_sys_processing_methodID) ? r_sub24_T_datain : 32'h0 ) ;
	assign w_sub24_T_r_w = ( (|r_sys_processing_methodID) ? r_sub24_T_r_w : 1'h0 ) ;
	assign w_sub24_V_addr = ( (|r_sys_processing_methodID) ? r_sub24_V_addr : 9'sh0 ) ;
	assign w_sub24_V_datain = ( (|r_sys_processing_methodID) ? r_sub24_V_datain : 32'h0 ) ;
	assign w_sub24_V_r_w = ( (|r_sys_processing_methodID) ? r_sub24_V_r_w : 1'h0 ) ;
	assign w_sub24_U_addr = ( (|r_sys_processing_methodID) ? r_sub24_U_addr : 9'sh0 ) ;
	assign w_sub24_U_datain = ( (|r_sys_processing_methodID) ? r_sub24_U_datain : 32'h0 ) ;
	assign w_sub24_U_r_w = ( (|r_sys_processing_methodID) ? r_sub24_U_r_w : 1'h0 ) ;
	assign w_sub24_result_addr = ( (|r_sys_processing_methodID) ? r_sub24_result_addr : 9'sh0 ) ;
	assign w_sub24_result_datain = ( (|r_sys_processing_methodID) ? r_sub24_result_datain : 32'h0 ) ;
	assign w_sub24_result_r_w = ( (|r_sys_processing_methodID) ? r_sub24_result_r_w : 1'h0 ) ;
	assign w_sub22_T_addr = ( (|r_sys_processing_methodID) ? r_sub22_T_addr : 9'sh0 ) ;
	assign w_sub22_T_datain = ( (|r_sys_processing_methodID) ? r_sub22_T_datain : 32'h0 ) ;
	assign w_sub22_T_r_w = ( (|r_sys_processing_methodID) ? r_sub22_T_r_w : 1'h0 ) ;
	assign w_sub22_V_addr = ( (|r_sys_processing_methodID) ? r_sub22_V_addr : 9'sh0 ) ;
	assign w_sub22_V_datain = ( (|r_sys_processing_methodID) ? r_sub22_V_datain : 32'h0 ) ;
	assign w_sub22_V_r_w = ( (|r_sys_processing_methodID) ? r_sub22_V_r_w : 1'h0 ) ;
	assign w_sub22_U_addr = ( (|r_sys_processing_methodID) ? r_sub22_U_addr : 9'sh0 ) ;
	assign w_sub22_U_datain = ( (|r_sys_processing_methodID) ? r_sub22_U_datain : 32'h0 ) ;
	assign w_sub22_U_r_w = ( (|r_sys_processing_methodID) ? r_sub22_U_r_w : 1'h0 ) ;
	assign w_sub22_result_addr = ( (|r_sys_processing_methodID) ? r_sub22_result_addr : 9'sh0 ) ;
	assign w_sub22_result_datain = ( (|r_sys_processing_methodID) ? r_sub22_result_datain : 32'h0 ) ;
	assign w_sub22_result_r_w = ( (|r_sys_processing_methodID) ? r_sub22_result_r_w : 1'h0 ) ;
	assign w_sub23_T_addr = ( (|r_sys_processing_methodID) ? r_sub23_T_addr : 9'sh0 ) ;
	assign w_sub23_T_datain = ( (|r_sys_processing_methodID) ? r_sub23_T_datain : 32'h0 ) ;
	assign w_sub23_T_r_w = ( (|r_sys_processing_methodID) ? r_sub23_T_r_w : 1'h0 ) ;
	assign w_sub23_V_addr = ( (|r_sys_processing_methodID) ? r_sub23_V_addr : 9'sh0 ) ;
	assign w_sub23_V_datain = ( (|r_sys_processing_methodID) ? r_sub23_V_datain : 32'h0 ) ;
	assign w_sub23_V_r_w = ( (|r_sys_processing_methodID) ? r_sub23_V_r_w : 1'h0 ) ;
	assign w_sub23_U_addr = ( (|r_sys_processing_methodID) ? r_sub23_U_addr : 9'sh0 ) ;
	assign w_sub23_U_datain = ( (|r_sys_processing_methodID) ? r_sub23_U_datain : 32'h0 ) ;
	assign w_sub23_U_r_w = ( (|r_sys_processing_methodID) ? r_sub23_U_r_w : 1'h0 ) ;
	assign w_sub23_result_addr = ( (|r_sys_processing_methodID) ? r_sub23_result_addr : 9'sh0 ) ;
	assign w_sub23_result_datain = ( (|r_sys_processing_methodID) ? r_sub23_result_datain : 32'h0 ) ;
	assign w_sub23_result_r_w = ( (|r_sys_processing_methodID) ? r_sub23_result_r_w : 1'h0 ) ;
	assign w_sub12_T_addr = ( (|r_sys_processing_methodID) ? r_sub12_T_addr : 9'sh0 ) ;
	assign w_sub12_T_datain = ( (|r_sys_processing_methodID) ? r_sub12_T_datain : 32'h0 ) ;
	assign w_sub12_T_r_w = ( (|r_sys_processing_methodID) ? r_sub12_T_r_w : 1'h0 ) ;
	assign w_sub12_V_addr = ( (|r_sys_processing_methodID) ? r_sub12_V_addr : 9'sh0 ) ;
	assign w_sub12_V_datain = ( (|r_sys_processing_methodID) ? r_sub12_V_datain : 32'h0 ) ;
	assign w_sub12_V_r_w = ( (|r_sys_processing_methodID) ? r_sub12_V_r_w : 1'h0 ) ;
	assign w_sub12_U_addr = ( (|r_sys_processing_methodID) ? r_sub12_U_addr : 9'sh0 ) ;
	assign w_sub12_U_datain = ( (|r_sys_processing_methodID) ? r_sub12_U_datain : 32'h0 ) ;
	assign w_sub12_U_r_w = ( (|r_sys_processing_methodID) ? r_sub12_U_r_w : 1'h0 ) ;
	assign w_sub12_result_addr = ( (|r_sys_processing_methodID) ? r_sub12_result_addr : 9'sh0 ) ;
	assign w_sub12_result_datain = ( (|r_sys_processing_methodID) ? r_sub12_result_datain : 32'h0 ) ;
	assign w_sub12_result_r_w = ( (|r_sys_processing_methodID) ? r_sub12_result_r_w : 1'h0 ) ;
	assign w_sub03_T_addr = ( (|r_sys_processing_methodID) ? r_sub03_T_addr : 9'sh0 ) ;
	assign w_sub03_T_datain = ( (|r_sys_processing_methodID) ? r_sub03_T_datain : 32'h0 ) ;
	assign w_sub03_T_r_w = ( (|r_sys_processing_methodID) ? r_sub03_T_r_w : 1'h0 ) ;
	assign w_sub03_V_addr = ( (|r_sys_processing_methodID) ? r_sub03_V_addr : 9'sh0 ) ;
	assign w_sub03_V_datain = ( (|r_sys_processing_methodID) ? r_sub03_V_datain : 32'h0 ) ;
	assign w_sub03_V_r_w = ( (|r_sys_processing_methodID) ? r_sub03_V_r_w : 1'h0 ) ;
	assign w_sub03_U_addr = ( (|r_sys_processing_methodID) ? r_sub03_U_addr : 9'sh0 ) ;
	assign w_sub03_U_datain = ( (|r_sys_processing_methodID) ? r_sub03_U_datain : 32'h0 ) ;
	assign w_sub03_U_r_w = ( (|r_sys_processing_methodID) ? r_sub03_U_r_w : 1'h0 ) ;
	assign w_sub03_result_addr = ( (|r_sys_processing_methodID) ? r_sub03_result_addr : 9'sh0 ) ;
	assign w_sub03_result_datain = ( (|r_sys_processing_methodID) ? r_sub03_result_datain : 32'h0 ) ;
	assign w_sub03_result_r_w = ( (|r_sys_processing_methodID) ? r_sub03_result_r_w : 1'h0 ) ;
	assign w_sub02_T_addr = ( (|r_sys_processing_methodID) ? r_sub02_T_addr : 9'sh0 ) ;
	assign w_sub02_T_datain = ( (|r_sys_processing_methodID) ? r_sub02_T_datain : 32'h0 ) ;
	assign w_sub02_T_r_w = ( (|r_sys_processing_methodID) ? r_sub02_T_r_w : 1'h0 ) ;
	assign w_sub02_V_addr = ( (|r_sys_processing_methodID) ? r_sub02_V_addr : 9'sh0 ) ;
	assign w_sub02_V_datain = ( (|r_sys_processing_methodID) ? r_sub02_V_datain : 32'h0 ) ;
	assign w_sub02_V_r_w = ( (|r_sys_processing_methodID) ? r_sub02_V_r_w : 1'h0 ) ;
	assign w_sub02_U_addr = ( (|r_sys_processing_methodID) ? r_sub02_U_addr : 9'sh0 ) ;
	assign w_sub02_U_datain = ( (|r_sys_processing_methodID) ? r_sub02_U_datain : 32'h0 ) ;
	assign w_sub02_U_r_w = ( (|r_sys_processing_methodID) ? r_sub02_U_r_w : 1'h0 ) ;
	assign w_sub02_result_addr = ( (|r_sys_processing_methodID) ? r_sub02_result_addr : 9'sh0 ) ;
	assign w_sub02_result_datain = ( (|r_sys_processing_methodID) ? r_sub02_result_datain : 32'h0 ) ;
	assign w_sub02_result_r_w = ( (|r_sys_processing_methodID) ? r_sub02_result_r_w : 1'h0 ) ;
	assign w_sub11_T_addr = ( (|r_sys_processing_methodID) ? r_sub11_T_addr : 9'sh0 ) ;
	assign w_sub11_T_datain = ( (|r_sys_processing_methodID) ? r_sub11_T_datain : 32'h0 ) ;
	assign w_sub11_T_r_w = ( (|r_sys_processing_methodID) ? r_sub11_T_r_w : 1'h0 ) ;
	assign w_sub11_V_addr = ( (|r_sys_processing_methodID) ? r_sub11_V_addr : 9'sh0 ) ;
	assign w_sub11_V_datain = ( (|r_sys_processing_methodID) ? r_sub11_V_datain : 32'h0 ) ;
	assign w_sub11_V_r_w = ( (|r_sys_processing_methodID) ? r_sub11_V_r_w : 1'h0 ) ;
	assign w_sub11_U_addr = ( (|r_sys_processing_methodID) ? r_sub11_U_addr : 9'sh0 ) ;
	assign w_sub11_U_datain = ( (|r_sys_processing_methodID) ? r_sub11_U_datain : 32'h0 ) ;
	assign w_sub11_U_r_w = ( (|r_sys_processing_methodID) ? r_sub11_U_r_w : 1'h0 ) ;
	assign w_sub11_result_addr = ( (|r_sys_processing_methodID) ? r_sub11_result_addr : 9'sh0 ) ;
	assign w_sub11_result_datain = ( (|r_sys_processing_methodID) ? r_sub11_result_datain : 32'h0 ) ;
	assign w_sub11_result_r_w = ( (|r_sys_processing_methodID) ? r_sub11_result_r_w : 1'h0 ) ;
	assign w_sub14_T_addr = ( (|r_sys_processing_methodID) ? r_sub14_T_addr : 9'sh0 ) ;
	assign w_sub14_T_datain = ( (|r_sys_processing_methodID) ? r_sub14_T_datain : 32'h0 ) ;
	assign w_sub14_T_r_w = ( (|r_sys_processing_methodID) ? r_sub14_T_r_w : 1'h0 ) ;
	assign w_sub14_V_addr = ( (|r_sys_processing_methodID) ? r_sub14_V_addr : 9'sh0 ) ;
	assign w_sub14_V_datain = ( (|r_sys_processing_methodID) ? r_sub14_V_datain : 32'h0 ) ;
	assign w_sub14_V_r_w = ( (|r_sys_processing_methodID) ? r_sub14_V_r_w : 1'h0 ) ;
	assign w_sub14_U_addr = ( (|r_sys_processing_methodID) ? r_sub14_U_addr : 9'sh0 ) ;
	assign w_sub14_U_datain = ( (|r_sys_processing_methodID) ? r_sub14_U_datain : 32'h0 ) ;
	assign w_sub14_U_r_w = ( (|r_sys_processing_methodID) ? r_sub14_U_r_w : 1'h0 ) ;
	assign w_sub14_result_addr = ( (|r_sys_processing_methodID) ? r_sub14_result_addr : 9'sh0 ) ;
	assign w_sub14_result_datain = ( (|r_sys_processing_methodID) ? r_sub14_result_datain : 32'h0 ) ;
	assign w_sub14_result_r_w = ( (|r_sys_processing_methodID) ? r_sub14_result_r_w : 1'h0 ) ;
	assign w_sub01_T_addr = ( (|r_sys_processing_methodID) ? r_sub01_T_addr : 9'sh0 ) ;
	assign w_sub01_T_datain = ( (|r_sys_processing_methodID) ? r_sub01_T_datain : 32'h0 ) ;
	assign w_sub01_T_r_w = ( (|r_sys_processing_methodID) ? r_sub01_T_r_w : 1'h0 ) ;
	assign w_sub01_V_addr = ( (|r_sys_processing_methodID) ? r_sub01_V_addr : 9'sh0 ) ;
	assign w_sub01_V_datain = ( (|r_sys_processing_methodID) ? r_sub01_V_datain : 32'h0 ) ;
	assign w_sub01_V_r_w = ( (|r_sys_processing_methodID) ? r_sub01_V_r_w : 1'h0 ) ;
	assign w_sub01_U_addr = ( (|r_sys_processing_methodID) ? r_sub01_U_addr : 9'sh0 ) ;
	assign w_sub01_U_datain = ( (|r_sys_processing_methodID) ? r_sub01_U_datain : 32'h0 ) ;
	assign w_sub01_U_r_w = ( (|r_sys_processing_methodID) ? r_sub01_U_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 9'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub00_T_addr = ( (|r_sys_processing_methodID) ? r_sub00_T_addr : 9'sh0 ) ;
	assign w_sub00_T_datain = ( (|r_sys_processing_methodID) ? r_sub00_T_datain : 32'h0 ) ;
	assign w_sub00_T_r_w = ( (|r_sys_processing_methodID) ? r_sub00_T_r_w : 1'h0 ) ;
	assign w_sub00_V_addr = ( (|r_sys_processing_methodID) ? r_sub00_V_addr : 9'sh0 ) ;
	assign w_sub00_V_datain = ( (|r_sys_processing_methodID) ? r_sub00_V_datain : 32'h0 ) ;
	assign w_sub00_V_r_w = ( (|r_sys_processing_methodID) ? r_sub00_V_r_w : 1'h0 ) ;
	assign w_sub00_U_addr = ( (|r_sys_processing_methodID) ? r_sub00_U_addr : 9'sh0 ) ;
	assign w_sub00_U_datain = ( (|r_sys_processing_methodID) ? r_sub00_U_datain : 32'h0 ) ;
	assign w_sub00_U_r_w = ( (|r_sys_processing_methodID) ? r_sub00_U_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 9'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sub13_T_addr = ( (|r_sys_processing_methodID) ? r_sub13_T_addr : 9'sh0 ) ;
	assign w_sub13_T_datain = ( (|r_sys_processing_methodID) ? r_sub13_T_datain : 32'h0 ) ;
	assign w_sub13_T_r_w = ( (|r_sys_processing_methodID) ? r_sub13_T_r_w : 1'h0 ) ;
	assign w_sub13_V_addr = ( (|r_sys_processing_methodID) ? r_sub13_V_addr : 9'sh0 ) ;
	assign w_sub13_V_datain = ( (|r_sys_processing_methodID) ? r_sub13_V_datain : 32'h0 ) ;
	assign w_sub13_V_r_w = ( (|r_sys_processing_methodID) ? r_sub13_V_r_w : 1'h0 ) ;
	assign w_sub13_U_addr = ( (|r_sys_processing_methodID) ? r_sub13_U_addr : 9'sh0 ) ;
	assign w_sub13_U_datain = ( (|r_sys_processing_methodID) ? r_sub13_U_datain : 32'h0 ) ;
	assign w_sub13_U_r_w = ( (|r_sys_processing_methodID) ? r_sub13_U_r_w : 1'h0 ) ;
	assign w_sub13_result_addr = ( (|r_sys_processing_methodID) ? r_sub13_result_addr : 9'sh0 ) ;
	assign w_sub13_result_datain = ( (|r_sys_processing_methodID) ? r_sub13_result_datain : 32'h0 ) ;
	assign w_sub13_result_r_w = ( (|r_sys_processing_methodID) ? r_sub13_result_r_w : 1'h0 ) ;
	assign w_sub07_T_addr = ( (|r_sys_processing_methodID) ? r_sub07_T_addr : 9'sh0 ) ;
	assign w_sub07_T_datain = ( (|r_sys_processing_methodID) ? r_sub07_T_datain : 32'h0 ) ;
	assign w_sub07_T_r_w = ( (|r_sys_processing_methodID) ? r_sub07_T_r_w : 1'h0 ) ;
	assign w_sub07_V_addr = ( (|r_sys_processing_methodID) ? r_sub07_V_addr : 9'sh0 ) ;
	assign w_sub07_V_datain = ( (|r_sys_processing_methodID) ? r_sub07_V_datain : 32'h0 ) ;
	assign w_sub07_V_r_w = ( (|r_sys_processing_methodID) ? r_sub07_V_r_w : 1'h0 ) ;
	assign w_sub07_U_addr = ( (|r_sys_processing_methodID) ? r_sub07_U_addr : 9'sh0 ) ;
	assign w_sub07_U_datain = ( (|r_sys_processing_methodID) ? r_sub07_U_datain : 32'h0 ) ;
	assign w_sub07_U_r_w = ( (|r_sys_processing_methodID) ? r_sub07_U_r_w : 1'h0 ) ;
	assign w_sub07_result_addr = ( (|r_sys_processing_methodID) ? r_sub07_result_addr : 9'sh0 ) ;
	assign w_sub07_result_datain = ( (|r_sys_processing_methodID) ? r_sub07_result_datain : 32'h0 ) ;
	assign w_sub07_result_r_w = ( (|r_sys_processing_methodID) ? r_sub07_result_r_w : 1'h0 ) ;
	assign w_sub16_T_addr = ( (|r_sys_processing_methodID) ? r_sub16_T_addr : 9'sh0 ) ;
	assign w_sub16_T_datain = ( (|r_sys_processing_methodID) ? r_sub16_T_datain : 32'h0 ) ;
	assign w_sub16_T_r_w = ( (|r_sys_processing_methodID) ? r_sub16_T_r_w : 1'h0 ) ;
	assign w_sub16_V_addr = ( (|r_sys_processing_methodID) ? r_sub16_V_addr : 9'sh0 ) ;
	assign w_sub16_V_datain = ( (|r_sys_processing_methodID) ? r_sub16_V_datain : 32'h0 ) ;
	assign w_sub16_V_r_w = ( (|r_sys_processing_methodID) ? r_sub16_V_r_w : 1'h0 ) ;
	assign w_sub16_U_addr = ( (|r_sys_processing_methodID) ? r_sub16_U_addr : 9'sh0 ) ;
	assign w_sub16_U_datain = ( (|r_sys_processing_methodID) ? r_sub16_U_datain : 32'h0 ) ;
	assign w_sub16_U_r_w = ( (|r_sys_processing_methodID) ? r_sub16_U_r_w : 1'h0 ) ;
	assign w_sub16_result_addr = ( (|r_sys_processing_methodID) ? r_sub16_result_addr : 9'sh0 ) ;
	assign w_sub16_result_datain = ( (|r_sys_processing_methodID) ? r_sub16_result_datain : 32'h0 ) ;
	assign w_sub16_result_r_w = ( (|r_sys_processing_methodID) ? r_sub16_result_r_w : 1'h0 ) ;
	assign w_sub06_T_addr = ( (|r_sys_processing_methodID) ? r_sub06_T_addr : 9'sh0 ) ;
	assign w_sub06_T_datain = ( (|r_sys_processing_methodID) ? r_sub06_T_datain : 32'h0 ) ;
	assign w_sub06_T_r_w = ( (|r_sys_processing_methodID) ? r_sub06_T_r_w : 1'h0 ) ;
	assign w_sub06_V_addr = ( (|r_sys_processing_methodID) ? r_sub06_V_addr : 9'sh0 ) ;
	assign w_sub06_V_datain = ( (|r_sys_processing_methodID) ? r_sub06_V_datain : 32'h0 ) ;
	assign w_sub06_V_r_w = ( (|r_sys_processing_methodID) ? r_sub06_V_r_w : 1'h0 ) ;
	assign w_sub06_U_addr = ( (|r_sys_processing_methodID) ? r_sub06_U_addr : 9'sh0 ) ;
	assign w_sub06_U_datain = ( (|r_sys_processing_methodID) ? r_sub06_U_datain : 32'h0 ) ;
	assign w_sub06_U_r_w = ( (|r_sys_processing_methodID) ? r_sub06_U_r_w : 1'h0 ) ;
	assign w_sub06_result_addr = ( (|r_sys_processing_methodID) ? r_sub06_result_addr : 9'sh0 ) ;
	assign w_sub06_result_datain = ( (|r_sys_processing_methodID) ? r_sub06_result_datain : 32'h0 ) ;
	assign w_sub06_result_r_w = ( (|r_sys_processing_methodID) ? r_sub06_result_r_w : 1'h0 ) ;
	assign w_sub15_T_addr = ( (|r_sys_processing_methodID) ? r_sub15_T_addr : 9'sh0 ) ;
	assign w_sub15_T_datain = ( (|r_sys_processing_methodID) ? r_sub15_T_datain : 32'h0 ) ;
	assign w_sub15_T_r_w = ( (|r_sys_processing_methodID) ? r_sub15_T_r_w : 1'h0 ) ;
	assign w_sub15_V_addr = ( (|r_sys_processing_methodID) ? r_sub15_V_addr : 9'sh0 ) ;
	assign w_sub15_V_datain = ( (|r_sys_processing_methodID) ? r_sub15_V_datain : 32'h0 ) ;
	assign w_sub15_V_r_w = ( (|r_sys_processing_methodID) ? r_sub15_V_r_w : 1'h0 ) ;
	assign w_sub15_U_addr = ( (|r_sys_processing_methodID) ? r_sub15_U_addr : 9'sh0 ) ;
	assign w_sub15_U_datain = ( (|r_sys_processing_methodID) ? r_sub15_U_datain : 32'h0 ) ;
	assign w_sub15_U_r_w = ( (|r_sys_processing_methodID) ? r_sub15_U_r_w : 1'h0 ) ;
	assign w_sub15_result_addr = ( (|r_sys_processing_methodID) ? r_sub15_result_addr : 9'sh0 ) ;
	assign w_sub15_result_datain = ( (|r_sys_processing_methodID) ? r_sub15_result_datain : 32'h0 ) ;
	assign w_sub15_result_r_w = ( (|r_sys_processing_methodID) ? r_sub15_result_r_w : 1'h0 ) ;
	assign w_sub05_T_addr = ( (|r_sys_processing_methodID) ? r_sub05_T_addr : 9'sh0 ) ;
	assign w_sub05_T_datain = ( (|r_sys_processing_methodID) ? r_sub05_T_datain : 32'h0 ) ;
	assign w_sub05_T_r_w = ( (|r_sys_processing_methodID) ? r_sub05_T_r_w : 1'h0 ) ;
	assign w_sub05_V_addr = ( (|r_sys_processing_methodID) ? r_sub05_V_addr : 9'sh0 ) ;
	assign w_sub05_V_datain = ( (|r_sys_processing_methodID) ? r_sub05_V_datain : 32'h0 ) ;
	assign w_sub05_V_r_w = ( (|r_sys_processing_methodID) ? r_sub05_V_r_w : 1'h0 ) ;
	assign w_sub05_U_addr = ( (|r_sys_processing_methodID) ? r_sub05_U_addr : 9'sh0 ) ;
	assign w_sub05_U_datain = ( (|r_sys_processing_methodID) ? r_sub05_U_datain : 32'h0 ) ;
	assign w_sub05_U_r_w = ( (|r_sys_processing_methodID) ? r_sub05_U_r_w : 1'h0 ) ;
	assign w_sub05_result_addr = ( (|r_sys_processing_methodID) ? r_sub05_result_addr : 9'sh0 ) ;
	assign w_sub05_result_datain = ( (|r_sys_processing_methodID) ? r_sub05_result_datain : 32'h0 ) ;
	assign w_sub05_result_r_w = ( (|r_sys_processing_methodID) ? r_sub05_result_r_w : 1'h0 ) ;
	assign w_sub18_T_addr = ( (|r_sys_processing_methodID) ? r_sub18_T_addr : 9'sh0 ) ;
	assign w_sub18_T_datain = ( (|r_sys_processing_methodID) ? r_sub18_T_datain : 32'h0 ) ;
	assign w_sub18_T_r_w = ( (|r_sys_processing_methodID) ? r_sub18_T_r_w : 1'h0 ) ;
	assign w_sub18_V_addr = ( (|r_sys_processing_methodID) ? r_sub18_V_addr : 9'sh0 ) ;
	assign w_sub18_V_datain = ( (|r_sys_processing_methodID) ? r_sub18_V_datain : 32'h0 ) ;
	assign w_sub18_V_r_w = ( (|r_sys_processing_methodID) ? r_sub18_V_r_w : 1'h0 ) ;
	assign w_sub18_U_addr = ( (|r_sys_processing_methodID) ? r_sub18_U_addr : 9'sh0 ) ;
	assign w_sub18_U_datain = ( (|r_sys_processing_methodID) ? r_sub18_U_datain : 32'h0 ) ;
	assign w_sub18_U_r_w = ( (|r_sys_processing_methodID) ? r_sub18_U_r_w : 1'h0 ) ;
	assign w_sub18_result_addr = ( (|r_sys_processing_methodID) ? r_sub18_result_addr : 9'sh0 ) ;
	assign w_sub18_result_datain = ( (|r_sys_processing_methodID) ? r_sub18_result_datain : 32'h0 ) ;
	assign w_sub18_result_r_w = ( (|r_sys_processing_methodID) ? r_sub18_result_r_w : 1'h0 ) ;
	assign w_sub04_T_addr = ( (|r_sys_processing_methodID) ? r_sub04_T_addr : 9'sh0 ) ;
	assign w_sub04_T_datain = ( (|r_sys_processing_methodID) ? r_sub04_T_datain : 32'h0 ) ;
	assign w_sub04_T_r_w = ( (|r_sys_processing_methodID) ? r_sub04_T_r_w : 1'h0 ) ;
	assign w_sub04_V_addr = ( (|r_sys_processing_methodID) ? r_sub04_V_addr : 9'sh0 ) ;
	assign w_sub04_V_datain = ( (|r_sys_processing_methodID) ? r_sub04_V_datain : 32'h0 ) ;
	assign w_sub04_V_r_w = ( (|r_sys_processing_methodID) ? r_sub04_V_r_w : 1'h0 ) ;
	assign w_sub04_U_addr = ( (|r_sys_processing_methodID) ? r_sub04_U_addr : 9'sh0 ) ;
	assign w_sub04_U_datain = ( (|r_sys_processing_methodID) ? r_sub04_U_datain : 32'h0 ) ;
	assign w_sub04_U_r_w = ( (|r_sys_processing_methodID) ? r_sub04_U_r_w : 1'h0 ) ;
	assign w_sub04_result_addr = ( (|r_sys_processing_methodID) ? r_sub04_result_addr : 9'sh0 ) ;
	assign w_sub04_result_datain = ( (|r_sys_processing_methodID) ? r_sub04_result_datain : 32'h0 ) ;
	assign w_sub04_result_r_w = ( (|r_sys_processing_methodID) ? r_sub04_result_r_w : 1'h0 ) ;
	assign w_sub17_T_addr = ( (|r_sys_processing_methodID) ? r_sub17_T_addr : 9'sh0 ) ;
	assign w_sub17_T_datain = ( (|r_sys_processing_methodID) ? r_sub17_T_datain : 32'h0 ) ;
	assign w_sub17_T_r_w = ( (|r_sys_processing_methodID) ? r_sub17_T_r_w : 1'h0 ) ;
	assign w_sub17_V_addr = ( (|r_sys_processing_methodID) ? r_sub17_V_addr : 9'sh0 ) ;
	assign w_sub17_V_datain = ( (|r_sys_processing_methodID) ? r_sub17_V_datain : 32'h0 ) ;
	assign w_sub17_V_r_w = ( (|r_sys_processing_methodID) ? r_sub17_V_r_w : 1'h0 ) ;
	assign w_sub17_U_addr = ( (|r_sys_processing_methodID) ? r_sub17_U_addr : 9'sh0 ) ;
	assign w_sub17_U_datain = ( (|r_sys_processing_methodID) ? r_sub17_U_datain : 32'h0 ) ;
	assign w_sub17_U_r_w = ( (|r_sys_processing_methodID) ? r_sub17_U_r_w : 1'h0 ) ;
	assign w_sub17_result_addr = ( (|r_sys_processing_methodID) ? r_sub17_result_addr : 9'sh0 ) ;
	assign w_sub17_result_datain = ( (|r_sys_processing_methodID) ? r_sub17_result_datain : 32'h0 ) ;
	assign w_sub17_result_r_w = ( (|r_sys_processing_methodID) ? r_sub17_result_r_w : 1'h0 ) ;
	assign w_sub10_T_addr = ( (|r_sys_processing_methodID) ? r_sub10_T_addr : 9'sh0 ) ;
	assign w_sub10_T_datain = ( (|r_sys_processing_methodID) ? r_sub10_T_datain : 32'h0 ) ;
	assign w_sub10_T_r_w = ( (|r_sys_processing_methodID) ? r_sub10_T_r_w : 1'h0 ) ;
	assign w_sub10_V_addr = ( (|r_sys_processing_methodID) ? r_sub10_V_addr : 9'sh0 ) ;
	assign w_sub10_V_datain = ( (|r_sys_processing_methodID) ? r_sub10_V_datain : 32'h0 ) ;
	assign w_sub10_V_r_w = ( (|r_sys_processing_methodID) ? r_sub10_V_r_w : 1'h0 ) ;
	assign w_sub10_U_addr = ( (|r_sys_processing_methodID) ? r_sub10_U_addr : 9'sh0 ) ;
	assign w_sub10_U_datain = ( (|r_sys_processing_methodID) ? r_sub10_U_datain : 32'h0 ) ;
	assign w_sub10_U_r_w = ( (|r_sys_processing_methodID) ? r_sub10_U_r_w : 1'h0 ) ;
	assign w_sub10_result_addr = ( (|r_sys_processing_methodID) ? r_sub10_result_addr : 9'sh0 ) ;
	assign w_sub10_result_datain = ( (|r_sys_processing_methodID) ? r_sub10_result_datain : 32'h0 ) ;
	assign w_sub10_result_r_w = ( (|r_sys_processing_methodID) ? r_sub10_result_r_w : 1'h0 ) ;
	assign w_sub20_T_addr = ( (|r_sys_processing_methodID) ? r_sub20_T_addr : 9'sh0 ) ;
	assign w_sub20_T_datain = ( (|r_sys_processing_methodID) ? r_sub20_T_datain : 32'h0 ) ;
	assign w_sub20_T_r_w = ( (|r_sys_processing_methodID) ? r_sub20_T_r_w : 1'h0 ) ;
	assign w_sub20_V_addr = ( (|r_sys_processing_methodID) ? r_sub20_V_addr : 9'sh0 ) ;
	assign w_sub20_V_datain = ( (|r_sys_processing_methodID) ? r_sub20_V_datain : 32'h0 ) ;
	assign w_sub20_V_r_w = ( (|r_sys_processing_methodID) ? r_sub20_V_r_w : 1'h0 ) ;
	assign w_sub20_U_addr = ( (|r_sys_processing_methodID) ? r_sub20_U_addr : 9'sh0 ) ;
	assign w_sub20_U_datain = ( (|r_sys_processing_methodID) ? r_sub20_U_datain : 32'h0 ) ;
	assign w_sub20_U_r_w = ( (|r_sys_processing_methodID) ? r_sub20_U_r_w : 1'h0 ) ;
	assign w_sub20_result_addr = ( (|r_sys_processing_methodID) ? r_sub20_result_addr : 9'sh0 ) ;
	assign w_sub20_result_datain = ( (|r_sys_processing_methodID) ? r_sub20_result_datain : 32'h0 ) ;
	assign w_sub20_result_r_w = ( (|r_sys_processing_methodID) ? r_sub20_result_r_w : 1'h0 ) ;
	assign w_sub21_T_addr = ( (|r_sys_processing_methodID) ? r_sub21_T_addr : 9'sh0 ) ;
	assign w_sub21_T_datain = ( (|r_sys_processing_methodID) ? r_sub21_T_datain : 32'h0 ) ;
	assign w_sub21_T_r_w = ( (|r_sys_processing_methodID) ? r_sub21_T_r_w : 1'h0 ) ;
	assign w_sub21_V_addr = ( (|r_sys_processing_methodID) ? r_sub21_V_addr : 9'sh0 ) ;
	assign w_sub21_V_datain = ( (|r_sys_processing_methodID) ? r_sub21_V_datain : 32'h0 ) ;
	assign w_sub21_V_r_w = ( (|r_sys_processing_methodID) ? r_sub21_V_r_w : 1'h0 ) ;
	assign w_sub21_U_addr = ( (|r_sys_processing_methodID) ? r_sub21_U_addr : 9'sh0 ) ;
	assign w_sub21_U_datain = ( (|r_sys_processing_methodID) ? r_sub21_U_datain : 32'h0 ) ;
	assign w_sub21_U_r_w = ( (|r_sys_processing_methodID) ? r_sub21_U_r_w : 1'h0 ) ;
	assign w_sub21_result_addr = ( (|r_sys_processing_methodID) ? r_sub21_result_addr : 9'sh0 ) ;
	assign w_sub21_result_datain = ( (|r_sys_processing_methodID) ? r_sub21_result_datain : 32'h0 ) ;
	assign w_sub21_result_r_w = ( (|r_sys_processing_methodID) ? r_sub21_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh00000014;
	assign w_sys_tmp3 = 32'sh00000015;
	assign w_sys_tmp5 = 32'h3a03126f;
	assign w_sys_tmp6 = 32'sh00000002;
	assign w_sys_tmp7 = 32'h3e4ccccd;
	assign w_sys_tmp8 = 32'h3d4ccccd;
	assign w_sys_tmp9 = 32'h3aa3d70b;
	assign w_sys_tmp10 = 32'h3ba3d70b;
	assign w_sys_tmp11 = 32'h3c4ccccc;
	assign w_sys_tmp12 = 32'h3e4ccccc;
	assign w_sys_tmp13 = ( !w_sys_tmp14 );
	assign w_sys_tmp14 = (r_run_my_33 < r_run_k_29);
	assign w_sys_tmp15 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp16 = ( !w_sys_tmp17 );
	assign w_sys_tmp17 = (r_run_mx_32 < r_run_j_30);
	assign w_sys_tmp19 = w_ip_MultFloat_product_0;
	assign w_sys_tmp20 = w_ip_FixedToFloat_floating_0;
	assign w_sys_tmp21 = (r_run_k_29 - w_sys_intOne);
	assign w_sys_tmp23 = (w_sys_tmp24 + r_run_k_29);
	assign w_sys_tmp24 = (r_run_j_30 * w_sys_tmp25);
	assign w_sys_tmp25 = 32'sh00000015;
	assign w_sys_tmp26 = 32'h0;
	assign w_sys_tmp28 = (w_sys_tmp29 + r_run_k_29);
	assign w_sys_tmp29 = (r_run_copy2_j_47 * w_sys_tmp25);
	assign w_sys_tmp33 = (w_sys_tmp34 + r_run_k_29);
	assign w_sys_tmp34 = (r_run_copy1_j_46 * w_sys_tmp25);
	assign w_sys_tmp37 = 32'h42200000;
	assign w_sys_tmp38 = w_sys_tmp19;
	assign w_sys_tmp39 = 32'h3f800000;
	assign w_sys_tmp42 = (w_sys_tmp43 + r_run_k_29);
	assign w_sys_tmp43 = (r_run_copy0_j_45 * w_sys_tmp25);
	assign w_sys_tmp46 = (r_run_copy0_j_45 + w_sys_intOne);
	assign w_sys_tmp47 = (r_run_copy1_j_46 + w_sys_intOne);
	assign w_sys_tmp48 = (r_run_copy2_j_47 + w_sys_intOne);
	assign w_sys_tmp49 = (r_run_j_30 + w_sys_intOne);
	assign w_sys_tmp129 = r_sys_tmp4_float;
	assign w_sys_tmp227 = ( !w_sys_tmp228 );
	assign w_sys_tmp228 = (w_sys_tmp229 < r_run_k_29);
	assign w_sys_tmp229 = 32'sh00000006;
	assign w_sys_tmp232 = (w_sys_tmp233 + r_run_k_29);
	assign w_sys_tmp233 = 32'sh00000015;
	assign w_sys_tmp234 = w_fld_U_2_dataout_1;
	assign w_sys_tmp238 = (w_sys_tmp239 + r_run_k_29);
	assign w_sys_tmp239 = 32'sh0000002a;
	assign w_sys_tmp244 = (w_sys_tmp245 + r_run_k_29);
	assign w_sys_tmp245 = 32'sh0000003f;
	assign w_sys_tmp250 = (w_sys_tmp251 + r_run_k_29);
	assign w_sys_tmp251 = 32'sh00000054;
	assign w_sys_tmp256 = (w_sys_tmp257 + r_run_k_29);
	assign w_sys_tmp257 = 32'sh00000069;
	assign w_sys_tmp262 = (w_sys_tmp263 + r_run_k_29);
	assign w_sys_tmp263 = 32'sh0000007e;
	assign w_sys_tmp280 = (w_sys_tmp281 + r_run_k_29);
	assign w_sys_tmp281 = 32'sh00000093;
	assign w_sys_tmp286 = (w_sys_tmp287 + r_run_k_29);
	assign w_sys_tmp287 = 32'sh000000a8;
	assign w_sys_tmp292 = (w_sys_tmp293 + r_run_k_29);
	assign w_sys_tmp293 = 32'sh000000bd;
	assign w_sys_tmp298 = (w_sys_tmp299 + r_run_k_29);
	assign w_sys_tmp299 = 32'sh000000d2;
	assign w_sys_tmp316 = (w_sys_tmp317 + r_run_k_29);
	assign w_sys_tmp317 = 32'sh000000e7;
	assign w_sys_tmp322 = (w_sys_tmp323 + r_run_k_29);
	assign w_sys_tmp323 = 32'sh000000fc;
	assign w_sys_tmp328 = (w_sys_tmp329 + r_run_k_29);
	assign w_sys_tmp329 = 32'sh00000111;
	assign w_sys_tmp334 = (w_sys_tmp335 + r_run_k_29);
	assign w_sys_tmp335 = 32'sh00000126;
	assign w_sys_tmp352 = (w_sys_tmp353 + r_run_k_29);
	assign w_sys_tmp353 = 32'sh0000013b;
	assign w_sys_tmp358 = (w_sys_tmp359 + r_run_k_29);
	assign w_sys_tmp359 = 32'sh00000150;
	assign w_sys_tmp364 = (w_sys_tmp365 + r_run_k_29);
	assign w_sys_tmp365 = 32'sh00000165;
	assign w_sys_tmp376 = (w_sys_tmp377 + r_run_k_29);
	assign w_sys_tmp377 = 32'sh0000017a;
	assign w_sys_tmp382 = (w_sys_tmp383 + r_run_k_29);
	assign w_sys_tmp383 = 32'sh0000018f;
	assign w_sys_tmp388 = (w_sys_tmp389 + r_run_k_29);
	assign w_sys_tmp389 = 32'sh000001a4;
	assign w_sys_tmp396 = w_fld_V_3_dataout_1;
	assign w_sys_tmp556 = (w_sys_tmp557 + r_run_k_29);
	assign w_sys_tmp557 = 32'sh00000019;
	assign w_sys_tmp562 = (w_sys_tmp563 + r_run_k_29);
	assign w_sys_tmp563 = 32'sh0000002e;
	assign w_sys_tmp568 = (w_sys_tmp569 + r_run_k_29);
	assign w_sys_tmp569 = 32'sh00000043;
	assign w_sys_tmp574 = (w_sys_tmp575 + r_run_k_29);
	assign w_sys_tmp575 = 32'sh00000058;
	assign w_sys_tmp580 = (w_sys_tmp581 + r_run_k_29);
	assign w_sys_tmp581 = 32'sh0000006d;
	assign w_sys_tmp586 = (w_sys_tmp587 + r_run_k_29);
	assign w_sys_tmp587 = 32'sh00000082;
	assign w_sys_tmp604 = (w_sys_tmp605 + r_run_k_29);
	assign w_sys_tmp605 = 32'sh00000097;
	assign w_sys_tmp610 = (w_sys_tmp611 + r_run_k_29);
	assign w_sys_tmp611 = 32'sh000000ac;
	assign w_sys_tmp616 = (w_sys_tmp617 + r_run_k_29);
	assign w_sys_tmp617 = 32'sh000000c1;
	assign w_sys_tmp622 = (w_sys_tmp623 + r_run_k_29);
	assign w_sys_tmp623 = 32'sh000000d6;
	assign w_sys_tmp640 = (w_sys_tmp641 + r_run_k_29);
	assign w_sys_tmp641 = 32'sh000000eb;
	assign w_sys_tmp646 = (w_sys_tmp647 + r_run_k_29);
	assign w_sys_tmp647 = 32'sh00000100;
	assign w_sys_tmp652 = (w_sys_tmp653 + r_run_k_29);
	assign w_sys_tmp653 = 32'sh00000115;
	assign w_sys_tmp658 = (w_sys_tmp659 + r_run_k_29);
	assign w_sys_tmp659 = 32'sh0000012a;
	assign w_sys_tmp676 = (w_sys_tmp677 + r_run_k_29);
	assign w_sys_tmp677 = 32'sh0000013f;
	assign w_sys_tmp682 = (w_sys_tmp683 + r_run_k_29);
	assign w_sys_tmp683 = 32'sh00000154;
	assign w_sys_tmp688 = (w_sys_tmp689 + r_run_k_29);
	assign w_sys_tmp689 = 32'sh00000169;
	assign w_sys_tmp700 = (w_sys_tmp701 + r_run_k_29);
	assign w_sys_tmp701 = 32'sh0000017e;
	assign w_sys_tmp706 = (w_sys_tmp707 + r_run_k_29);
	assign w_sys_tmp707 = 32'sh00000193;
	assign w_sys_tmp712 = (w_sys_tmp713 + r_run_k_29);
	assign w_sys_tmp713 = 32'sh000001a8;
	assign w_sys_tmp880 = (w_sys_tmp881 + r_run_k_29);
	assign w_sys_tmp881 = 32'sh0000001d;
	assign w_sys_tmp886 = (w_sys_tmp887 + r_run_k_29);
	assign w_sys_tmp887 = 32'sh00000032;
	assign w_sys_tmp892 = (w_sys_tmp893 + r_run_k_29);
	assign w_sys_tmp893 = 32'sh00000047;
	assign w_sys_tmp898 = (w_sys_tmp899 + r_run_k_29);
	assign w_sys_tmp899 = 32'sh0000005c;
	assign w_sys_tmp904 = (w_sys_tmp905 + r_run_k_29);
	assign w_sys_tmp905 = 32'sh00000071;
	assign w_sys_tmp910 = (w_sys_tmp911 + r_run_k_29);
	assign w_sys_tmp911 = 32'sh00000086;
	assign w_sys_tmp928 = (w_sys_tmp929 + r_run_k_29);
	assign w_sys_tmp929 = 32'sh0000009b;
	assign w_sys_tmp934 = (w_sys_tmp935 + r_run_k_29);
	assign w_sys_tmp935 = 32'sh000000b0;
	assign w_sys_tmp940 = (w_sys_tmp941 + r_run_k_29);
	assign w_sys_tmp941 = 32'sh000000c5;
	assign w_sys_tmp946 = (w_sys_tmp947 + r_run_k_29);
	assign w_sys_tmp947 = 32'sh000000da;
	assign w_sys_tmp964 = (w_sys_tmp965 + r_run_k_29);
	assign w_sys_tmp965 = 32'sh000000ef;
	assign w_sys_tmp970 = (w_sys_tmp971 + r_run_k_29);
	assign w_sys_tmp971 = 32'sh00000104;
	assign w_sys_tmp976 = (w_sys_tmp977 + r_run_k_29);
	assign w_sys_tmp977 = 32'sh00000119;
	assign w_sys_tmp982 = (w_sys_tmp983 + r_run_k_29);
	assign w_sys_tmp983 = 32'sh0000012e;
	assign w_sys_tmp1000 = (w_sys_tmp1001 + r_run_k_29);
	assign w_sys_tmp1001 = 32'sh00000143;
	assign w_sys_tmp1006 = (w_sys_tmp1007 + r_run_k_29);
	assign w_sys_tmp1007 = 32'sh00000158;
	assign w_sys_tmp1012 = (w_sys_tmp1013 + r_run_k_29);
	assign w_sys_tmp1013 = 32'sh0000016d;
	assign w_sys_tmp1024 = (w_sys_tmp1025 + r_run_k_29);
	assign w_sys_tmp1025 = 32'sh00000182;
	assign w_sys_tmp1030 = (w_sys_tmp1031 + r_run_k_29);
	assign w_sys_tmp1031 = 32'sh00000197;
	assign w_sys_tmp1036 = (w_sys_tmp1037 + r_run_k_29);
	assign w_sys_tmp1037 = 32'sh000001ac;
	assign w_sys_tmp1204 = (w_sys_tmp1205 + r_run_k_29);
	assign w_sys_tmp1205 = 32'sh00000021;
	assign w_sys_tmp1210 = (w_sys_tmp1211 + r_run_k_29);
	assign w_sys_tmp1211 = 32'sh00000036;
	assign w_sys_tmp1216 = (w_sys_tmp1217 + r_run_k_29);
	assign w_sys_tmp1217 = 32'sh0000004b;
	assign w_sys_tmp1222 = (w_sys_tmp1223 + r_run_k_29);
	assign w_sys_tmp1223 = 32'sh00000060;
	assign w_sys_tmp1228 = (w_sys_tmp1229 + r_run_k_29);
	assign w_sys_tmp1229 = 32'sh00000075;
	assign w_sys_tmp1234 = (w_sys_tmp1235 + r_run_k_29);
	assign w_sys_tmp1235 = 32'sh0000008a;
	assign w_sys_tmp1252 = (w_sys_tmp1253 + r_run_k_29);
	assign w_sys_tmp1253 = 32'sh0000009f;
	assign w_sys_tmp1258 = (w_sys_tmp1259 + r_run_k_29);
	assign w_sys_tmp1259 = 32'sh000000b4;
	assign w_sys_tmp1264 = (w_sys_tmp1265 + r_run_k_29);
	assign w_sys_tmp1265 = 32'sh000000c9;
	assign w_sys_tmp1270 = (w_sys_tmp1271 + r_run_k_29);
	assign w_sys_tmp1271 = 32'sh000000de;
	assign w_sys_tmp1288 = (w_sys_tmp1289 + r_run_k_29);
	assign w_sys_tmp1289 = 32'sh000000f3;
	assign w_sys_tmp1294 = (w_sys_tmp1295 + r_run_k_29);
	assign w_sys_tmp1295 = 32'sh00000108;
	assign w_sys_tmp1300 = (w_sys_tmp1301 + r_run_k_29);
	assign w_sys_tmp1301 = 32'sh0000011d;
	assign w_sys_tmp1306 = (w_sys_tmp1307 + r_run_k_29);
	assign w_sys_tmp1307 = 32'sh00000132;
	assign w_sys_tmp1324 = (w_sys_tmp1325 + r_run_k_29);
	assign w_sys_tmp1325 = 32'sh00000147;
	assign w_sys_tmp1330 = (w_sys_tmp1331 + r_run_k_29);
	assign w_sys_tmp1331 = 32'sh0000015c;
	assign w_sys_tmp1336 = (w_sys_tmp1337 + r_run_k_29);
	assign w_sys_tmp1337 = 32'sh00000171;
	assign w_sys_tmp1348 = (w_sys_tmp1349 + r_run_k_29);
	assign w_sys_tmp1349 = 32'sh00000186;
	assign w_sys_tmp1354 = (w_sys_tmp1355 + r_run_k_29);
	assign w_sys_tmp1355 = 32'sh0000019b;
	assign w_sys_tmp1360 = (w_sys_tmp1361 + r_run_k_29);
	assign w_sys_tmp1361 = 32'sh000001b0;
	assign w_sys_tmp1527 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp1528 = 32'sh00000011;
	assign w_sys_tmp1529 = ( !w_sys_tmp1530 );
	assign w_sys_tmp1530 = (w_sys_tmp1531 < r_run_k_29);
	assign w_sys_tmp1531 = 32'sh00000015;
	assign w_sys_tmp1534 = (w_sys_tmp1535 + r_run_k_29);
	assign w_sys_tmp1535 = 32'sh00000015;
	assign w_sys_tmp1536 = w_fld_U_2_dataout_1;
	assign w_sys_tmp1540 = (w_sys_tmp1541 + r_run_k_29);
	assign w_sys_tmp1541 = 32'sh0000002a;
	assign w_sys_tmp1546 = (w_sys_tmp1547 + r_run_k_29);
	assign w_sys_tmp1547 = 32'sh0000003f;
	assign w_sys_tmp1552 = (w_sys_tmp1553 + r_run_k_29);
	assign w_sys_tmp1553 = 32'sh00000054;
	assign w_sys_tmp1558 = (w_sys_tmp1559 + r_run_k_29);
	assign w_sys_tmp1559 = 32'sh00000069;
	assign w_sys_tmp1564 = (w_sys_tmp1565 + r_run_k_29);
	assign w_sys_tmp1565 = 32'sh0000007e;
	assign w_sys_tmp1582 = (w_sys_tmp1583 + r_run_k_29);
	assign w_sys_tmp1583 = 32'sh00000093;
	assign w_sys_tmp1588 = (w_sys_tmp1589 + r_run_k_29);
	assign w_sys_tmp1589 = 32'sh000000a8;
	assign w_sys_tmp1594 = (w_sys_tmp1595 + r_run_k_29);
	assign w_sys_tmp1595 = 32'sh000000bd;
	assign w_sys_tmp1600 = (w_sys_tmp1601 + r_run_k_29);
	assign w_sys_tmp1601 = 32'sh000000d2;
	assign w_sys_tmp1618 = (w_sys_tmp1619 + r_run_k_29);
	assign w_sys_tmp1619 = 32'sh000000e7;
	assign w_sys_tmp1624 = (w_sys_tmp1625 + r_run_k_29);
	assign w_sys_tmp1625 = 32'sh000000fc;
	assign w_sys_tmp1630 = (w_sys_tmp1631 + r_run_k_29);
	assign w_sys_tmp1631 = 32'sh00000111;
	assign w_sys_tmp1636 = (w_sys_tmp1637 + r_run_k_29);
	assign w_sys_tmp1637 = 32'sh00000126;
	assign w_sys_tmp1654 = (w_sys_tmp1655 + r_run_k_29);
	assign w_sys_tmp1655 = 32'sh0000013b;
	assign w_sys_tmp1660 = (w_sys_tmp1661 + r_run_k_29);
	assign w_sys_tmp1661 = 32'sh00000150;
	assign w_sys_tmp1666 = (w_sys_tmp1667 + r_run_k_29);
	assign w_sys_tmp1667 = 32'sh00000165;
	assign w_sys_tmp1678 = (w_sys_tmp1679 + r_run_k_29);
	assign w_sys_tmp1679 = 32'sh0000017a;
	assign w_sys_tmp1684 = (w_sys_tmp1685 + r_run_k_29);
	assign w_sys_tmp1685 = 32'sh0000018f;
	assign w_sys_tmp1690 = (w_sys_tmp1691 + r_run_k_29);
	assign w_sys_tmp1691 = 32'sh000001a4;
	assign w_sys_tmp1698 = w_fld_V_3_dataout_1;
	assign w_sys_tmp1857 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp1858 = ( !w_sys_tmp1859 );
	assign w_sys_tmp1859 = (r_run_nlast_44 < r_run_n_31);
	assign w_sys_tmp1860 = (r_run_n_31 + w_sys_intOne);
	assign w_sys_tmp1861 = ( !w_sys_tmp1862 );
	assign w_sys_tmp1862 = (r_run_my_33 < r_run_k_29);
	assign w_sys_tmp1865 = (w_sys_tmp1866 + r_run_k_29);
	assign w_sys_tmp1866 = 32'sh00000015;
	assign w_sys_tmp1867 = 32'h0;
	assign w_sys_tmp1869 = (w_sys_tmp1870 + r_run_k_29);
	assign w_sys_tmp1870 = (r_run_mx_32 * w_sys_tmp1866);
	assign w_sys_tmp1872 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1873 = (w_sys_tmp1874 + r_run_k_29);
	assign w_sys_tmp1874 = (w_sys_tmp1875 * w_sys_tmp1866);
	assign w_sys_tmp1875 = (r_run_mx_32 - w_sys_intOne);
	assign w_sys_tmp1877 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp1878 = ( !w_sys_tmp1879 );
	assign w_sys_tmp1879 = (r_run_mx_32 < r_run_j_30);
	assign w_sys_tmp1882 = (w_sys_tmp1883 + w_sys_intOne);
	assign w_sys_tmp1883 = (r_run_j_30 * w_sys_tmp1884);
	assign w_sys_tmp1884 = 32'sh00000015;
	assign w_sys_tmp1885 = 32'h0;
	assign w_sys_tmp1887 = (w_sys_tmp1888 + r_run_my_33);
	assign w_sys_tmp1888 = (r_run_copy0_j_48 * w_sys_tmp1884);
	assign w_sys_tmp1891 = (r_run_copy0_j_48 + w_sys_intOne);
	assign w_sys_tmp1892 = (r_run_j_30 + w_sys_intOne);
	assign w_sys_tmp1965 = w_ip_DivInt_quotient_0;
	assign w_sys_tmp1966 = 32'sh00000004;
	assign w_sys_tmp1967 = ( !w_sys_tmp1968 );
	assign w_sys_tmp1968 = (w_sys_tmp1969 < r_run_j_30);
	assign w_sys_tmp1969 = w_ip_DivInt_quotient_0;
	assign w_sys_tmp1970 = 32'sh00000002;
	assign w_sys_tmp1973 = (w_sys_tmp1974 + w_sys_intOne);
	assign w_sys_tmp1974 = (r_run_j_30 * w_sys_tmp1975);
	assign w_sys_tmp1975 = 32'sh00000015;
	assign w_sys_tmp1976 = 32'h3f800000;
	assign w_sys_tmp1977 = (r_run_j_30 + w_sys_intOne);
	assign w_sys_tmp2014 = ( !w_sys_tmp2015 );
	assign w_sys_tmp2015 = (w_sys_tmp2016 < r_run_k_29);
	assign w_sys_tmp2016 = 32'sh00000006;
	assign w_sys_tmp2019 = (w_sys_tmp2020 + r_run_k_29);
	assign w_sys_tmp2020 = 32'sh00000015;
	assign w_sys_tmp2021 = w_fld_T_0_dataout_1;
	assign w_sys_tmp2025 = (w_sys_tmp2026 + r_run_k_29);
	assign w_sys_tmp2026 = 32'sh0000002a;
	assign w_sys_tmp2031 = (w_sys_tmp2032 + r_run_k_29);
	assign w_sys_tmp2032 = 32'sh0000003f;
	assign w_sys_tmp2037 = (w_sys_tmp2038 + r_run_k_29);
	assign w_sys_tmp2038 = 32'sh00000054;
	assign w_sys_tmp2043 = (w_sys_tmp2044 + r_run_k_29);
	assign w_sys_tmp2044 = 32'sh00000069;
	assign w_sys_tmp2049 = (w_sys_tmp2050 + r_run_k_29);
	assign w_sys_tmp2050 = 32'sh0000007e;
	assign w_sys_tmp2067 = (w_sys_tmp2068 + r_run_k_29);
	assign w_sys_tmp2068 = 32'sh00000093;
	assign w_sys_tmp2073 = (w_sys_tmp2074 + r_run_k_29);
	assign w_sys_tmp2074 = 32'sh000000a8;
	assign w_sys_tmp2079 = (w_sys_tmp2080 + r_run_k_29);
	assign w_sys_tmp2080 = 32'sh000000bd;
	assign w_sys_tmp2085 = (w_sys_tmp2086 + r_run_k_29);
	assign w_sys_tmp2086 = 32'sh000000d2;
	assign w_sys_tmp2103 = (w_sys_tmp2104 + r_run_k_29);
	assign w_sys_tmp2104 = 32'sh000000e7;
	assign w_sys_tmp2109 = (w_sys_tmp2110 + r_run_k_29);
	assign w_sys_tmp2110 = 32'sh000000fc;
	assign w_sys_tmp2115 = (w_sys_tmp2116 + r_run_k_29);
	assign w_sys_tmp2116 = 32'sh00000111;
	assign w_sys_tmp2121 = (w_sys_tmp2122 + r_run_k_29);
	assign w_sys_tmp2122 = 32'sh00000126;
	assign w_sys_tmp2139 = (w_sys_tmp2140 + r_run_k_29);
	assign w_sys_tmp2140 = 32'sh0000013b;
	assign w_sys_tmp2145 = (w_sys_tmp2146 + r_run_k_29);
	assign w_sys_tmp2146 = 32'sh00000150;
	assign w_sys_tmp2151 = (w_sys_tmp2152 + r_run_k_29);
	assign w_sys_tmp2152 = 32'sh00000165;
	assign w_sys_tmp2163 = (w_sys_tmp2164 + r_run_k_29);
	assign w_sys_tmp2164 = 32'sh0000017a;
	assign w_sys_tmp2169 = (w_sys_tmp2170 + r_run_k_29);
	assign w_sys_tmp2170 = 32'sh0000018f;
	assign w_sys_tmp2175 = (w_sys_tmp2176 + r_run_k_29);
	assign w_sys_tmp2176 = 32'sh000001a4;
	assign w_sys_tmp2181 = (w_sys_tmp2182 + r_run_k_29);
	assign w_sys_tmp2182 = 32'sh00000019;
	assign w_sys_tmp2187 = (w_sys_tmp2188 + r_run_k_29);
	assign w_sys_tmp2188 = 32'sh0000002e;
	assign w_sys_tmp2193 = (w_sys_tmp2194 + r_run_k_29);
	assign w_sys_tmp2194 = 32'sh00000043;
	assign w_sys_tmp2199 = (w_sys_tmp2200 + r_run_k_29);
	assign w_sys_tmp2200 = 32'sh00000058;
	assign w_sys_tmp2205 = (w_sys_tmp2206 + r_run_k_29);
	assign w_sys_tmp2206 = 32'sh0000006d;
	assign w_sys_tmp2211 = (w_sys_tmp2212 + r_run_k_29);
	assign w_sys_tmp2212 = 32'sh00000082;
	assign w_sys_tmp2229 = (w_sys_tmp2230 + r_run_k_29);
	assign w_sys_tmp2230 = 32'sh00000097;
	assign w_sys_tmp2235 = (w_sys_tmp2236 + r_run_k_29);
	assign w_sys_tmp2236 = 32'sh000000ac;
	assign w_sys_tmp2241 = (w_sys_tmp2242 + r_run_k_29);
	assign w_sys_tmp2242 = 32'sh000000c1;
	assign w_sys_tmp2247 = (w_sys_tmp2248 + r_run_k_29);
	assign w_sys_tmp2248 = 32'sh000000d6;
	assign w_sys_tmp2265 = (w_sys_tmp2266 + r_run_k_29);
	assign w_sys_tmp2266 = 32'sh000000eb;
	assign w_sys_tmp2271 = (w_sys_tmp2272 + r_run_k_29);
	assign w_sys_tmp2272 = 32'sh00000100;
	assign w_sys_tmp2277 = (w_sys_tmp2278 + r_run_k_29);
	assign w_sys_tmp2278 = 32'sh00000115;
	assign w_sys_tmp2283 = (w_sys_tmp2284 + r_run_k_29);
	assign w_sys_tmp2284 = 32'sh0000012a;
	assign w_sys_tmp2301 = (w_sys_tmp2302 + r_run_k_29);
	assign w_sys_tmp2302 = 32'sh0000013f;
	assign w_sys_tmp2307 = (w_sys_tmp2308 + r_run_k_29);
	assign w_sys_tmp2308 = 32'sh00000154;
	assign w_sys_tmp2313 = (w_sys_tmp2314 + r_run_k_29);
	assign w_sys_tmp2314 = 32'sh00000169;
	assign w_sys_tmp2325 = (w_sys_tmp2326 + r_run_k_29);
	assign w_sys_tmp2326 = 32'sh0000017e;
	assign w_sys_tmp2331 = (w_sys_tmp2332 + r_run_k_29);
	assign w_sys_tmp2332 = 32'sh00000193;
	assign w_sys_tmp2337 = (w_sys_tmp2338 + r_run_k_29);
	assign w_sys_tmp2338 = 32'sh000001a8;
	assign w_sys_tmp2343 = (w_sys_tmp2344 + r_run_k_29);
	assign w_sys_tmp2344 = 32'sh0000001d;
	assign w_sys_tmp2349 = (w_sys_tmp2350 + r_run_k_29);
	assign w_sys_tmp2350 = 32'sh00000032;
	assign w_sys_tmp2355 = (w_sys_tmp2356 + r_run_k_29);
	assign w_sys_tmp2356 = 32'sh00000047;
	assign w_sys_tmp2361 = (w_sys_tmp2362 + r_run_k_29);
	assign w_sys_tmp2362 = 32'sh0000005c;
	assign w_sys_tmp2367 = (w_sys_tmp2368 + r_run_k_29);
	assign w_sys_tmp2368 = 32'sh00000071;
	assign w_sys_tmp2373 = (w_sys_tmp2374 + r_run_k_29);
	assign w_sys_tmp2374 = 32'sh00000086;
	assign w_sys_tmp2391 = (w_sys_tmp2392 + r_run_k_29);
	assign w_sys_tmp2392 = 32'sh0000009b;
	assign w_sys_tmp2397 = (w_sys_tmp2398 + r_run_k_29);
	assign w_sys_tmp2398 = 32'sh000000b0;
	assign w_sys_tmp2403 = (w_sys_tmp2404 + r_run_k_29);
	assign w_sys_tmp2404 = 32'sh000000c5;
	assign w_sys_tmp2409 = (w_sys_tmp2410 + r_run_k_29);
	assign w_sys_tmp2410 = 32'sh000000da;
	assign w_sys_tmp2427 = (w_sys_tmp2428 + r_run_k_29);
	assign w_sys_tmp2428 = 32'sh000000ef;
	assign w_sys_tmp2433 = (w_sys_tmp2434 + r_run_k_29);
	assign w_sys_tmp2434 = 32'sh00000104;
	assign w_sys_tmp2439 = (w_sys_tmp2440 + r_run_k_29);
	assign w_sys_tmp2440 = 32'sh00000119;
	assign w_sys_tmp2445 = (w_sys_tmp2446 + r_run_k_29);
	assign w_sys_tmp2446 = 32'sh0000012e;
	assign w_sys_tmp2463 = (w_sys_tmp2464 + r_run_k_29);
	assign w_sys_tmp2464 = 32'sh00000143;
	assign w_sys_tmp2469 = (w_sys_tmp2470 + r_run_k_29);
	assign w_sys_tmp2470 = 32'sh00000158;
	assign w_sys_tmp2475 = (w_sys_tmp2476 + r_run_k_29);
	assign w_sys_tmp2476 = 32'sh0000016d;
	assign w_sys_tmp2487 = (w_sys_tmp2488 + r_run_k_29);
	assign w_sys_tmp2488 = 32'sh00000182;
	assign w_sys_tmp2493 = (w_sys_tmp2494 + r_run_k_29);
	assign w_sys_tmp2494 = 32'sh00000197;
	assign w_sys_tmp2499 = (w_sys_tmp2500 + r_run_k_29);
	assign w_sys_tmp2500 = 32'sh000001ac;
	assign w_sys_tmp2505 = (w_sys_tmp2506 + r_run_k_29);
	assign w_sys_tmp2506 = 32'sh00000021;
	assign w_sys_tmp2511 = (w_sys_tmp2512 + r_run_k_29);
	assign w_sys_tmp2512 = 32'sh00000036;
	assign w_sys_tmp2517 = (w_sys_tmp2518 + r_run_k_29);
	assign w_sys_tmp2518 = 32'sh0000004b;
	assign w_sys_tmp2523 = (w_sys_tmp2524 + r_run_k_29);
	assign w_sys_tmp2524 = 32'sh00000060;
	assign w_sys_tmp2529 = (w_sys_tmp2530 + r_run_k_29);
	assign w_sys_tmp2530 = 32'sh00000075;
	assign w_sys_tmp2535 = (w_sys_tmp2536 + r_run_k_29);
	assign w_sys_tmp2536 = 32'sh0000008a;
	assign w_sys_tmp2553 = (w_sys_tmp2554 + r_run_k_29);
	assign w_sys_tmp2554 = 32'sh0000009f;
	assign w_sys_tmp2559 = (w_sys_tmp2560 + r_run_k_29);
	assign w_sys_tmp2560 = 32'sh000000b4;
	assign w_sys_tmp2565 = (w_sys_tmp2566 + r_run_k_29);
	assign w_sys_tmp2566 = 32'sh000000c9;
	assign w_sys_tmp2571 = (w_sys_tmp2572 + r_run_k_29);
	assign w_sys_tmp2572 = 32'sh000000de;
	assign w_sys_tmp2589 = (w_sys_tmp2590 + r_run_k_29);
	assign w_sys_tmp2590 = 32'sh000000f3;
	assign w_sys_tmp2595 = (w_sys_tmp2596 + r_run_k_29);
	assign w_sys_tmp2596 = 32'sh00000108;
	assign w_sys_tmp2601 = (w_sys_tmp2602 + r_run_k_29);
	assign w_sys_tmp2602 = 32'sh0000011d;
	assign w_sys_tmp2607 = (w_sys_tmp2608 + r_run_k_29);
	assign w_sys_tmp2608 = 32'sh00000132;
	assign w_sys_tmp2625 = (w_sys_tmp2626 + r_run_k_29);
	assign w_sys_tmp2626 = 32'sh00000147;
	assign w_sys_tmp2631 = (w_sys_tmp2632 + r_run_k_29);
	assign w_sys_tmp2632 = 32'sh0000015c;
	assign w_sys_tmp2637 = (w_sys_tmp2638 + r_run_k_29);
	assign w_sys_tmp2638 = 32'sh00000171;
	assign w_sys_tmp2649 = (w_sys_tmp2650 + r_run_k_29);
	assign w_sys_tmp2650 = 32'sh00000186;
	assign w_sys_tmp2655 = (w_sys_tmp2656 + r_run_k_29);
	assign w_sys_tmp2656 = 32'sh0000019b;
	assign w_sys_tmp2661 = (w_sys_tmp2662 + r_run_k_29);
	assign w_sys_tmp2662 = 32'sh000001b0;
	assign w_sys_tmp2666 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp2667 = 32'sh00000011;
	assign w_sys_tmp2668 = ( !w_sys_tmp2669 );
	assign w_sys_tmp2669 = (w_sys_tmp2670 < r_run_k_29);
	assign w_sys_tmp2670 = 32'sh00000015;
	assign w_sys_tmp2673 = (w_sys_tmp2674 + r_run_k_29);
	assign w_sys_tmp2674 = 32'sh00000015;
	assign w_sys_tmp2675 = w_fld_T_0_dataout_1;
	assign w_sys_tmp2679 = (w_sys_tmp2680 + r_run_k_29);
	assign w_sys_tmp2680 = 32'sh0000002a;
	assign w_sys_tmp2685 = (w_sys_tmp2686 + r_run_k_29);
	assign w_sys_tmp2686 = 32'sh0000003f;
	assign w_sys_tmp2691 = (w_sys_tmp2692 + r_run_k_29);
	assign w_sys_tmp2692 = 32'sh00000054;
	assign w_sys_tmp2697 = (w_sys_tmp2698 + r_run_k_29);
	assign w_sys_tmp2698 = 32'sh00000069;
	assign w_sys_tmp2703 = (w_sys_tmp2704 + r_run_k_29);
	assign w_sys_tmp2704 = 32'sh0000007e;
	assign w_sys_tmp2721 = (w_sys_tmp2722 + r_run_k_29);
	assign w_sys_tmp2722 = 32'sh00000093;
	assign w_sys_tmp2727 = (w_sys_tmp2728 + r_run_k_29);
	assign w_sys_tmp2728 = 32'sh000000a8;
	assign w_sys_tmp2733 = (w_sys_tmp2734 + r_run_k_29);
	assign w_sys_tmp2734 = 32'sh000000bd;
	assign w_sys_tmp2739 = (w_sys_tmp2740 + r_run_k_29);
	assign w_sys_tmp2740 = 32'sh000000d2;
	assign w_sys_tmp2757 = (w_sys_tmp2758 + r_run_k_29);
	assign w_sys_tmp2758 = 32'sh000000e7;
	assign w_sys_tmp2763 = (w_sys_tmp2764 + r_run_k_29);
	assign w_sys_tmp2764 = 32'sh000000fc;
	assign w_sys_tmp2769 = (w_sys_tmp2770 + r_run_k_29);
	assign w_sys_tmp2770 = 32'sh00000111;
	assign w_sys_tmp2775 = (w_sys_tmp2776 + r_run_k_29);
	assign w_sys_tmp2776 = 32'sh00000126;
	assign w_sys_tmp2793 = (w_sys_tmp2794 + r_run_k_29);
	assign w_sys_tmp2794 = 32'sh0000013b;
	assign w_sys_tmp2799 = (w_sys_tmp2800 + r_run_k_29);
	assign w_sys_tmp2800 = 32'sh00000150;
	assign w_sys_tmp2805 = (w_sys_tmp2806 + r_run_k_29);
	assign w_sys_tmp2806 = 32'sh00000165;
	assign w_sys_tmp2817 = (w_sys_tmp2818 + r_run_k_29);
	assign w_sys_tmp2818 = 32'sh0000017a;
	assign w_sys_tmp2823 = (w_sys_tmp2824 + r_run_k_29);
	assign w_sys_tmp2824 = 32'sh0000018f;
	assign w_sys_tmp2829 = (w_sys_tmp2830 + r_run_k_29);
	assign w_sys_tmp2830 = 32'sh000001a4;
	assign w_sys_tmp2834 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp2835 = 32'sh00000002;
	assign w_sys_tmp2836 = ( !w_sys_tmp2837 );
	assign w_sys_tmp2837 = (w_sys_tmp2838 < r_run_k_29);
	assign w_sys_tmp2838 = 32'sh00000005;
	assign w_sys_tmp2841 = (w_sys_tmp2842 + r_run_k_29);
	assign w_sys_tmp2842 = 32'sh0000002a;
	assign w_sys_tmp2843 = w_sub00_result_dataout;
	assign w_sys_tmp2847 = (w_sys_tmp2848 + r_run_k_29);
	assign w_sys_tmp2848 = 32'sh0000003f;
	assign w_sys_tmp2853 = (w_sys_tmp2854 + r_run_k_29);
	assign w_sys_tmp2854 = 32'sh00000054;
	assign w_sys_tmp2859 = (w_sys_tmp2860 + r_run_k_29);
	assign w_sys_tmp2860 = 32'sh00000069;
	assign w_sys_tmp2865 = (w_sys_tmp2866 + r_run_k_29);
	assign w_sys_tmp2866 = 32'sh0000007e;
	assign w_sys_tmp2870 = (w_sys_tmp2871 + r_run_k_29);
	assign w_sys_tmp2871 = 32'sh00000093;
	assign w_sys_tmp2875 = (w_sys_tmp2876 + r_run_k_29);
	assign w_sys_tmp2876 = 32'sh000000a8;
	assign w_sys_tmp2880 = (w_sys_tmp2881 + r_run_k_29);
	assign w_sys_tmp2881 = 32'sh000000bd;
	assign w_sys_tmp2885 = (w_sys_tmp2886 + r_run_k_29);
	assign w_sys_tmp2886 = 32'sh000000d2;
	assign w_sys_tmp2890 = (w_sys_tmp2891 + r_run_k_29);
	assign w_sys_tmp2891 = 32'sh000000e7;
	assign w_sys_tmp2895 = (w_sys_tmp2896 + r_run_k_29);
	assign w_sys_tmp2896 = 32'sh000000fc;
	assign w_sys_tmp2900 = (w_sys_tmp2901 + r_run_k_29);
	assign w_sys_tmp2901 = 32'sh00000111;
	assign w_sys_tmp2905 = (w_sys_tmp2906 + r_run_k_29);
	assign w_sys_tmp2906 = 32'sh00000126;
	assign w_sys_tmp2910 = (w_sys_tmp2911 + r_run_k_29);
	assign w_sys_tmp2911 = 32'sh0000013b;
	assign w_sys_tmp2915 = (w_sys_tmp2916 + r_run_k_29);
	assign w_sys_tmp2916 = 32'sh00000150;
	assign w_sys_tmp2920 = (w_sys_tmp2921 + r_run_k_29);
	assign w_sys_tmp2921 = 32'sh00000165;
	assign w_sys_tmp2925 = (w_sys_tmp2926 + r_run_k_29);
	assign w_sys_tmp2926 = 32'sh0000017a;
	assign w_sys_tmp2930 = (w_sys_tmp2931 + r_run_k_29);
	assign w_sys_tmp2931 = 32'sh0000018f;
	assign w_sys_tmp2935 = (w_sys_tmp2936 + r_run_k_29);
	assign w_sys_tmp2936 = 32'sh000001a4;
	assign w_sys_tmp2940 = (w_sys_tmp2941 + r_run_k_29);
	assign w_sys_tmp2941 = 32'sh0000002e;
	assign w_sys_tmp2945 = (w_sys_tmp2946 + r_run_k_29);
	assign w_sys_tmp2946 = 32'sh00000043;
	assign w_sys_tmp2950 = (w_sys_tmp2951 + r_run_k_29);
	assign w_sys_tmp2951 = 32'sh00000058;
	assign w_sys_tmp2955 = (w_sys_tmp2956 + r_run_k_29);
	assign w_sys_tmp2956 = 32'sh0000006d;
	assign w_sys_tmp2960 = (w_sys_tmp2961 + r_run_k_29);
	assign w_sys_tmp2961 = 32'sh00000082;
	assign w_sys_tmp2965 = (w_sys_tmp2966 + r_run_k_29);
	assign w_sys_tmp2966 = 32'sh00000097;
	assign w_sys_tmp2970 = (w_sys_tmp2971 + r_run_k_29);
	assign w_sys_tmp2971 = 32'sh000000ac;
	assign w_sys_tmp2975 = (w_sys_tmp2976 + r_run_k_29);
	assign w_sys_tmp2976 = 32'sh000000c1;
	assign w_sys_tmp2980 = (w_sys_tmp2981 + r_run_k_29);
	assign w_sys_tmp2981 = 32'sh000000d6;
	assign w_sys_tmp2985 = (w_sys_tmp2986 + r_run_k_29);
	assign w_sys_tmp2986 = 32'sh000000eb;
	assign w_sys_tmp2990 = (w_sys_tmp2991 + r_run_k_29);
	assign w_sys_tmp2991 = 32'sh00000100;
	assign w_sys_tmp2995 = (w_sys_tmp2996 + r_run_k_29);
	assign w_sys_tmp2996 = 32'sh00000115;
	assign w_sys_tmp3000 = (w_sys_tmp3001 + r_run_k_29);
	assign w_sys_tmp3001 = 32'sh0000012a;
	assign w_sys_tmp3005 = (w_sys_tmp3006 + r_run_k_29);
	assign w_sys_tmp3006 = 32'sh0000013f;
	assign w_sys_tmp3010 = (w_sys_tmp3011 + r_run_k_29);
	assign w_sys_tmp3011 = 32'sh00000154;
	assign w_sys_tmp3015 = (w_sys_tmp3016 + r_run_k_29);
	assign w_sys_tmp3016 = 32'sh00000169;
	assign w_sys_tmp3020 = (w_sys_tmp3021 + r_run_k_29);
	assign w_sys_tmp3021 = 32'sh0000017e;
	assign w_sys_tmp3025 = (w_sys_tmp3026 + r_run_k_29);
	assign w_sys_tmp3026 = 32'sh00000193;
	assign w_sys_tmp3030 = (w_sys_tmp3031 + r_run_k_29);
	assign w_sys_tmp3031 = 32'sh000001a8;
	assign w_sys_tmp3035 = (w_sys_tmp3036 + r_run_k_29);
	assign w_sys_tmp3036 = 32'sh00000032;
	assign w_sys_tmp3040 = (w_sys_tmp3041 + r_run_k_29);
	assign w_sys_tmp3041 = 32'sh00000047;
	assign w_sys_tmp3045 = (w_sys_tmp3046 + r_run_k_29);
	assign w_sys_tmp3046 = 32'sh0000005c;
	assign w_sys_tmp3050 = (w_sys_tmp3051 + r_run_k_29);
	assign w_sys_tmp3051 = 32'sh00000071;
	assign w_sys_tmp3055 = (w_sys_tmp3056 + r_run_k_29);
	assign w_sys_tmp3056 = 32'sh00000086;
	assign w_sys_tmp3060 = (w_sys_tmp3061 + r_run_k_29);
	assign w_sys_tmp3061 = 32'sh0000009b;
	assign w_sys_tmp3065 = (w_sys_tmp3066 + r_run_k_29);
	assign w_sys_tmp3066 = 32'sh000000b0;
	assign w_sys_tmp3070 = (w_sys_tmp3071 + r_run_k_29);
	assign w_sys_tmp3071 = 32'sh000000c5;
	assign w_sys_tmp3075 = (w_sys_tmp3076 + r_run_k_29);
	assign w_sys_tmp3076 = 32'sh000000da;
	assign w_sys_tmp3080 = (w_sys_tmp3081 + r_run_k_29);
	assign w_sys_tmp3081 = 32'sh000000ef;
	assign w_sys_tmp3085 = (w_sys_tmp3086 + r_run_k_29);
	assign w_sys_tmp3086 = 32'sh00000104;
	assign w_sys_tmp3090 = (w_sys_tmp3091 + r_run_k_29);
	assign w_sys_tmp3091 = 32'sh00000119;
	assign w_sys_tmp3095 = (w_sys_tmp3096 + r_run_k_29);
	assign w_sys_tmp3096 = 32'sh0000012e;
	assign w_sys_tmp3100 = (w_sys_tmp3101 + r_run_k_29);
	assign w_sys_tmp3101 = 32'sh00000143;
	assign w_sys_tmp3105 = (w_sys_tmp3106 + r_run_k_29);
	assign w_sys_tmp3106 = 32'sh00000158;
	assign w_sys_tmp3110 = (w_sys_tmp3111 + r_run_k_29);
	assign w_sys_tmp3111 = 32'sh0000016d;
	assign w_sys_tmp3115 = (w_sys_tmp3116 + r_run_k_29);
	assign w_sys_tmp3116 = 32'sh00000182;
	assign w_sys_tmp3120 = (w_sys_tmp3121 + r_run_k_29);
	assign w_sys_tmp3121 = 32'sh00000197;
	assign w_sys_tmp3125 = (w_sys_tmp3126 + r_run_k_29);
	assign w_sys_tmp3126 = 32'sh000001ac;
	assign w_sys_tmp3130 = (w_sys_tmp3131 + r_run_k_29);
	assign w_sys_tmp3131 = 32'sh00000036;
	assign w_sys_tmp3135 = (w_sys_tmp3136 + r_run_k_29);
	assign w_sys_tmp3136 = 32'sh0000004b;
	assign w_sys_tmp3140 = (w_sys_tmp3141 + r_run_k_29);
	assign w_sys_tmp3141 = 32'sh00000060;
	assign w_sys_tmp3145 = (w_sys_tmp3146 + r_run_k_29);
	assign w_sys_tmp3146 = 32'sh00000075;
	assign w_sys_tmp3150 = (w_sys_tmp3151 + r_run_k_29);
	assign w_sys_tmp3151 = 32'sh0000008a;
	assign w_sys_tmp3155 = (w_sys_tmp3156 + r_run_k_29);
	assign w_sys_tmp3156 = 32'sh0000009f;
	assign w_sys_tmp3160 = (w_sys_tmp3161 + r_run_k_29);
	assign w_sys_tmp3161 = 32'sh000000b4;
	assign w_sys_tmp3165 = (w_sys_tmp3166 + r_run_k_29);
	assign w_sys_tmp3166 = 32'sh000000c9;
	assign w_sys_tmp3170 = (w_sys_tmp3171 + r_run_k_29);
	assign w_sys_tmp3171 = 32'sh000000de;
	assign w_sys_tmp3175 = (w_sys_tmp3176 + r_run_k_29);
	assign w_sys_tmp3176 = 32'sh000000f3;
	assign w_sys_tmp3180 = (w_sys_tmp3181 + r_run_k_29);
	assign w_sys_tmp3181 = 32'sh00000108;
	assign w_sys_tmp3185 = (w_sys_tmp3186 + r_run_k_29);
	assign w_sys_tmp3186 = 32'sh0000011d;
	assign w_sys_tmp3190 = (w_sys_tmp3191 + r_run_k_29);
	assign w_sys_tmp3191 = 32'sh00000132;
	assign w_sys_tmp3195 = (w_sys_tmp3196 + r_run_k_29);
	assign w_sys_tmp3196 = 32'sh00000147;
	assign w_sys_tmp3200 = (w_sys_tmp3201 + r_run_k_29);
	assign w_sys_tmp3201 = 32'sh0000015c;
	assign w_sys_tmp3205 = (w_sys_tmp3206 + r_run_k_29);
	assign w_sys_tmp3206 = 32'sh00000171;
	assign w_sys_tmp3210 = (w_sys_tmp3211 + r_run_k_29);
	assign w_sys_tmp3211 = 32'sh00000186;
	assign w_sys_tmp3215 = (w_sys_tmp3216 + r_run_k_29);
	assign w_sys_tmp3216 = 32'sh0000019b;
	assign w_sys_tmp3220 = (w_sys_tmp3221 + r_run_k_29);
	assign w_sys_tmp3221 = 32'sh000001b0;
	assign w_sys_tmp3224 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp3225 = 32'sh00000012;
	assign w_sys_tmp3226 = ( !w_sys_tmp3227 );
	assign w_sys_tmp3227 = (w_sys_tmp3228 < r_run_k_29);
	assign w_sys_tmp3228 = 32'sh00000014;
	assign w_sys_tmp3231 = (w_sys_tmp3232 + r_run_k_29);
	assign w_sys_tmp3232 = 32'sh0000002a;
	assign w_sys_tmp3233 = w_sub20_result_dataout;
	assign w_sys_tmp3237 = (w_sys_tmp3238 + r_run_k_29);
	assign w_sys_tmp3238 = 32'sh0000003f;
	assign w_sys_tmp3243 = (w_sys_tmp3244 + r_run_k_29);
	assign w_sys_tmp3244 = 32'sh00000054;
	assign w_sys_tmp3249 = (w_sys_tmp3250 + r_run_k_29);
	assign w_sys_tmp3250 = 32'sh00000069;
	assign w_sys_tmp3255 = (w_sys_tmp3256 + r_run_k_29);
	assign w_sys_tmp3256 = 32'sh0000007e;
	assign w_sys_tmp3260 = (w_sys_tmp3261 + r_run_k_29);
	assign w_sys_tmp3261 = 32'sh00000093;
	assign w_sys_tmp3265 = (w_sys_tmp3266 + r_run_k_29);
	assign w_sys_tmp3266 = 32'sh000000a8;
	assign w_sys_tmp3270 = (w_sys_tmp3271 + r_run_k_29);
	assign w_sys_tmp3271 = 32'sh000000bd;
	assign w_sys_tmp3275 = (w_sys_tmp3276 + r_run_k_29);
	assign w_sys_tmp3276 = 32'sh000000d2;
	assign w_sys_tmp3280 = (w_sys_tmp3281 + r_run_k_29);
	assign w_sys_tmp3281 = 32'sh000000e7;
	assign w_sys_tmp3285 = (w_sys_tmp3286 + r_run_k_29);
	assign w_sys_tmp3286 = 32'sh000000fc;
	assign w_sys_tmp3290 = (w_sys_tmp3291 + r_run_k_29);
	assign w_sys_tmp3291 = 32'sh00000111;
	assign w_sys_tmp3295 = (w_sys_tmp3296 + r_run_k_29);
	assign w_sys_tmp3296 = 32'sh00000126;
	assign w_sys_tmp3300 = (w_sys_tmp3301 + r_run_k_29);
	assign w_sys_tmp3301 = 32'sh0000013b;
	assign w_sys_tmp3305 = (w_sys_tmp3306 + r_run_k_29);
	assign w_sys_tmp3306 = 32'sh00000150;
	assign w_sys_tmp3310 = (w_sys_tmp3311 + r_run_k_29);
	assign w_sys_tmp3311 = 32'sh00000165;
	assign w_sys_tmp3315 = (w_sys_tmp3316 + r_run_k_29);
	assign w_sys_tmp3316 = 32'sh0000017a;
	assign w_sys_tmp3320 = (w_sys_tmp3321 + r_run_k_29);
	assign w_sys_tmp3321 = 32'sh0000018f;
	assign w_sys_tmp3325 = (w_sys_tmp3326 + r_run_k_29);
	assign w_sys_tmp3326 = 32'sh000001a4;
	assign w_sys_tmp3329 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp3330 = w_fld_T_0_dataout_1;
	assign w_sys_tmp3331 = 32'sh000000dc;


	sub19
		sub19_inst(
			.i_fld_T_0_addr_0 (w_sub19_T_addr),
			.i_fld_T_0_datain_0 (w_sub19_T_datain),
			.o_fld_T_0_dataout_0 (w_sub19_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub19_T_r_w),
			.i_fld_U_2_addr_0 (w_sub19_U_addr),
			.i_fld_U_2_datain_0 (w_sub19_U_datain),
			.o_fld_U_2_dataout_0 (w_sub19_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub19_U_r_w),
			.i_fld_V_1_addr_0 (w_sub19_V_addr),
			.i_fld_V_1_datain_0 (w_sub19_V_datain),
			.o_fld_V_1_dataout_0 (w_sub19_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub19_V_r_w),
			.i_fld_result_3_addr_0 (w_sub19_result_addr),
			.i_fld_result_3_datain_0 (w_sub19_result_datain),
			.o_fld_result_3_dataout_0 (w_sub19_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub19_result_r_w),
			.o_run_busy (w_sub19_run_busy),
			.i_run_req (r_sub19_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub09
		sub09_inst(
			.i_fld_T_0_addr_0 (w_sub09_T_addr),
			.i_fld_T_0_datain_0 (w_sub09_T_datain),
			.o_fld_T_0_dataout_0 (w_sub09_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub09_T_r_w),
			.i_fld_U_2_addr_0 (w_sub09_U_addr),
			.i_fld_U_2_datain_0 (w_sub09_U_datain),
			.o_fld_U_2_dataout_0 (w_sub09_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub09_U_r_w),
			.i_fld_V_1_addr_0 (w_sub09_V_addr),
			.i_fld_V_1_datain_0 (w_sub09_V_datain),
			.o_fld_V_1_dataout_0 (w_sub09_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub09_V_r_w),
			.i_fld_result_3_addr_0 (w_sub09_result_addr),
			.i_fld_result_3_datain_0 (w_sub09_result_datain),
			.o_fld_result_3_dataout_0 (w_sub09_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub09_result_r_w),
			.o_run_busy (w_sub09_run_busy),
			.i_run_req (r_sub09_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub08
		sub08_inst(
			.i_fld_T_0_addr_0 (w_sub08_T_addr),
			.i_fld_T_0_datain_0 (w_sub08_T_datain),
			.o_fld_T_0_dataout_0 (w_sub08_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub08_T_r_w),
			.i_fld_U_2_addr_0 (w_sub08_U_addr),
			.i_fld_U_2_datain_0 (w_sub08_U_datain),
			.o_fld_U_2_dataout_0 (w_sub08_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub08_U_r_w),
			.i_fld_V_1_addr_0 (w_sub08_V_addr),
			.i_fld_V_1_datain_0 (w_sub08_V_datain),
			.o_fld_V_1_dataout_0 (w_sub08_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub08_V_r_w),
			.i_fld_result_3_addr_0 (w_sub08_result_addr),
			.i_fld_result_3_datain_0 (w_sub08_result_datain),
			.o_fld_result_3_dataout_0 (w_sub08_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub08_result_r_w),
			.o_run_busy (w_sub08_run_busy),
			.i_run_req (r_sub08_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub24
		sub24_inst(
			.i_fld_T_0_addr_0 (w_sub24_T_addr),
			.i_fld_T_0_datain_0 (w_sub24_T_datain),
			.o_fld_T_0_dataout_0 (w_sub24_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub24_T_r_w),
			.i_fld_U_2_addr_0 (w_sub24_U_addr),
			.i_fld_U_2_datain_0 (w_sub24_U_datain),
			.o_fld_U_2_dataout_0 (w_sub24_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub24_U_r_w),
			.i_fld_V_1_addr_0 (w_sub24_V_addr),
			.i_fld_V_1_datain_0 (w_sub24_V_datain),
			.o_fld_V_1_dataout_0 (w_sub24_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub24_V_r_w),
			.i_fld_result_3_addr_0 (w_sub24_result_addr),
			.i_fld_result_3_datain_0 (w_sub24_result_datain),
			.o_fld_result_3_dataout_0 (w_sub24_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub24_result_r_w),
			.o_run_busy (w_sub24_run_busy),
			.i_run_req (r_sub24_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub22
		sub22_inst(
			.i_fld_T_0_addr_0 (w_sub22_T_addr),
			.i_fld_T_0_datain_0 (w_sub22_T_datain),
			.o_fld_T_0_dataout_0 (w_sub22_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub22_T_r_w),
			.i_fld_U_2_addr_0 (w_sub22_U_addr),
			.i_fld_U_2_datain_0 (w_sub22_U_datain),
			.o_fld_U_2_dataout_0 (w_sub22_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub22_U_r_w),
			.i_fld_V_1_addr_0 (w_sub22_V_addr),
			.i_fld_V_1_datain_0 (w_sub22_V_datain),
			.o_fld_V_1_dataout_0 (w_sub22_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub22_V_r_w),
			.i_fld_result_3_addr_0 (w_sub22_result_addr),
			.i_fld_result_3_datain_0 (w_sub22_result_datain),
			.o_fld_result_3_dataout_0 (w_sub22_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub22_result_r_w),
			.o_run_busy (w_sub22_run_busy),
			.i_run_req (r_sub22_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub23
		sub23_inst(
			.i_fld_T_0_addr_0 (w_sub23_T_addr),
			.i_fld_T_0_datain_0 (w_sub23_T_datain),
			.o_fld_T_0_dataout_0 (w_sub23_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub23_T_r_w),
			.i_fld_U_2_addr_0 (w_sub23_U_addr),
			.i_fld_U_2_datain_0 (w_sub23_U_datain),
			.o_fld_U_2_dataout_0 (w_sub23_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub23_U_r_w),
			.i_fld_V_1_addr_0 (w_sub23_V_addr),
			.i_fld_V_1_datain_0 (w_sub23_V_datain),
			.o_fld_V_1_dataout_0 (w_sub23_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub23_V_r_w),
			.i_fld_result_3_addr_0 (w_sub23_result_addr),
			.i_fld_result_3_datain_0 (w_sub23_result_datain),
			.o_fld_result_3_dataout_0 (w_sub23_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub23_result_r_w),
			.o_run_busy (w_sub23_run_busy),
			.i_run_req (r_sub23_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub12
		sub12_inst(
			.i_fld_T_0_addr_0 (w_sub12_T_addr),
			.i_fld_T_0_datain_0 (w_sub12_T_datain),
			.o_fld_T_0_dataout_0 (w_sub12_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub12_T_r_w),
			.i_fld_U_2_addr_0 (w_sub12_U_addr),
			.i_fld_U_2_datain_0 (w_sub12_U_datain),
			.o_fld_U_2_dataout_0 (w_sub12_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub12_U_r_w),
			.i_fld_V_1_addr_0 (w_sub12_V_addr),
			.i_fld_V_1_datain_0 (w_sub12_V_datain),
			.o_fld_V_1_dataout_0 (w_sub12_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub12_V_r_w),
			.i_fld_result_3_addr_0 (w_sub12_result_addr),
			.i_fld_result_3_datain_0 (w_sub12_result_datain),
			.o_fld_result_3_dataout_0 (w_sub12_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub12_result_r_w),
			.o_run_busy (w_sub12_run_busy),
			.i_run_req (r_sub12_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub03
		sub03_inst(
			.i_fld_T_0_addr_0 (w_sub03_T_addr),
			.i_fld_T_0_datain_0 (w_sub03_T_datain),
			.o_fld_T_0_dataout_0 (w_sub03_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub03_T_r_w),
			.i_fld_U_2_addr_0 (w_sub03_U_addr),
			.i_fld_U_2_datain_0 (w_sub03_U_datain),
			.o_fld_U_2_dataout_0 (w_sub03_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub03_U_r_w),
			.i_fld_V_1_addr_0 (w_sub03_V_addr),
			.i_fld_V_1_datain_0 (w_sub03_V_datain),
			.o_fld_V_1_dataout_0 (w_sub03_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub03_V_r_w),
			.i_fld_result_3_addr_0 (w_sub03_result_addr),
			.i_fld_result_3_datain_0 (w_sub03_result_datain),
			.o_fld_result_3_dataout_0 (w_sub03_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub03_result_r_w),
			.o_run_busy (w_sub03_run_busy),
			.i_run_req (r_sub03_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub02
		sub02_inst(
			.i_fld_T_0_addr_0 (w_sub02_T_addr),
			.i_fld_T_0_datain_0 (w_sub02_T_datain),
			.o_fld_T_0_dataout_0 (w_sub02_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub02_T_r_w),
			.i_fld_U_2_addr_0 (w_sub02_U_addr),
			.i_fld_U_2_datain_0 (w_sub02_U_datain),
			.o_fld_U_2_dataout_0 (w_sub02_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub02_U_r_w),
			.i_fld_V_1_addr_0 (w_sub02_V_addr),
			.i_fld_V_1_datain_0 (w_sub02_V_datain),
			.o_fld_V_1_dataout_0 (w_sub02_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub02_V_r_w),
			.i_fld_result_3_addr_0 (w_sub02_result_addr),
			.i_fld_result_3_datain_0 (w_sub02_result_datain),
			.o_fld_result_3_dataout_0 (w_sub02_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub02_result_r_w),
			.o_run_busy (w_sub02_run_busy),
			.i_run_req (r_sub02_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub11
		sub11_inst(
			.i_fld_T_0_addr_0 (w_sub11_T_addr),
			.i_fld_T_0_datain_0 (w_sub11_T_datain),
			.o_fld_T_0_dataout_0 (w_sub11_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub11_T_r_w),
			.i_fld_U_2_addr_0 (w_sub11_U_addr),
			.i_fld_U_2_datain_0 (w_sub11_U_datain),
			.o_fld_U_2_dataout_0 (w_sub11_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub11_U_r_w),
			.i_fld_V_1_addr_0 (w_sub11_V_addr),
			.i_fld_V_1_datain_0 (w_sub11_V_datain),
			.o_fld_V_1_dataout_0 (w_sub11_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub11_V_r_w),
			.i_fld_result_3_addr_0 (w_sub11_result_addr),
			.i_fld_result_3_datain_0 (w_sub11_result_datain),
			.o_fld_result_3_dataout_0 (w_sub11_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub11_result_r_w),
			.o_run_busy (w_sub11_run_busy),
			.i_run_req (r_sub11_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub14
		sub14_inst(
			.i_fld_T_0_addr_0 (w_sub14_T_addr),
			.i_fld_T_0_datain_0 (w_sub14_T_datain),
			.o_fld_T_0_dataout_0 (w_sub14_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub14_T_r_w),
			.i_fld_U_2_addr_0 (w_sub14_U_addr),
			.i_fld_U_2_datain_0 (w_sub14_U_datain),
			.o_fld_U_2_dataout_0 (w_sub14_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub14_U_r_w),
			.i_fld_V_1_addr_0 (w_sub14_V_addr),
			.i_fld_V_1_datain_0 (w_sub14_V_datain),
			.o_fld_V_1_dataout_0 (w_sub14_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub14_V_r_w),
			.i_fld_result_3_addr_0 (w_sub14_result_addr),
			.i_fld_result_3_datain_0 (w_sub14_result_datain),
			.o_fld_result_3_dataout_0 (w_sub14_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub14_result_r_w),
			.o_run_busy (w_sub14_run_busy),
			.i_run_req (r_sub14_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub01
		sub01_inst(
			.i_fld_T_0_addr_0 (w_sub01_T_addr),
			.i_fld_T_0_datain_0 (w_sub01_T_datain),
			.o_fld_T_0_dataout_0 (w_sub01_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub01_T_r_w),
			.i_fld_U_2_addr_0 (w_sub01_U_addr),
			.i_fld_U_2_datain_0 (w_sub01_U_datain),
			.o_fld_U_2_dataout_0 (w_sub01_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub01_U_r_w),
			.i_fld_V_1_addr_0 (w_sub01_V_addr),
			.i_fld_V_1_datain_0 (w_sub01_V_datain),
			.o_fld_V_1_dataout_0 (w_sub01_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub01_V_r_w),
			.i_fld_result_3_addr_0 (w_sub01_result_addr),
			.i_fld_result_3_datain_0 (w_sub01_result_datain),
			.o_fld_result_3_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub01_result_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub00
		sub00_inst(
			.i_fld_T_0_addr_0 (w_sub00_T_addr),
			.i_fld_T_0_datain_0 (w_sub00_T_datain),
			.o_fld_T_0_dataout_0 (w_sub00_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub00_T_r_w),
			.i_fld_U_2_addr_0 (w_sub00_U_addr),
			.i_fld_U_2_datain_0 (w_sub00_U_datain),
			.o_fld_U_2_dataout_0 (w_sub00_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub00_U_r_w),
			.i_fld_V_1_addr_0 (w_sub00_V_addr),
			.i_fld_V_1_datain_0 (w_sub00_V_datain),
			.o_fld_V_1_dataout_0 (w_sub00_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub00_V_r_w),
			.i_fld_result_3_addr_0 (w_sub00_result_addr),
			.i_fld_result_3_datain_0 (w_sub00_result_datain),
			.o_fld_result_3_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub00_result_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub13
		sub13_inst(
			.i_fld_T_0_addr_0 (w_sub13_T_addr),
			.i_fld_T_0_datain_0 (w_sub13_T_datain),
			.o_fld_T_0_dataout_0 (w_sub13_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub13_T_r_w),
			.i_fld_U_2_addr_0 (w_sub13_U_addr),
			.i_fld_U_2_datain_0 (w_sub13_U_datain),
			.o_fld_U_2_dataout_0 (w_sub13_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub13_U_r_w),
			.i_fld_V_1_addr_0 (w_sub13_V_addr),
			.i_fld_V_1_datain_0 (w_sub13_V_datain),
			.o_fld_V_1_dataout_0 (w_sub13_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub13_V_r_w),
			.i_fld_result_3_addr_0 (w_sub13_result_addr),
			.i_fld_result_3_datain_0 (w_sub13_result_datain),
			.o_fld_result_3_dataout_0 (w_sub13_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub13_result_r_w),
			.o_run_busy (w_sub13_run_busy),
			.i_run_req (r_sub13_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub07
		sub07_inst(
			.i_fld_T_0_addr_0 (w_sub07_T_addr),
			.i_fld_T_0_datain_0 (w_sub07_T_datain),
			.o_fld_T_0_dataout_0 (w_sub07_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub07_T_r_w),
			.i_fld_U_2_addr_0 (w_sub07_U_addr),
			.i_fld_U_2_datain_0 (w_sub07_U_datain),
			.o_fld_U_2_dataout_0 (w_sub07_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub07_U_r_w),
			.i_fld_V_1_addr_0 (w_sub07_V_addr),
			.i_fld_V_1_datain_0 (w_sub07_V_datain),
			.o_fld_V_1_dataout_0 (w_sub07_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub07_V_r_w),
			.i_fld_result_3_addr_0 (w_sub07_result_addr),
			.i_fld_result_3_datain_0 (w_sub07_result_datain),
			.o_fld_result_3_dataout_0 (w_sub07_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub07_result_r_w),
			.o_run_busy (w_sub07_run_busy),
			.i_run_req (r_sub07_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub16
		sub16_inst(
			.i_fld_T_0_addr_0 (w_sub16_T_addr),
			.i_fld_T_0_datain_0 (w_sub16_T_datain),
			.o_fld_T_0_dataout_0 (w_sub16_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub16_T_r_w),
			.i_fld_U_2_addr_0 (w_sub16_U_addr),
			.i_fld_U_2_datain_0 (w_sub16_U_datain),
			.o_fld_U_2_dataout_0 (w_sub16_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub16_U_r_w),
			.i_fld_V_1_addr_0 (w_sub16_V_addr),
			.i_fld_V_1_datain_0 (w_sub16_V_datain),
			.o_fld_V_1_dataout_0 (w_sub16_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub16_V_r_w),
			.i_fld_result_3_addr_0 (w_sub16_result_addr),
			.i_fld_result_3_datain_0 (w_sub16_result_datain),
			.o_fld_result_3_dataout_0 (w_sub16_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub16_result_r_w),
			.o_run_busy (w_sub16_run_busy),
			.i_run_req (r_sub16_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub06
		sub06_inst(
			.i_fld_T_0_addr_0 (w_sub06_T_addr),
			.i_fld_T_0_datain_0 (w_sub06_T_datain),
			.o_fld_T_0_dataout_0 (w_sub06_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub06_T_r_w),
			.i_fld_U_2_addr_0 (w_sub06_U_addr),
			.i_fld_U_2_datain_0 (w_sub06_U_datain),
			.o_fld_U_2_dataout_0 (w_sub06_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub06_U_r_w),
			.i_fld_V_1_addr_0 (w_sub06_V_addr),
			.i_fld_V_1_datain_0 (w_sub06_V_datain),
			.o_fld_V_1_dataout_0 (w_sub06_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub06_V_r_w),
			.i_fld_result_3_addr_0 (w_sub06_result_addr),
			.i_fld_result_3_datain_0 (w_sub06_result_datain),
			.o_fld_result_3_dataout_0 (w_sub06_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub06_result_r_w),
			.o_run_busy (w_sub06_run_busy),
			.i_run_req (r_sub06_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub15
		sub15_inst(
			.i_fld_T_0_addr_0 (w_sub15_T_addr),
			.i_fld_T_0_datain_0 (w_sub15_T_datain),
			.o_fld_T_0_dataout_0 (w_sub15_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub15_T_r_w),
			.i_fld_U_2_addr_0 (w_sub15_U_addr),
			.i_fld_U_2_datain_0 (w_sub15_U_datain),
			.o_fld_U_2_dataout_0 (w_sub15_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub15_U_r_w),
			.i_fld_V_1_addr_0 (w_sub15_V_addr),
			.i_fld_V_1_datain_0 (w_sub15_V_datain),
			.o_fld_V_1_dataout_0 (w_sub15_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub15_V_r_w),
			.i_fld_result_3_addr_0 (w_sub15_result_addr),
			.i_fld_result_3_datain_0 (w_sub15_result_datain),
			.o_fld_result_3_dataout_0 (w_sub15_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub15_result_r_w),
			.o_run_busy (w_sub15_run_busy),
			.i_run_req (r_sub15_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub05
		sub05_inst(
			.i_fld_T_0_addr_0 (w_sub05_T_addr),
			.i_fld_T_0_datain_0 (w_sub05_T_datain),
			.o_fld_T_0_dataout_0 (w_sub05_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub05_T_r_w),
			.i_fld_U_2_addr_0 (w_sub05_U_addr),
			.i_fld_U_2_datain_0 (w_sub05_U_datain),
			.o_fld_U_2_dataout_0 (w_sub05_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub05_U_r_w),
			.i_fld_V_1_addr_0 (w_sub05_V_addr),
			.i_fld_V_1_datain_0 (w_sub05_V_datain),
			.o_fld_V_1_dataout_0 (w_sub05_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub05_V_r_w),
			.i_fld_result_3_addr_0 (w_sub05_result_addr),
			.i_fld_result_3_datain_0 (w_sub05_result_datain),
			.o_fld_result_3_dataout_0 (w_sub05_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub05_result_r_w),
			.o_run_busy (w_sub05_run_busy),
			.i_run_req (r_sub05_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub18
		sub18_inst(
			.i_fld_T_0_addr_0 (w_sub18_T_addr),
			.i_fld_T_0_datain_0 (w_sub18_T_datain),
			.o_fld_T_0_dataout_0 (w_sub18_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub18_T_r_w),
			.i_fld_U_2_addr_0 (w_sub18_U_addr),
			.i_fld_U_2_datain_0 (w_sub18_U_datain),
			.o_fld_U_2_dataout_0 (w_sub18_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub18_U_r_w),
			.i_fld_V_1_addr_0 (w_sub18_V_addr),
			.i_fld_V_1_datain_0 (w_sub18_V_datain),
			.o_fld_V_1_dataout_0 (w_sub18_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub18_V_r_w),
			.i_fld_result_3_addr_0 (w_sub18_result_addr),
			.i_fld_result_3_datain_0 (w_sub18_result_datain),
			.o_fld_result_3_dataout_0 (w_sub18_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub18_result_r_w),
			.o_run_busy (w_sub18_run_busy),
			.i_run_req (r_sub18_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub04
		sub04_inst(
			.i_fld_T_0_addr_0 (w_sub04_T_addr),
			.i_fld_T_0_datain_0 (w_sub04_T_datain),
			.o_fld_T_0_dataout_0 (w_sub04_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub04_T_r_w),
			.i_fld_U_2_addr_0 (w_sub04_U_addr),
			.i_fld_U_2_datain_0 (w_sub04_U_datain),
			.o_fld_U_2_dataout_0 (w_sub04_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub04_U_r_w),
			.i_fld_V_1_addr_0 (w_sub04_V_addr),
			.i_fld_V_1_datain_0 (w_sub04_V_datain),
			.o_fld_V_1_dataout_0 (w_sub04_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub04_V_r_w),
			.i_fld_result_3_addr_0 (w_sub04_result_addr),
			.i_fld_result_3_datain_0 (w_sub04_result_datain),
			.o_fld_result_3_dataout_0 (w_sub04_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub04_result_r_w),
			.o_run_busy (w_sub04_run_busy),
			.i_run_req (r_sub04_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub17
		sub17_inst(
			.i_fld_T_0_addr_0 (w_sub17_T_addr),
			.i_fld_T_0_datain_0 (w_sub17_T_datain),
			.o_fld_T_0_dataout_0 (w_sub17_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub17_T_r_w),
			.i_fld_U_2_addr_0 (w_sub17_U_addr),
			.i_fld_U_2_datain_0 (w_sub17_U_datain),
			.o_fld_U_2_dataout_0 (w_sub17_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub17_U_r_w),
			.i_fld_V_1_addr_0 (w_sub17_V_addr),
			.i_fld_V_1_datain_0 (w_sub17_V_datain),
			.o_fld_V_1_dataout_0 (w_sub17_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub17_V_r_w),
			.i_fld_result_3_addr_0 (w_sub17_result_addr),
			.i_fld_result_3_datain_0 (w_sub17_result_datain),
			.o_fld_result_3_dataout_0 (w_sub17_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub17_result_r_w),
			.o_run_busy (w_sub17_run_busy),
			.i_run_req (r_sub17_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub10
		sub10_inst(
			.i_fld_T_0_addr_0 (w_sub10_T_addr),
			.i_fld_T_0_datain_0 (w_sub10_T_datain),
			.o_fld_T_0_dataout_0 (w_sub10_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub10_T_r_w),
			.i_fld_U_2_addr_0 (w_sub10_U_addr),
			.i_fld_U_2_datain_0 (w_sub10_U_datain),
			.o_fld_U_2_dataout_0 (w_sub10_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub10_U_r_w),
			.i_fld_V_1_addr_0 (w_sub10_V_addr),
			.i_fld_V_1_datain_0 (w_sub10_V_datain),
			.o_fld_V_1_dataout_0 (w_sub10_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub10_V_r_w),
			.i_fld_result_3_addr_0 (w_sub10_result_addr),
			.i_fld_result_3_datain_0 (w_sub10_result_datain),
			.o_fld_result_3_dataout_0 (w_sub10_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub10_result_r_w),
			.o_run_busy (w_sub10_run_busy),
			.i_run_req (r_sub10_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub20
		sub20_inst(
			.i_fld_T_0_addr_0 (w_sub20_T_addr),
			.i_fld_T_0_datain_0 (w_sub20_T_datain),
			.o_fld_T_0_dataout_0 (w_sub20_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub20_T_r_w),
			.i_fld_U_2_addr_0 (w_sub20_U_addr),
			.i_fld_U_2_datain_0 (w_sub20_U_datain),
			.o_fld_U_2_dataout_0 (w_sub20_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub20_U_r_w),
			.i_fld_V_1_addr_0 (w_sub20_V_addr),
			.i_fld_V_1_datain_0 (w_sub20_V_datain),
			.o_fld_V_1_dataout_0 (w_sub20_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub20_V_r_w),
			.i_fld_result_3_addr_0 (w_sub20_result_addr),
			.i_fld_result_3_datain_0 (w_sub20_result_datain),
			.o_fld_result_3_dataout_0 (w_sub20_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub20_result_r_w),
			.o_run_busy (w_sub20_run_busy),
			.i_run_req (r_sub20_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub21
		sub21_inst(
			.i_fld_T_0_addr_0 (w_sub21_T_addr),
			.i_fld_T_0_datain_0 (w_sub21_T_datain),
			.o_fld_T_0_dataout_0 (w_sub21_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub21_T_r_w),
			.i_fld_U_2_addr_0 (w_sub21_U_addr),
			.i_fld_U_2_datain_0 (w_sub21_U_datain),
			.o_fld_U_2_dataout_0 (w_sub21_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub21_U_r_w),
			.i_fld_V_1_addr_0 (w_sub21_V_addr),
			.i_fld_V_1_datain_0 (w_sub21_V_datain),
			.o_fld_V_1_dataout_0 (w_sub21_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub21_V_r_w),
			.i_fld_result_3_addr_0 (w_sub21_result_addr),
			.i_fld_result_3_datain_0 (w_sub21_result_datain),
			.o_fld_result_3_dataout_0 (w_sub21_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub21_result_r_w),
			.o_run_busy (w_sub21_run_busy),
			.i_run_req (r_sub21_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(9), .WORDS(484) )
		dpram_T_0(
			.clk (clock),
			.ce_0 (w_fld_T_0_ce_0),
			.addr_0 (w_fld_T_0_addr_0),
			.datain_0 (w_fld_T_0_datain_0),
			.dataout_0 (w_fld_T_0_dataout_0),
			.r_w_0 (w_fld_T_0_r_w_0),
			.ce_1 (w_fld_T_0_ce_1),
			.addr_1 (r_fld_T_0_addr_1),
			.datain_1 (r_fld_T_0_datain_1),
			.dataout_1 (w_fld_T_0_dataout_1),
			.r_w_1 (r_fld_T_0_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(9), .WORDS(484) )
		dpram_TT_1(
			.clk (clock),
			.ce_0 (w_fld_TT_1_ce_0),
			.addr_0 (w_fld_TT_1_addr_0),
			.datain_0 (w_fld_TT_1_datain_0),
			.dataout_0 (w_fld_TT_1_dataout_0),
			.r_w_0 (w_fld_TT_1_r_w_0),
			.ce_1 (w_fld_TT_1_ce_1),
			.addr_1 (r_fld_TT_1_addr_1),
			.datain_1 (r_fld_TT_1_datain_1),
			.dataout_1 (w_fld_TT_1_dataout_1),
			.r_w_1 (r_fld_TT_1_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(9), .WORDS(484) )
		dpram_U_2(
			.clk (clock),
			.ce_0 (w_fld_U_2_ce_0),
			.addr_0 (w_fld_U_2_addr_0),
			.datain_0 (w_fld_U_2_datain_0),
			.dataout_0 (w_fld_U_2_dataout_0),
			.r_w_0 (w_fld_U_2_r_w_0),
			.ce_1 (w_fld_U_2_ce_1),
			.addr_1 (r_fld_U_2_addr_1),
			.datain_1 (r_fld_U_2_datain_1),
			.dataout_1 (w_fld_U_2_dataout_1),
			.r_w_1 (r_fld_U_2_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(9), .WORDS(484) )
		dpram_V_3(
			.clk (clock),
			.ce_0 (w_fld_V_3_ce_0),
			.addr_0 (w_fld_V_3_addr_0),
			.datain_0 (w_fld_V_3_datain_0),
			.dataout_0 (w_fld_V_3_dataout_0),
			.r_w_0 (w_fld_V_3_r_w_0),
			.ce_1 (w_fld_V_3_ce_1),
			.addr_1 (r_fld_V_3_addr_1),
			.datain_1 (r_fld_V_3_datain_1),
			.dataout_1 (w_fld_V_3_dataout_1),
			.r_w_1 (r_fld_V_3_r_w_1)
		);

	DivInt
		DivInt_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.dividend (r_ip_DivInt_dividend_0),
			.divisor (r_ip_DivInt_divisor_0),
			.fractional (w_ip_DivInt_fractional_0),
			.quotient (w_ip_DivInt_quotient_0)
		);

	AddFloat
		AddFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_AddFloat_portA_0),
			.b (r_ip_AddFloat_portB_0),
			.result (w_ip_AddFloat_result_0)
		);

	MultFloat
		MultFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_MultFloat_multiplicand_0),
			.b (r_ip_MultFloat_multiplier_0),
			.result (w_ip_MultFloat_product_0)
		);

	FixedToFloat
		FixedToFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_FixedToFloat_fixed_0),
			.result (w_ip_FixedToFloat_floating_0)
		);

	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_ip_DivInt_dividend_0 <= r_run_mx_32;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_ip_DivInt_dividend_0 <= r_run_mx_32;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_ip_DivInt_divisor_0 <= w_sys_tmp1966;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_ip_DivInt_divisor_0 <= w_sys_tmp1970;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hc) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h14)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp39;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp38[31], w_sys_tmp38[30:0] };

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp129[31], w_sys_tmp129[30:0] };

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp38[31], w_sys_tmp38[30:0] };

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp129[31], w_sys_tmp129[30:0] };

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp38[31], w_sys_tmp38[30:0] };

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp38[31], w_sys_tmp38[30:0] };

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp38[31], w_sys_tmp38[30:0] };

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1b)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp19;

									end
									else
									if((r_sys_run_step==7'hc) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h16)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp37;

									end
									else
									if((r_sys_run_step==7'h13) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h1a)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp4_float;

									end
									else
									if((7'h7<=r_sys_run_step && r_sys_run_step<=7'hb) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'hf)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_dy_36;

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp0_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h15) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h1b)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==7'h13) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h1a)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==7'he) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h16)) begin
										r_ip_MultFloat_multiplier_0 <= r_run_YY_41;

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp38;

									end
									else
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'hf)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp4_float;

									end
									else
									if((7'h7<=r_sys_run_step && r_sys_run_step<=7'hb)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp20;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_ip_FixedToFloat_fixed_0 <= w_sys_tmp21;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						7'h4f: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_return <= 32'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4c: begin
							r_sys_run_return <= r_sys_tmp21_float;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 7'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h0: begin
							r_sys_run_phase <= 7'h2;
						end

						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h4;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h5;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp13) ? 7'h9 : 7'hf);

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h5;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'ha;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp16) ? 7'hd : 7'h6);

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h20)) begin
										r_sys_run_phase <= 7'ha;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h10;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp227) ? 7'h13 : 7'h15);

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6d)) begin
										r_sys_run_phase <= 7'h10;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h16;

									end
								end

							endcase
						end

						7'h16: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1529) ? 7'h19 : 7'h1b);

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1c)) begin
										r_sys_run_phase <= 7'h16;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h1c;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1858) ? 7'h20 : 7'h4d);

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h1c;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h21;

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1861) ? 7'h24 : 7'h26);

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_run_phase <= 7'h21;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h27;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1878) ? 7'h2a : 7'h2c);

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_phase <= 7'h27;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h2d;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h25)) begin
										r_sys_run_phase <= ((w_sys_tmp1967) ? 7'h30 : 7'h32);

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_run_phase <= 7'h2d;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h33;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2014) ? 7'h36 : 7'h38);

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6d)) begin
										r_sys_run_phase <= 7'h33;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h39;

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2668) ? 7'h3c : 7'h3d);

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1c)) begin
										r_sys_run_phase <= 7'h39;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h18: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_phase <= 7'h3f;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h18: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_phase <= 7'h41;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h42;

									end
								end

							endcase
						end

						7'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2836) ? 7'h45 : 7'h47);

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4d)) begin
										r_sys_run_phase <= 7'h42;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h48;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3226) ? 7'h4b : 7'h1d);

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h14)) begin
										r_sys_run_phase <= 7'h48;

									end
								end

							endcase
						end

						7'h4c: begin
							r_sys_run_phase <= 7'h4f;
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_run_phase <= 7'h4c;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sys_run_phase <= 7'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 5'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h20)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h16: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1c)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h25)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h25)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1c)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h14)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 7'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h20)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h1f)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6d)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h16: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1c)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h1b)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h1) || (r_sys_run_step==7'h2)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'hc)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h25)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h24)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h25)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h24)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h5)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6d)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1c)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h1b)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4d)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h4c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h14)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h1)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						7'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						7'h4f: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_T_0_addr_1 <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp23[8:0] );

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1865[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1869[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1873[8:0] );

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1) || (r_sys_run_step==7'h3) || (r_sys_run_step==7'h5) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'h9) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'hd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1887[8:0] );

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h2) || (r_sys_run_step==7'h4) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'hc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1882[8:0] );

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1973[8:0] );

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h62) || (r_sys_run_step==7'h64)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2607[8:0] );

									end
									else
									if((r_sys_run_step==7'h59)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2553[8:0] );

									end
									else
									if((r_sys_run_step==7'h44)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2427[8:0] );

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2049[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2067[8:0] );

									end
									else
									if((r_sys_run_step==7'h1f) || (r_sys_run_step==7'h21)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2205[8:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2145[8:0] );

									end
									else
									if((r_sys_run_step==7'h51)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2505[8:0] );

									end
									else
									if((r_sys_run_step==7'h39)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2361[8:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2193[8:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2169[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2019[8:0] );

									end
									else
									if((r_sys_run_step==7'h3f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2397[8:0] );

									end
									else
									if((r_sys_run_step==7'h50)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2499[8:0] );

									end
									else
									if((r_sys_run_step==7'h69)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2649[8:0] );

									end
									else
									if((r_sys_run_step==7'h5b) || (r_sys_run_step==7'h5d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2565[8:0] );

									end
									else
									if((r_sys_run_step==7'h4b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2469[8:0] );

									end
									else
									if((r_sys_run_step==7'h4a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2463[8:0] );

									end
									else
									if((r_sys_run_step==7'h34)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2331[8:0] );

									end
									else
									if((r_sys_run_step==7'h23)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2229[8:0] );

									end
									else
									if((r_sys_run_step==7'h5c) || (r_sys_run_step==7'h5e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2571[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2073[8:0] );

									end
									else
									if((r_sys_run_step==7'h33)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2325[8:0] );

									end
									else
									if((r_sys_run_step==7'h2c) || (r_sys_run_step==7'h2e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2283[8:0] );

									end
									else
									if((r_sys_run_step==7'h37)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2349[8:0] );

									end
									else
									if((r_sys_run_step==7'h60)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2595[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2031[8:0] );

									end
									else
									if((r_sys_run_step==7'h25) || (r_sys_run_step==7'h27)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2241[8:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2199[8:0] );

									end
									else
									if((r_sys_run_step==7'h53)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2517[8:0] );

									end
									else
									if((r_sys_run_step==7'h45)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2433[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2175[8:0] );

									end
									else
									if((r_sys_run_step==7'h4f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2493[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2025[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2109[8:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2163[8:0] );

									end
									else
									if((r_sys_run_step==7'h4e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2487[8:0] );

									end
									else
									if((r_sys_run_step==7'h36)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2343[8:0] );

									end
									else
									if((r_sys_run_step==7'hb) || (r_sys_run_step==7'hd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2085[8:0] );

									end
									else
									if((r_sys_run_step==7'h40) || (r_sys_run_step==7'h42)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2403[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2181[8:0] );

									end
									else
									if((r_sys_run_step==7'h20) || (r_sys_run_step==7'h22)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2211[8:0] );

									end
									else
									if((r_sys_run_step==7'h38)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2355[8:0] );

									end
									else
									if((r_sys_run_step==7'h29)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2265[8:0] );

									end
									else
									if((r_sys_run_step==7'h31) || (r_sys_run_step==7'h32)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2313[8:0] );

									end
									else
									if((r_sys_run_step==7'h61) || (r_sys_run_step==7'h63)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2601[8:0] );

									end
									else
									if((r_sys_run_step==7'h16) || (r_sys_run_step==7'h17)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2151[8:0] );

									end
									else
									if((r_sys_run_step==7'h56) || (r_sys_run_step==7'h58)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2535[8:0] );

									end
									else
									if((r_sys_run_step==7'h26) || (r_sys_run_step==7'h28)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2247[8:0] );

									end
									else
									if((r_sys_run_step==7'h24)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2235[8:0] );

									end
									else
									if((r_sys_run_step==7'h52)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2511[8:0] );

									end
									else
									if((r_sys_run_step==7'h2b) || (r_sys_run_step==7'h2d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2277[8:0] );

									end
									else
									if((r_sys_run_step==7'h41) || (r_sys_run_step==7'h43)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2409[8:0] );

									end
									else
									if((r_sys_run_step==7'h46) || (r_sys_run_step==7'h48)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2439[8:0] );

									end
									else
									if((r_sys_run_step==7'h6b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2661[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2103[8:0] );

									end
									else
									if((r_sys_run_step==7'h3a) || (r_sys_run_step==7'h3c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2367[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2139[8:0] );

									end
									else
									if((r_sys_run_step==7'h5f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2589[8:0] );

									end
									else
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'hc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2079[8:0] );

									end
									else
									if((r_sys_run_step==7'h65)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2625[8:0] );

									end
									else
									if((r_sys_run_step==7'h3e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2391[8:0] );

									end
									else
									if((r_sys_run_step==7'h10) || (r_sys_run_step==7'h12)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2115[8:0] );

									end
									else
									if((r_sys_run_step==7'h6a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2655[8:0] );

									end
									else
									if((r_sys_run_step==7'h3b) || (r_sys_run_step==7'h3d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2373[8:0] );

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2337[8:0] );

									end
									else
									if((r_sys_run_step==7'h5a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2559[8:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2187[8:0] );

									end
									else
									if((r_sys_run_step==7'h67) || (r_sys_run_step==7'h68)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2637[8:0] );

									end
									else
									if((r_sys_run_step==7'h4c) || (r_sys_run_step==7'h4d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2475[8:0] );

									end
									else
									if((r_sys_run_step==7'h55) || (r_sys_run_step==7'h57)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2529[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2037[8:0] );

									end
									else
									if((r_sys_run_step==7'h2f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2301[8:0] );

									end
									else
									if((r_sys_run_step==7'h47) || (r_sys_run_step==7'h49)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2445[8:0] );

									end
									else
									if((r_sys_run_step==7'h2a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2271[8:0] );

									end
									else
									if((r_sys_run_step==7'h11) || (r_sys_run_step==7'h13)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2121[8:0] );

									end
									else
									if((r_sys_run_step==7'h66)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2631[8:0] );

									end
									else
									if((r_sys_run_step==7'h4) || (r_sys_run_step==7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2043[8:0] );

									end
									else
									if((r_sys_run_step==7'h54)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2523[8:0] );

									end
									else
									if((r_sys_run_step==7'h30)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2307[8:0] );

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4) || (r_sys_run_step==7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2697[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2757[8:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2799[8:0] );

									end
									else
									if((r_sys_run_step==7'h16) || (r_sys_run_step==7'h17)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2805[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2685[8:0] );

									end
									else
									if((r_sys_run_step==7'h11) || (r_sys_run_step==7'h13)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2775[8:0] );

									end
									else
									if((r_sys_run_step==7'h10) || (r_sys_run_step==7'h12)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2769[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2763[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2727[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2721[8:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2817[8:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2823[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2673[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2679[8:0] );

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2703[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2691[8:0] );

									end
									else
									if((r_sys_run_step==7'hb) || (r_sys_run_step==7'hd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2739[8:0] );

									end
									else
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'hc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2733[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2829[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2793[8:0] );

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2885[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2910[8:0] );

									end
									else
									if((r_sys_run_step==7'h32)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3085[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2841[8:0] );

									end
									else
									if((r_sys_run_step==7'h49)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3200[8:0] );

									end
									else
									if((r_sys_run_step==7'h2c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3055[8:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2955[8:0] );

									end
									else
									if((r_sys_run_step==7'h2f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3070[8:0] );

									end
									else
									if((r_sys_run_step==7'h46)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3185[8:0] );

									end
									else
									if((r_sys_run_step==7'h3a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3125[8:0] );

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3100[8:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2995[8:0] );

									end
									else
									if((r_sys_run_step==7'h23)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3010[8:0] );

									end
									else
									if((r_sys_run_step==7'h37)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3110[8:0] );

									end
									else
									if((r_sys_run_step==7'h33)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3090[8:0] );

									end
									else
									if((r_sys_run_step==7'h41)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3160[8:0] );

									end
									else
									if((r_sys_run_step==7'h24)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3015[8:0] );

									end
									else
									if((r_sys_run_step==7'h28)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3035[8:0] );

									end
									else
									if((r_sys_run_step==7'h3d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3140[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2930[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2865[8:0] );

									end
									else
									if((r_sys_run_step==7'h3b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3130[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2915[8:0] );

									end
									else
									if((r_sys_run_step==7'h3e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3145[8:0] );

									end
									else
									if((r_sys_run_step==7'h43)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3170[8:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2895[8:0] );

									end
									else
									if((r_sys_run_step==7'h22)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3005[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2875[8:0] );

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3000[8:0] );

									end
									else
									if((r_sys_run_step==7'h36)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3105[8:0] );

									end
									else
									if((r_sys_run_step==7'h44)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3175[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2859[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2905[8:0] );

									end
									else
									if((r_sys_run_step==7'h25)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3020[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2880[8:0] );

									end
									else
									if((r_sys_run_step==7'h4c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3215[8:0] );

									end
									else
									if((r_sys_run_step==7'h34)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3095[8:0] );

									end
									else
									if((r_sys_run_step==7'h26)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3025[8:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2975[8:0] );

									end
									else
									if((r_sys_run_step==7'h2b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3050[8:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2980[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2925[8:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2940[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2920[8:0] );

									end
									else
									if((r_sys_run_step==7'h30)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3075[8:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2890[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2970[8:0] );

									end
									else
									if((r_sys_run_step==7'h2d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3060[8:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2985[8:0] );

									end
									else
									if((r_sys_run_step==7'h4b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3210[8:0] );

									end
									else
									if((r_sys_run_step==7'h2e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3065[8:0] );

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2945[8:0] );

									end
									else
									if((r_sys_run_step==7'h2a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3045[8:0] );

									end
									else
									if((r_sys_run_step==7'h39)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3120[8:0] );

									end
									else
									if((r_sys_run_step==7'h4a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3205[8:0] );

									end
									else
									if((r_sys_run_step==7'h27)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3030[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2853[8:0] );

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2950[8:0] );

									end
									else
									if((r_sys_run_step==7'h3c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3135[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2870[8:0] );

									end
									else
									if((r_sys_run_step==7'h29)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3040[8:0] );

									end
									else
									if((r_sys_run_step==7'h40)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3155[8:0] );

									end
									else
									if((r_sys_run_step==7'h42)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3165[8:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2960[8:0] );

									end
									else
									if((r_sys_run_step==7'h38)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3115[8:0] );

									end
									else
									if((r_sys_run_step==7'h4d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3220[8:0] );

									end
									else
									if((r_sys_run_step==7'h45)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3180[8:0] );

									end
									else
									if((r_sys_run_step==7'h31)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3080[8:0] );

									end
									else
									if((r_sys_run_step==7'h48)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3195[8:0] );

									end
									else
									if((r_sys_run_step==7'h47)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3190[8:0] );

									end
									else
									if((r_sys_run_step==7'h3f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3150[8:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2990[8:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2900[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2965[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2935[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2847[8:0] );

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3285[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3310[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3243[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3320[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3325[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3260[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3265[8:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3290[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3295[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3231[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3249[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3270[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3315[8:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3280[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3305[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3300[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3255[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3237[8:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3275[8:0] );

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3331[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp26;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp1872;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp1867;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp1885;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp1976;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h14)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp67_float;

									end
									else
									if((r_sys_run_step==7'h31)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp42_float;

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp69_float;

									end
									else
									if((r_sys_run_step==7'h25)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp52_float;

									end
									else
									if((r_sys_run_step==7'h29)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp44_float;

									end
									else
									if((r_sys_run_step==7'h43)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp55_float;

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp34_float;

									end
									else
									if((r_sys_run_step==7'h2a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp26_float;

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp47_float;

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==7'h4b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp53_float;

									end
									else
									if((r_sys_run_step==7'h39)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp35_float;

									end
									else
									if((r_sys_run_step==7'h4c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp36_float;

									end
									else
									if((r_sys_run_step==7'h32)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp24_float;

									end
									else
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h5)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp2843;

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp31_float;

									end
									else
									if((r_sys_run_step==7'h30)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp60_float;

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp64_float;

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp32_float;

									end
									else
									if((r_sys_run_step==7'h49)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp18_float;

									end
									else
									if((r_sys_run_step==7'h34)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp59_float;

									end
									else
									if((r_sys_run_step==7'h2c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp61_float;

									end
									else
									if((r_sys_run_step==7'h4a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==7'h3c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp40_float;

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp29_float;

									end
									else
									if((r_sys_run_step==7'h45)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp19_float;

									end
									else
									if((r_sys_run_step==7'h36)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp23_float;

									end
									else
									if((r_sys_run_step==7'h42)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==7'h40)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp39_float;

									end
									else
									if((r_sys_run_step==7'h3d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp21_float;

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==7'h3e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==7'h38)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp58_float;

									end
									else
									if((r_sys_run_step==7'h46)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp51_float;

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp50_float;

									end
									else
									if((r_sys_run_step==7'h3a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp22_float;

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp63_float;

									end
									else
									if((r_sys_run_step==7'h2b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==7'h2d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp43_float;

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp28_float;

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp68_float;

									end
									else
									if((r_sys_run_step==7'h23)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp27_float;

									end
									else
									if((r_sys_run_step==7'h26)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp45_float;

									end
									else
									if((r_sys_run_step==7'h47)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp54_float;

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp65_float;

									end
									else
									if((r_sys_run_step==7'h48)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp37_float;

									end
									else
									if((r_sys_run_step==7'h44)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp38_float;

									end
									else
									if((r_sys_run_step==7'h33)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp33_float;

									end
									else
									if((r_sys_run_step==7'h2e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp25_float;

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp14_float;

									end
									else
									if((r_sys_run_step==7'h22)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp46_float;

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp30_float;

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp49_float;

									end
									else
									if((r_sys_run_step==7'h24)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp41_float;

									end
									else
									if((r_sys_run_step==7'h41)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp20_float;

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==7'h28)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp62_float;

									end
									else
									if((r_sys_run_step==7'h27)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==7'h3b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp57_float;

									end
									else
									if((r_sys_run_step==7'h6) || (r_sys_run_step==7'h2f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp70_float;

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp48_float;

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp66_float;

									end
									else
									if((r_sys_run_step==7'h4d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==7'h3f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp56_float;

									end
									else
									if((r_sys_run_step==7'h37)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp6_float;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hb)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp18_float;

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp19_float;

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp9_float;

									end
									else
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h5)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp3233;

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp14_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_T_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h3)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6b)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h1a)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h4d)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h14)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_fld_T_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_TT_1_addr_1 <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_TT_1_addr_1 <= $signed( w_sys_tmp28[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_TT_1_datain_1 <= w_sys_tmp26;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_TT_1_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_TT_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4f: begin
							r_fld_TT_1_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_U_2_addr_1 <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h18) || (r_sys_run_step==7'h1a) || (7'h1c<=r_sys_run_step && r_sys_run_step<=7'h20)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp33[8:0] );

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h44)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp964[8:0] );

									end
									else
									if((r_sys_run_step==7'h36)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp880[8:0] );

									end
									else
									if((r_sys_run_step==7'h69)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1348[8:0] );

									end
									else
									if((r_sys_run_step==7'h29)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp640[8:0] );

									end
									else
									if((r_sys_run_step==7'h60)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1294[8:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp568[8:0] );

									end
									else
									if((r_sys_run_step==7'h5f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1288[8:0] );

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h7)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp262[8:0] );

									end
									else
									if((r_sys_run_step==7'h34)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp706[8:0] );

									end
									else
									if((r_sys_run_step==7'h6a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1354[8:0] );

									end
									else
									if((r_sys_run_step==7'h2f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp676[8:0] );

									end
									else
									if((r_sys_run_step==7'h4b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1006[8:0] );

									end
									else
									if((r_sys_run_step==7'h5b) || (r_sys_run_step==7'h5d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1264[8:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp376[8:0] );

									end
									else
									if((r_sys_run_step==7'h4e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1024[8:0] );

									end
									else
									if((r_sys_run_step==7'h20) || (r_sys_run_step==7'h22)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp586[8:0] );

									end
									else
									if((r_sys_run_step==7'h67) || (r_sys_run_step==7'h68)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1336[8:0] );

									end
									else
									if((r_sys_run_step==7'h26) || (r_sys_run_step==7'h28)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp622[8:0] );

									end
									else
									if((r_sys_run_step==7'h10) || (r_sys_run_step==7'h12)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp328[8:0] );

									end
									else
									if((r_sys_run_step==7'h54)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1222[8:0] );

									end
									else
									if((r_sys_run_step==7'h52)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1210[8:0] );

									end
									else
									if((r_sys_run_step==7'h61) || (r_sys_run_step==7'h63)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1300[8:0] );

									end
									else
									if((r_sys_run_step==7'h56) || (r_sys_run_step==7'h58)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1234[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp238[8:0] );

									end
									else
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'hc)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp292[8:0] );

									end
									else
									if((r_sys_run_step==7'h30)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp682[8:0] );

									end
									else
									if((r_sys_run_step==7'h3e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp928[8:0] );

									end
									else
									if((r_sys_run_step==7'h50)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1036[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp322[8:0] );

									end
									else
									if((r_sys_run_step==7'h53)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1216[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp388[8:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp382[8:0] );

									end
									else
									if((r_sys_run_step==7'h37)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp886[8:0] );

									end
									else
									if((r_sys_run_step==7'h6b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1360[8:0] );

									end
									else
									if((r_sys_run_step==7'h62) || (r_sys_run_step==7'h64)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1306[8:0] );

									end
									else
									if((r_sys_run_step==7'h2c) || (r_sys_run_step==7'h2e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp658[8:0] );

									end
									else
									if((r_sys_run_step==7'h39)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp898[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp250[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp280[8:0] );

									end
									else
									if((r_sys_run_step==7'h2a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp646[8:0] );

									end
									else
									if((r_sys_run_step==7'h38)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp892[8:0] );

									end
									else
									if((r_sys_run_step==7'h3f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp934[8:0] );

									end
									else
									if((r_sys_run_step==7'h4a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1000[8:0] );

									end
									else
									if((r_sys_run_step==7'h51)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1204[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp352[8:0] );

									end
									else
									if((r_sys_run_step==7'h66)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1330[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp316[8:0] );

									end
									else
									if((r_sys_run_step==7'h3a) || (r_sys_run_step==7'h3c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp904[8:0] );

									end
									else
									if((r_sys_run_step==7'h33)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp700[8:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp574[8:0] );

									end
									else
									if((r_sys_run_step==7'h5c) || (r_sys_run_step==7'h5e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1270[8:0] );

									end
									else
									if((r_sys_run_step==7'h25) || (r_sys_run_step==7'h27)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp616[8:0] );

									end
									else
									if((r_sys_run_step==7'h46) || (r_sys_run_step==7'h48)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp976[8:0] );

									end
									else
									if((r_sys_run_step==7'h11) || (r_sys_run_step==7'h13)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp334[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp286[8:0] );

									end
									else
									if((r_sys_run_step==7'h1f) || (r_sys_run_step==7'h21)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp580[8:0] );

									end
									else
									if((r_sys_run_step==7'h4c) || (r_sys_run_step==7'h4d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1012[8:0] );

									end
									else
									if((r_sys_run_step==7'h23)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp604[8:0] );

									end
									else
									if((r_sys_run_step==7'h5a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1258[8:0] );

									end
									else
									if((r_sys_run_step==7'h3b) || (r_sys_run_step==7'h3d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp910[8:0] );

									end
									else
									if((r_sys_run_step==7'h16) || (r_sys_run_step==7'h17)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp364[8:0] );

									end
									else
									if((r_sys_run_step==7'h45)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp970[8:0] );

									end
									else
									if((r_sys_run_step==7'h40) || (r_sys_run_step==7'h42)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp940[8:0] );

									end
									else
									if((r_sys_run_step==7'h47) || (r_sys_run_step==7'h49)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp982[8:0] );

									end
									else
									if((r_sys_run_step==7'hb) || (r_sys_run_step==7'hd)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp298[8:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp358[8:0] );

									end
									else
									if((r_sys_run_step==7'h4f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1030[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp556[8:0] );

									end
									else
									if((r_sys_run_step==7'h24)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp610[8:0] );

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp712[8:0] );

									end
									else
									if((r_sys_run_step==7'h65)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1324[8:0] );

									end
									else
									if((r_sys_run_step==7'h59)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1252[8:0] );

									end
									else
									if((r_sys_run_step==7'h2b) || (r_sys_run_step==7'h2d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp652[8:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp562[8:0] );

									end
									else
									if((r_sys_run_step==7'h31) || (r_sys_run_step==7'h32)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp688[8:0] );

									end
									else
									if((r_sys_run_step==7'h55) || (r_sys_run_step==7'h57)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1228[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp244[8:0] );

									end
									else
									if((r_sys_run_step==7'h41) || (r_sys_run_step==7'h43)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp946[8:0] );

									end
									else
									if((r_sys_run_step==7'h4) || (r_sys_run_step==7'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp256[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp232[8:0] );

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h15)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1660[8:0] );

									end
									else
									if((r_sys_run_step==7'h10) || (r_sys_run_step==7'h12)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1630[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1582[8:0] );

									end
									else
									if((r_sys_run_step==7'h16) || (r_sys_run_step==7'h17)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1666[8:0] );

									end
									else
									if((r_sys_run_step==7'h4) || (r_sys_run_step==7'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1558[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1588[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1534[8:0] );

									end
									else
									if((r_sys_run_step==7'h11) || (r_sys_run_step==7'h13)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1636[8:0] );

									end
									else
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'hc)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1594[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1546[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1624[8:0] );

									end
									else
									if((r_sys_run_step==7'hb) || (r_sys_run_step==7'hd)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1600[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1690[8:0] );

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h7)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1564[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1540[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1552[8:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1678[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1654[8:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1684[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1618[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h18) || (r_sys_run_step==7'h1a) || (7'h1c<=r_sys_run_step && r_sys_run_step<=7'h20)) begin
										r_fld_U_2_datain_1 <= w_sys_tmp19;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_U_2_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h18) || (r_sys_run_step==7'h1a) || (7'h1c<=r_sys_run_step && r_sys_run_step<=7'h20)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6b)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h1a)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_fld_U_2_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_V_3_addr_1 <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp42[8:0] );

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h44)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp964[8:0] );

									end
									else
									if((r_sys_run_step==7'h36)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp880[8:0] );

									end
									else
									if((r_sys_run_step==7'h69)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1348[8:0] );

									end
									else
									if((r_sys_run_step==7'h29)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp640[8:0] );

									end
									else
									if((r_sys_run_step==7'h60)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1294[8:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp568[8:0] );

									end
									else
									if((r_sys_run_step==7'h5f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1288[8:0] );

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h7)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp262[8:0] );

									end
									else
									if((r_sys_run_step==7'h34)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp706[8:0] );

									end
									else
									if((r_sys_run_step==7'h6a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1354[8:0] );

									end
									else
									if((r_sys_run_step==7'h2f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp676[8:0] );

									end
									else
									if((r_sys_run_step==7'h4b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1006[8:0] );

									end
									else
									if((r_sys_run_step==7'h5b) || (r_sys_run_step==7'h5d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1264[8:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp376[8:0] );

									end
									else
									if((r_sys_run_step==7'h4e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1024[8:0] );

									end
									else
									if((r_sys_run_step==7'h20) || (r_sys_run_step==7'h22)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp586[8:0] );

									end
									else
									if((r_sys_run_step==7'h67) || (r_sys_run_step==7'h68)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1336[8:0] );

									end
									else
									if((r_sys_run_step==7'h26) || (r_sys_run_step==7'h28)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp622[8:0] );

									end
									else
									if((r_sys_run_step==7'h10) || (r_sys_run_step==7'h12)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp328[8:0] );

									end
									else
									if((r_sys_run_step==7'h54)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1222[8:0] );

									end
									else
									if((r_sys_run_step==7'h52)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1210[8:0] );

									end
									else
									if((r_sys_run_step==7'h61) || (r_sys_run_step==7'h63)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1300[8:0] );

									end
									else
									if((r_sys_run_step==7'h56) || (r_sys_run_step==7'h58)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1234[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp238[8:0] );

									end
									else
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'hc)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp292[8:0] );

									end
									else
									if((r_sys_run_step==7'h30)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp682[8:0] );

									end
									else
									if((r_sys_run_step==7'h3e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp928[8:0] );

									end
									else
									if((r_sys_run_step==7'h50)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1036[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp322[8:0] );

									end
									else
									if((r_sys_run_step==7'h53)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1216[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp388[8:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp382[8:0] );

									end
									else
									if((r_sys_run_step==7'h37)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp886[8:0] );

									end
									else
									if((r_sys_run_step==7'h6b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1360[8:0] );

									end
									else
									if((r_sys_run_step==7'h62) || (r_sys_run_step==7'h64)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1306[8:0] );

									end
									else
									if((r_sys_run_step==7'h2c) || (r_sys_run_step==7'h2e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp658[8:0] );

									end
									else
									if((r_sys_run_step==7'h39)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp898[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp250[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp280[8:0] );

									end
									else
									if((r_sys_run_step==7'h2a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp646[8:0] );

									end
									else
									if((r_sys_run_step==7'h38)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp892[8:0] );

									end
									else
									if((r_sys_run_step==7'h3f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp934[8:0] );

									end
									else
									if((r_sys_run_step==7'h4a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1000[8:0] );

									end
									else
									if((r_sys_run_step==7'h51)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1204[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp352[8:0] );

									end
									else
									if((r_sys_run_step==7'h66)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1330[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp316[8:0] );

									end
									else
									if((r_sys_run_step==7'h3a) || (r_sys_run_step==7'h3c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp904[8:0] );

									end
									else
									if((r_sys_run_step==7'h33)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp700[8:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp574[8:0] );

									end
									else
									if((r_sys_run_step==7'h5c) || (r_sys_run_step==7'h5e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1270[8:0] );

									end
									else
									if((r_sys_run_step==7'h25) || (r_sys_run_step==7'h27)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp616[8:0] );

									end
									else
									if((r_sys_run_step==7'h46) || (r_sys_run_step==7'h48)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp976[8:0] );

									end
									else
									if((r_sys_run_step==7'h11) || (r_sys_run_step==7'h13)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp334[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp286[8:0] );

									end
									else
									if((r_sys_run_step==7'h1f) || (r_sys_run_step==7'h21)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp580[8:0] );

									end
									else
									if((r_sys_run_step==7'h4c) || (r_sys_run_step==7'h4d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1012[8:0] );

									end
									else
									if((r_sys_run_step==7'h23)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp604[8:0] );

									end
									else
									if((r_sys_run_step==7'h5a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1258[8:0] );

									end
									else
									if((r_sys_run_step==7'h3b) || (r_sys_run_step==7'h3d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp910[8:0] );

									end
									else
									if((r_sys_run_step==7'h16) || (r_sys_run_step==7'h17)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp364[8:0] );

									end
									else
									if((r_sys_run_step==7'h45)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp970[8:0] );

									end
									else
									if((r_sys_run_step==7'h40) || (r_sys_run_step==7'h42)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp940[8:0] );

									end
									else
									if((r_sys_run_step==7'h47) || (r_sys_run_step==7'h49)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp982[8:0] );

									end
									else
									if((r_sys_run_step==7'hb) || (r_sys_run_step==7'hd)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp298[8:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp358[8:0] );

									end
									else
									if((r_sys_run_step==7'h4f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1030[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp556[8:0] );

									end
									else
									if((r_sys_run_step==7'h24)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp610[8:0] );

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp712[8:0] );

									end
									else
									if((r_sys_run_step==7'h65)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1324[8:0] );

									end
									else
									if((r_sys_run_step==7'h59)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1252[8:0] );

									end
									else
									if((r_sys_run_step==7'h2b) || (r_sys_run_step==7'h2d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp652[8:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp562[8:0] );

									end
									else
									if((r_sys_run_step==7'h31) || (r_sys_run_step==7'h32)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp688[8:0] );

									end
									else
									if((r_sys_run_step==7'h55) || (r_sys_run_step==7'h57)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1228[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp244[8:0] );

									end
									else
									if((r_sys_run_step==7'h41) || (r_sys_run_step==7'h43)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp946[8:0] );

									end
									else
									if((r_sys_run_step==7'h4) || (r_sys_run_step==7'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp256[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp232[8:0] );

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h15)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1660[8:0] );

									end
									else
									if((r_sys_run_step==7'h10) || (r_sys_run_step==7'h12)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1630[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1582[8:0] );

									end
									else
									if((r_sys_run_step==7'h16) || (r_sys_run_step==7'h17)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1666[8:0] );

									end
									else
									if((r_sys_run_step==7'h4) || (r_sys_run_step==7'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1558[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1588[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1534[8:0] );

									end
									else
									if((r_sys_run_step==7'h11) || (r_sys_run_step==7'h13)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1636[8:0] );

									end
									else
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'hc)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1594[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1546[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1624[8:0] );

									end
									else
									if((r_sys_run_step==7'hb) || (r_sys_run_step==7'hd)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1600[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1690[8:0] );

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h7)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1564[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1540[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1552[8:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1678[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1654[8:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1684[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1618[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_datain_1 <= w_sys_tmp26;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_V_3_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6b)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h1a)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_fld_V_3_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_29 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_29 <= w_sys_tmp15;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_29 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6d)) begin
										r_run_k_29 <= w_sys_tmp1527;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_29 <= w_sys_tmp1528;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1c)) begin
										r_run_k_29 <= w_sys_tmp1857;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_29 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_run_k_29 <= w_sys_tmp1877;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_29 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6d)) begin
										r_run_k_29 <= w_sys_tmp2666;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_29 <= w_sys_tmp2667;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1c)) begin
										r_run_k_29 <= w_sys_tmp2834;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_29 <= w_sys_tmp2835;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4d)) begin
										r_run_k_29 <= w_sys_tmp3224;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_29 <= w_sys_tmp3225;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h14)) begin
										r_run_k_29 <= w_sys_tmp3329;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_30 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_30 <= w_sys_tmp49;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_30 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h2) || (r_sys_run_step==7'h4) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'hc)) begin
										r_run_j_30 <= w_sys_tmp1892;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h25)) begin
										r_run_j_30 <= w_sys_tmp1965;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_30 <= w_sys_tmp1977;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_n_31 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_n_31 <= w_sys_tmp1860;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_mx_32 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_my_33 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_dt_34 <= w_sys_tmp5;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_dx_35 <= w_sys_tmp7;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_dy_36 <= w_sys_tmp8;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_r1_37 <= w_sys_tmp9;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_r2_38 <= w_sys_tmp10;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_r3_39 <= w_sys_tmp11;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_r4_40 <= w_sys_tmp12;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hc) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h14)) begin
										r_run_YY_41 <= w_sys_tmp19;

									end
									else
									if((r_sys_run_step==7'h10) || (r_sys_run_step==7'h11)) begin
										r_run_YY_41 <= r_sys_tmp4_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_kx_42 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_ky_43 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_nlast_44 <= w_sys_tmp6;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_45 <= r_run_j_30;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_45 <= w_sys_tmp46;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_46 <= r_run_j_30;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h18) || (r_sys_run_step==7'h1a) || (7'h1c<=r_sys_run_step && r_sys_run_step<=7'h20)) begin
										r_run_copy1_j_46 <= w_sys_tmp47;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy2_j_47 <= r_run_j_30;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy2_j_47 <= w_sys_tmp48;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_48 <= r_run_j_30;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1) || (r_sys_run_step==7'h3) || (r_sys_run_step==7'h5) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'h9) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'hd)) begin
										r_run_copy0_j_48 <= w_sys_tmp1891;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub19_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub19_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6a)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp2637[8:0] );

									end
									else
									if((r_sys_run_step==7'h6c)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp2655[8:0] );

									end
									else
									if((r_sys_run_step==7'h6b)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp2649[8:0] );

									end
									else
									if((r_sys_run_step==7'h6d)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp2661[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h6a<=r_sys_run_step && r_sys_run_step<=7'h6d)) begin
										r_sub19_T_datain <= w_sys_tmp2021;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h6a<=r_sys_run_step && r_sys_run_step<=7'h6d)) begin
										r_sub19_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub19_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6b)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp1348[8:0] );

									end
									else
									if((r_sys_run_step==7'h6a)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp1336[8:0] );

									end
									else
									if((r_sys_run_step==7'h6d)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp1360[8:0] );

									end
									else
									if((r_sys_run_step==7'h6c)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp1354[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h6a<=r_sys_run_step && r_sys_run_step<=7'h6d)) begin
										r_sub19_V_datain <= w_sys_tmp396;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h6a<=r_sys_run_step && r_sys_run_step<=7'h6d)) begin
										r_sub19_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub19_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6b)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp1348[8:0] );

									end
									else
									if((r_sys_run_step==7'h6a)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp1336[8:0] );

									end
									else
									if((r_sys_run_step==7'h6d)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp1360[8:0] );

									end
									else
									if((r_sys_run_step==7'h6c)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp1354[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h6a<=r_sys_run_step && r_sys_run_step<=7'h6d)) begin
										r_sub19_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h6a<=r_sys_run_step && r_sys_run_step<=7'h6d)) begin
										r_sub19_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub19_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp3220[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp3215[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp3210[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h1) || (r_sys_run_step==7'h2)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub19_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub09_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub09_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h37)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp2337[8:0] );

									end
									else
									if((r_sys_run_step==7'h34)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp2313[8:0] );

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp2325[8:0] );

									end
									else
									if((r_sys_run_step==7'h36)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp2331[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h34<=r_sys_run_step && r_sys_run_step<=7'h37)) begin
										r_sub09_T_datain <= w_sys_tmp2021;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h34<=r_sys_run_step && r_sys_run_step<=7'h37)) begin
										r_sub09_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub09_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h34)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp688[8:0] );

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp700[8:0] );

									end
									else
									if((r_sys_run_step==7'h36)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp706[8:0] );

									end
									else
									if((r_sys_run_step==7'h37)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp712[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h34<=r_sys_run_step && r_sys_run_step<=7'h37)) begin
										r_sub09_V_datain <= w_sys_tmp396;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h34<=r_sys_run_step && r_sys_run_step<=7'h37)) begin
										r_sub09_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub09_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h34)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp688[8:0] );

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp700[8:0] );

									end
									else
									if((r_sys_run_step==7'h36)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp706[8:0] );

									end
									else
									if((r_sys_run_step==7'h37)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp712[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h34<=r_sys_run_step && r_sys_run_step<=7'h37)) begin
										r_sub09_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h34<=r_sys_run_step && r_sys_run_step<=7'h37)) begin
										r_sub09_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub09_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp3030[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp3020[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp3025[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h1) || (r_sys_run_step==7'h2)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub09_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub08_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub08_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h33)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp2313[8:0] );

									end
									else
									if((r_sys_run_step==7'h30)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp2283[8:0] );

									end
									else
									if((r_sys_run_step==7'h2f)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp2277[8:0] );

									end
									else
									if((r_sys_run_step==7'h31)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp2301[8:0] );

									end
									else
									if((r_sys_run_step==7'h32)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp2307[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2f<=r_sys_run_step && r_sys_run_step<=7'h33)) begin
										r_sub08_T_datain <= w_sys_tmp2021;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2f<=r_sys_run_step && r_sys_run_step<=7'h33)) begin
										r_sub08_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub08_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h33)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp688[8:0] );

									end
									else
									if((r_sys_run_step==7'h32)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp682[8:0] );

									end
									else
									if((r_sys_run_step==7'h31)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp676[8:0] );

									end
									else
									if((r_sys_run_step==7'h30)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp658[8:0] );

									end
									else
									if((r_sys_run_step==7'h2f)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp652[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2f<=r_sys_run_step && r_sys_run_step<=7'h33)) begin
										r_sub08_V_datain <= w_sys_tmp396;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2f<=r_sys_run_step && r_sys_run_step<=7'h33)) begin
										r_sub08_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub08_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h33)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp688[8:0] );

									end
									else
									if((r_sys_run_step==7'h32)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp682[8:0] );

									end
									else
									if((r_sys_run_step==7'h31)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp676[8:0] );

									end
									else
									if((r_sys_run_step==7'h30)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp658[8:0] );

									end
									else
									if((r_sys_run_step==7'h2f)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp652[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2f<=r_sys_run_step && r_sys_run_step<=7'h33)) begin
										r_sub08_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2f<=r_sys_run_step && r_sys_run_step<=7'h33)) begin
										r_sub08_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub08_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp3015[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp3005[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp3000[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp3010[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub08_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub24_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub24_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1a)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp2817[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp2823[8:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp2805[8:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp2829[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h19<=r_sys_run_step && r_sys_run_step<=7'h1c)) begin
										r_sub24_T_datain <= w_sys_tmp2675;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h19<=r_sys_run_step && r_sys_run_step<=7'h1c)) begin
										r_sub24_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub24_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h19)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp1666[8:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp1690[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp1678[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp1684[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h19<=r_sys_run_step && r_sys_run_step<=7'h1c)) begin
										r_sub24_V_datain <= w_sys_tmp1698;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h19<=r_sys_run_step && r_sys_run_step<=7'h1c)) begin
										r_sub24_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub24_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h19)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp1666[8:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp1690[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp1678[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp1684[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h19<=r_sys_run_step && r_sys_run_step<=7'h1c)) begin
										r_sub24_U_datain <= w_sys_tmp1536;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h19<=r_sys_run_step && r_sys_run_step<=7'h1c)) begin
										r_sub24_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub24_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp3320[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp3315[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp3325[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h1) || (r_sys_run_step==7'h2)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub24_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub22_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub22_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h10)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp2757[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp2775[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp2769[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp2763[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp2739[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp2733[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_sub22_T_datain <= w_sys_tmp2675;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_sub22_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub22_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h11)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp1624[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp1630[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp1600[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp1636[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp1594[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp1618[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_sub22_V_datain <= w_sys_tmp1698;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_sub22_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub22_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h11)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp1624[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp1630[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp1600[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp1636[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp1594[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp1618[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_sub22_U_datain <= w_sys_tmp1536;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_sub22_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub22_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp3290[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp3285[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp3280[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp3275[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub22_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub23_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub23_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h17)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp2799[8:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp2805[8:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp2775[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp2769[8:0] );

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp2793[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h14<=r_sys_run_step && r_sys_run_step<=7'h18)) begin
										r_sub23_T_datain <= w_sys_tmp2675;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h14<=r_sys_run_step && r_sys_run_step<=7'h18)) begin
										r_sub23_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub23_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h17)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp1660[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp1630[8:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp1666[8:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp1636[8:0] );

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp1654[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h14<=r_sys_run_step && r_sys_run_step<=7'h18)) begin
										r_sub23_V_datain <= w_sys_tmp1698;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h14<=r_sys_run_step && r_sys_run_step<=7'h18)) begin
										r_sub23_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub23_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h17)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp1660[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp1630[8:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp1666[8:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp1636[8:0] );

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp1654[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h14<=r_sys_run_step && r_sys_run_step<=7'h18)) begin
										r_sub23_U_datain <= w_sys_tmp1536;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h14<=r_sys_run_step && r_sys_run_step<=7'h18)) begin
										r_sub23_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub23_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp3310[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp3295[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp3305[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp3300[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub23_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub12_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub12_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h46)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp2427[8:0] );

									end
									else
									if((r_sys_run_step==7'h44)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp2403[8:0] );

									end
									else
									if((r_sys_run_step==7'h47)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp2433[8:0] );

									end
									else
									if((r_sys_run_step==7'h45)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp2409[8:0] );

									end
									else
									if((r_sys_run_step==7'h49)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp2445[8:0] );

									end
									else
									if((r_sys_run_step==7'h48)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp2439[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h44<=r_sys_run_step && r_sys_run_step<=7'h49)) begin
										r_sub12_T_datain <= w_sys_tmp2021;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h44<=r_sys_run_step && r_sys_run_step<=7'h49)) begin
										r_sub12_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub12_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h48)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp976[8:0] );

									end
									else
									if((r_sys_run_step==7'h46)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp964[8:0] );

									end
									else
									if((r_sys_run_step==7'h49)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp982[8:0] );

									end
									else
									if((r_sys_run_step==7'h45)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp946[8:0] );

									end
									else
									if((r_sys_run_step==7'h47)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp970[8:0] );

									end
									else
									if((r_sys_run_step==7'h44)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp940[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h44<=r_sys_run_step && r_sys_run_step<=7'h49)) begin
										r_sub12_V_datain <= w_sys_tmp396;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h44<=r_sys_run_step && r_sys_run_step<=7'h49)) begin
										r_sub12_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub12_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h48)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp976[8:0] );

									end
									else
									if((r_sys_run_step==7'h46)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp964[8:0] );

									end
									else
									if((r_sys_run_step==7'h49)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp982[8:0] );

									end
									else
									if((r_sys_run_step==7'h45)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp946[8:0] );

									end
									else
									if((r_sys_run_step==7'h47)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp970[8:0] );

									end
									else
									if((r_sys_run_step==7'h44)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp940[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h44<=r_sys_run_step && r_sys_run_step<=7'h49)) begin
										r_sub12_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h44<=r_sys_run_step && r_sys_run_step<=7'h49)) begin
										r_sub12_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub12_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp3090[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp3085[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp3075[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp3080[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub12_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h16)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp2139[8:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp2121[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp2115[8:0] );

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp2145[8:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp2151[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h14<=r_sys_run_step && r_sys_run_step<=7'h18)) begin
										r_sub03_T_datain <= w_sys_tmp2021;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h14<=r_sys_run_step && r_sys_run_step<=7'h18)) begin
										r_sub03_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub03_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h15)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp334[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp328[8:0] );

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp358[8:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp364[8:0] );

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp352[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h14<=r_sys_run_step && r_sys_run_step<=7'h18)) begin
										r_sub03_V_datain <= w_sys_tmp396;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h14<=r_sys_run_step && r_sys_run_step<=7'h18)) begin
										r_sub03_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub03_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h15)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp334[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp328[8:0] );

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp358[8:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp364[8:0] );

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp352[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h14<=r_sys_run_step && r_sys_run_step<=7'h18)) begin
										r_sub03_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h14<=r_sys_run_step && r_sys_run_step<=7'h18)) begin
										r_sub03_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub03_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2910[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2905[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2915[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2920[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub03_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'he)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp2079[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp2121[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp2085[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp2115[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp2109[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp2103[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_sub02_T_datain <= w_sys_tmp2021;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_sub02_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub02_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h11)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp322[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp334[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp328[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp316[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp298[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp292[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_sub02_V_datain <= w_sys_tmp396;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_sub02_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub02_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h11)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp322[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp334[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp328[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp316[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp298[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp292[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_sub02_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_sub02_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub02_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2885[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2895[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2890[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2900[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub02_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub11_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub11_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h40)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp2391[8:0] );

									end
									else
									if((r_sys_run_step==7'h42)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp2403[8:0] );

									end
									else
									if((r_sys_run_step==7'h43)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp2409[8:0] );

									end
									else
									if((r_sys_run_step==7'h41)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp2397[8:0] );

									end
									else
									if((r_sys_run_step==7'h3f)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp2373[8:0] );

									end
									else
									if((r_sys_run_step==7'h3e)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp2367[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h3e<=r_sys_run_step && r_sys_run_step<=7'h43)) begin
										r_sub11_T_datain <= w_sys_tmp2021;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h3e<=r_sys_run_step && r_sys_run_step<=7'h43)) begin
										r_sub11_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub11_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3e)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp904[8:0] );

									end
									else
									if((r_sys_run_step==7'h43)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp946[8:0] );

									end
									else
									if((r_sys_run_step==7'h3f)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp910[8:0] );

									end
									else
									if((r_sys_run_step==7'h41)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp934[8:0] );

									end
									else
									if((r_sys_run_step==7'h40)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp928[8:0] );

									end
									else
									if((r_sys_run_step==7'h42)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp940[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h3e<=r_sys_run_step && r_sys_run_step<=7'h43)) begin
										r_sub11_V_datain <= w_sys_tmp396;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h3e<=r_sys_run_step && r_sys_run_step<=7'h43)) begin
										r_sub11_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub11_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3e)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp904[8:0] );

									end
									else
									if((r_sys_run_step==7'h43)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp946[8:0] );

									end
									else
									if((r_sys_run_step==7'h3f)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp910[8:0] );

									end
									else
									if((r_sys_run_step==7'h41)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp934[8:0] );

									end
									else
									if((r_sys_run_step==7'h40)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp928[8:0] );

									end
									else
									if((r_sys_run_step==7'h42)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp940[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h3e<=r_sys_run_step && r_sys_run_step<=7'h43)) begin
										r_sub11_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h3e<=r_sys_run_step && r_sys_run_step<=7'h43)) begin
										r_sub11_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub11_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp3065[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp3055[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp3060[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h1) || (r_sys_run_step==7'h2)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub11_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub14_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub14_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h50)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp2487[8:0] );

									end
									else
									if((r_sys_run_step==7'h4f)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp2475[8:0] );

									end
									else
									if((r_sys_run_step==7'h51)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp2493[8:0] );

									end
									else
									if((r_sys_run_step==7'h52)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp2499[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h4f<=r_sys_run_step && r_sys_run_step<=7'h52)) begin
										r_sub14_T_datain <= w_sys_tmp2021;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h4f<=r_sys_run_step && r_sys_run_step<=7'h52)) begin
										r_sub14_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub14_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h52)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp1036[8:0] );

									end
									else
									if((r_sys_run_step==7'h50)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp1024[8:0] );

									end
									else
									if((r_sys_run_step==7'h4f)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp1012[8:0] );

									end
									else
									if((r_sys_run_step==7'h51)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp1030[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h4f<=r_sys_run_step && r_sys_run_step<=7'h52)) begin
										r_sub14_V_datain <= w_sys_tmp396;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h4f<=r_sys_run_step && r_sys_run_step<=7'h52)) begin
										r_sub14_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub14_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h52)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp1036[8:0] );

									end
									else
									if((r_sys_run_step==7'h50)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp1024[8:0] );

									end
									else
									if((r_sys_run_step==7'h4f)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp1012[8:0] );

									end
									else
									if((r_sys_run_step==7'h51)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp1030[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h4f<=r_sys_run_step && r_sys_run_step<=7'h52)) begin
										r_sub14_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h4f<=r_sys_run_step && r_sys_run_step<=7'h52)) begin
										r_sub14_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub14_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp3120[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp3125[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp3115[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h1) || (r_sys_run_step==7'h2)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub14_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hc)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp2079[8:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp2067[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp2049[8:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp2085[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp2043[8:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp2073[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h8<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub01_T_datain <= w_sys_tmp2021;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h8<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub01_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub01_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hb)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp286[8:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp280[8:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp298[8:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp292[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp262[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp256[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h8<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub01_V_datain <= w_sys_tmp396;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h8<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub01_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub01_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hb)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp286[8:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp280[8:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp298[8:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp292[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp262[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp256[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h8<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub01_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h8<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub01_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub01_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2865[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2870[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2875[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2880[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp2031[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp2049[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp2043[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp2037[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp2025[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp2019[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sub00_T_datain <= w_sys_tmp2021;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sub00_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub00_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp250[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp244[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp262[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp238[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp256[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp232[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sub00_V_datain <= w_sys_tmp396;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sub00_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub00_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp250[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp244[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp262[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp238[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp256[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp232[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sub00_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sub00_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub00_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp2841[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp2853[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp2859[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp2847[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub13_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub13_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4e)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp2475[8:0] );

									end
									else
									if((r_sys_run_step==7'h4b)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp2445[8:0] );

									end
									else
									if((r_sys_run_step==7'h4a)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp2439[8:0] );

									end
									else
									if((r_sys_run_step==7'h4d)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp2469[8:0] );

									end
									else
									if((r_sys_run_step==7'h4c)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp2463[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h4a<=r_sys_run_step && r_sys_run_step<=7'h4e)) begin
										r_sub13_T_datain <= w_sys_tmp2021;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h4a<=r_sys_run_step && r_sys_run_step<=7'h4e)) begin
										r_sub13_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub13_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4a)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp976[8:0] );

									end
									else
									if((r_sys_run_step==7'h4b)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp982[8:0] );

									end
									else
									if((r_sys_run_step==7'h4e)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp1012[8:0] );

									end
									else
									if((r_sys_run_step==7'h4d)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp1006[8:0] );

									end
									else
									if((r_sys_run_step==7'h4c)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp1000[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h4a<=r_sys_run_step && r_sys_run_step<=7'h4e)) begin
										r_sub13_V_datain <= w_sys_tmp396;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h4a<=r_sys_run_step && r_sys_run_step<=7'h4e)) begin
										r_sub13_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub13_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4a)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp976[8:0] );

									end
									else
									if((r_sys_run_step==7'h4b)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp982[8:0] );

									end
									else
									if((r_sys_run_step==7'h4e)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp1012[8:0] );

									end
									else
									if((r_sys_run_step==7'h4d)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp1006[8:0] );

									end
									else
									if((r_sys_run_step==7'h4c)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp1000[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h4a<=r_sys_run_step && r_sys_run_step<=7'h4e)) begin
										r_sub13_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h4a<=r_sys_run_step && r_sys_run_step<=7'h4e)) begin
										r_sub13_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub13_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp3100[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp3105[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp3110[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp3095[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub13_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub07_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub07_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2c)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp2271[8:0] );

									end
									else
									if((r_sys_run_step==7'h29)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp2241[8:0] );

									end
									else
									if((r_sys_run_step==7'h2b)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp2265[8:0] );

									end
									else
									if((r_sys_run_step==7'h2a)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp2247[8:0] );

									end
									else
									if((r_sys_run_step==7'h2e)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp2283[8:0] );

									end
									else
									if((r_sys_run_step==7'h2d)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp2277[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h29<=r_sys_run_step && r_sys_run_step<=7'h2e)) begin
										r_sub07_T_datain <= w_sys_tmp2021;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h29<=r_sys_run_step && r_sys_run_step<=7'h2e)) begin
										r_sub07_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub07_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2b)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp640[8:0] );

									end
									else
									if((r_sys_run_step==7'h2a)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp622[8:0] );

									end
									else
									if((r_sys_run_step==7'h2c)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp646[8:0] );

									end
									else
									if((r_sys_run_step==7'h2e)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp658[8:0] );

									end
									else
									if((r_sys_run_step==7'h29)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp616[8:0] );

									end
									else
									if((r_sys_run_step==7'h2d)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp652[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h29<=r_sys_run_step && r_sys_run_step<=7'h2e)) begin
										r_sub07_V_datain <= w_sys_tmp396;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h29<=r_sys_run_step && r_sys_run_step<=7'h2e)) begin
										r_sub07_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub07_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2b)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp640[8:0] );

									end
									else
									if((r_sys_run_step==7'h2a)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp622[8:0] );

									end
									else
									if((r_sys_run_step==7'h2c)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp646[8:0] );

									end
									else
									if((r_sys_run_step==7'h2e)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp658[8:0] );

									end
									else
									if((r_sys_run_step==7'h29)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp616[8:0] );

									end
									else
									if((r_sys_run_step==7'h2d)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp652[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h29<=r_sys_run_step && r_sys_run_step<=7'h2e)) begin
										r_sub07_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h29<=r_sys_run_step && r_sys_run_step<=7'h2e)) begin
										r_sub07_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub07_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2980[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2990[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2995[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2985[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub07_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub16_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub16_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5b)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp2553[8:0] );

									end
									else
									if((r_sys_run_step==7'h5c)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp2559[8:0] );

									end
									else
									if((r_sys_run_step==7'h5e)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp2571[8:0] );

									end
									else
									if((r_sys_run_step==7'h5a)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp2535[8:0] );

									end
									else
									if((r_sys_run_step==7'h59)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp2529[8:0] );

									end
									else
									if((r_sys_run_step==7'h5d)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp2565[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h59<=r_sys_run_step && r_sys_run_step<=7'h5e)) begin
										r_sub16_T_datain <= w_sys_tmp2021;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h59<=r_sys_run_step && r_sys_run_step<=7'h5e)) begin
										r_sub16_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub16_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h59)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp1228[8:0] );

									end
									else
									if((r_sys_run_step==7'h5a)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp1234[8:0] );

									end
									else
									if((r_sys_run_step==7'h5e)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp1270[8:0] );

									end
									else
									if((r_sys_run_step==7'h5c)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp1258[8:0] );

									end
									else
									if((r_sys_run_step==7'h5d)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp1264[8:0] );

									end
									else
									if((r_sys_run_step==7'h5b)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp1252[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h59<=r_sys_run_step && r_sys_run_step<=7'h5e)) begin
										r_sub16_V_datain <= w_sys_tmp396;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h59<=r_sys_run_step && r_sys_run_step<=7'h5e)) begin
										r_sub16_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub16_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h59)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp1228[8:0] );

									end
									else
									if((r_sys_run_step==7'h5a)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp1234[8:0] );

									end
									else
									if((r_sys_run_step==7'h5e)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp1270[8:0] );

									end
									else
									if((r_sys_run_step==7'h5c)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp1258[8:0] );

									end
									else
									if((r_sys_run_step==7'h5d)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp1264[8:0] );

									end
									else
									if((r_sys_run_step==7'h5b)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp1252[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h59<=r_sys_run_step && r_sys_run_step<=7'h5e)) begin
										r_sub16_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h59<=r_sys_run_step && r_sys_run_step<=7'h5e)) begin
										r_sub16_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub16_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp3150[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp3160[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp3155[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp3165[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub16_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub06_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub06_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h27)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp2241[8:0] );

									end
									else
									if((r_sys_run_step==7'h25)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp2229[8:0] );

									end
									else
									if((r_sys_run_step==7'h23)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp2205[8:0] );

									end
									else
									if((r_sys_run_step==7'h28)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp2247[8:0] );

									end
									else
									if((r_sys_run_step==7'h24)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp2211[8:0] );

									end
									else
									if((r_sys_run_step==7'h26)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp2235[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h23<=r_sys_run_step && r_sys_run_step<=7'h28)) begin
										r_sub06_T_datain <= w_sys_tmp2021;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h23<=r_sys_run_step && r_sys_run_step<=7'h28)) begin
										r_sub06_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub06_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h24)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp586[8:0] );

									end
									else
									if((r_sys_run_step==7'h28)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp622[8:0] );

									end
									else
									if((r_sys_run_step==7'h23)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp580[8:0] );

									end
									else
									if((r_sys_run_step==7'h25)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp604[8:0] );

									end
									else
									if((r_sys_run_step==7'h27)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp616[8:0] );

									end
									else
									if((r_sys_run_step==7'h26)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp610[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h23<=r_sys_run_step && r_sys_run_step<=7'h28)) begin
										r_sub06_V_datain <= w_sys_tmp396;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h23<=r_sys_run_step && r_sys_run_step<=7'h28)) begin
										r_sub06_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub06_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h24)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp586[8:0] );

									end
									else
									if((r_sys_run_step==7'h28)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp622[8:0] );

									end
									else
									if((r_sys_run_step==7'h23)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp580[8:0] );

									end
									else
									if((r_sys_run_step==7'h25)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp604[8:0] );

									end
									else
									if((r_sys_run_step==7'h27)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp616[8:0] );

									end
									else
									if((r_sys_run_step==7'h26)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp610[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h23<=r_sys_run_step && r_sys_run_step<=7'h28)) begin
										r_sub06_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h23<=r_sys_run_step && r_sys_run_step<=7'h28)) begin
										r_sub06_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub06_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2975[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2960[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2970[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2965[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub06_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub15_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub15_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h55)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp2517[8:0] );

									end
									else
									if((r_sys_run_step==7'h58)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp2535[8:0] );

									end
									else
									if((r_sys_run_step==7'h56)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp2523[8:0] );

									end
									else
									if((r_sys_run_step==7'h53)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp2505[8:0] );

									end
									else
									if((r_sys_run_step==7'h54)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp2511[8:0] );

									end
									else
									if((r_sys_run_step==7'h57)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp2529[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h53<=r_sys_run_step && r_sys_run_step<=7'h58)) begin
										r_sub15_T_datain <= w_sys_tmp2021;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h53<=r_sys_run_step && r_sys_run_step<=7'h58)) begin
										r_sub15_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub15_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h55)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp1216[8:0] );

									end
									else
									if((r_sys_run_step==7'h57)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp1228[8:0] );

									end
									else
									if((r_sys_run_step==7'h56)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp1222[8:0] );

									end
									else
									if((r_sys_run_step==7'h54)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp1210[8:0] );

									end
									else
									if((r_sys_run_step==7'h58)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp1234[8:0] );

									end
									else
									if((r_sys_run_step==7'h53)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp1204[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h53<=r_sys_run_step && r_sys_run_step<=7'h58)) begin
										r_sub15_V_datain <= w_sys_tmp396;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h53<=r_sys_run_step && r_sys_run_step<=7'h58)) begin
										r_sub15_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub15_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h55)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp1216[8:0] );

									end
									else
									if((r_sys_run_step==7'h57)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp1228[8:0] );

									end
									else
									if((r_sys_run_step==7'h56)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp1222[8:0] );

									end
									else
									if((r_sys_run_step==7'h54)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp1210[8:0] );

									end
									else
									if((r_sys_run_step==7'h58)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp1234[8:0] );

									end
									else
									if((r_sys_run_step==7'h53)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp1204[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h53<=r_sys_run_step && r_sys_run_step<=7'h58)) begin
										r_sub15_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h53<=r_sys_run_step && r_sys_run_step<=7'h58)) begin
										r_sub15_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub15_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp3140[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp3130[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp3145[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp3135[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub15_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub05_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub05_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1e)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp2187[8:0] );

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp2205[8:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp2199[8:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp2181[8:0] );

									end
									else
									if((r_sys_run_step==7'h22)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp2211[8:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp2193[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h1d<=r_sys_run_step && r_sys_run_step<=7'h22)) begin
										r_sub05_T_datain <= w_sys_tmp2021;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h1d<=r_sys_run_step && r_sys_run_step<=7'h22)) begin
										r_sub05_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub05_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h22)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp586[8:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp562[8:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp568[8:0] );

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp580[8:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp574[8:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp556[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h1d<=r_sys_run_step && r_sys_run_step<=7'h22)) begin
										r_sub05_V_datain <= w_sys_tmp396;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h1d<=r_sys_run_step && r_sys_run_step<=7'h22)) begin
										r_sub05_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub05_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h22)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp586[8:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp562[8:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp568[8:0] );

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp580[8:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp574[8:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp556[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h1d<=r_sys_run_step && r_sys_run_step<=7'h22)) begin
										r_sub05_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h1d<=r_sys_run_step && r_sys_run_step<=7'h22)) begin
										r_sub05_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub05_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2945[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2955[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2950[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2940[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub05_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub18_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub18_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h66)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp2607[8:0] );

									end
									else
									if((r_sys_run_step==7'h67)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp2625[8:0] );

									end
									else
									if((r_sys_run_step==7'h68)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp2631[8:0] );

									end
									else
									if((r_sys_run_step==7'h69)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp2637[8:0] );

									end
									else
									if((r_sys_run_step==7'h65)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp2601[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h65<=r_sys_run_step && r_sys_run_step<=7'h69)) begin
										r_sub18_T_datain <= w_sys_tmp2021;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h65<=r_sys_run_step && r_sys_run_step<=7'h69)) begin
										r_sub18_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub18_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h69)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp1336[8:0] );

									end
									else
									if((r_sys_run_step==7'h68)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp1330[8:0] );

									end
									else
									if((r_sys_run_step==7'h65)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp1300[8:0] );

									end
									else
									if((r_sys_run_step==7'h66)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp1306[8:0] );

									end
									else
									if((r_sys_run_step==7'h67)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp1324[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h65<=r_sys_run_step && r_sys_run_step<=7'h69)) begin
										r_sub18_V_datain <= w_sys_tmp396;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h65<=r_sys_run_step && r_sys_run_step<=7'h69)) begin
										r_sub18_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub18_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h69)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp1336[8:0] );

									end
									else
									if((r_sys_run_step==7'h68)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp1330[8:0] );

									end
									else
									if((r_sys_run_step==7'h65)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp1300[8:0] );

									end
									else
									if((r_sys_run_step==7'h66)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp1306[8:0] );

									end
									else
									if((r_sys_run_step==7'h67)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp1324[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h65<=r_sys_run_step && r_sys_run_step<=7'h69)) begin
										r_sub18_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h65<=r_sys_run_step && r_sys_run_step<=7'h69)) begin
										r_sub18_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub18_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp3190[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp3205[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp3200[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp3195[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub18_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub04_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub04_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h19)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp2151[8:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp2175[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp2169[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp2163[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h19<=r_sys_run_step && r_sys_run_step<=7'h1c)) begin
										r_sub04_T_datain <= w_sys_tmp2021;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h19<=r_sys_run_step && r_sys_run_step<=7'h1c)) begin
										r_sub04_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub04_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1c)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp388[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp382[8:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp364[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp376[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h19<=r_sys_run_step && r_sys_run_step<=7'h1c)) begin
										r_sub04_V_datain <= w_sys_tmp396;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h19<=r_sys_run_step && r_sys_run_step<=7'h1c)) begin
										r_sub04_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub04_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1c)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp388[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp382[8:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp364[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp376[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h19<=r_sys_run_step && r_sys_run_step<=7'h1c)) begin
										r_sub04_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h19<=r_sys_run_step && r_sys_run_step<=7'h1c)) begin
										r_sub04_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub04_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2930[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2925[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2935[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h1) || (r_sys_run_step==7'h2)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub04_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub17_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub17_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h64)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp2607[8:0] );

									end
									else
									if((r_sys_run_step==7'h62)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp2595[8:0] );

									end
									else
									if((r_sys_run_step==7'h61)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp2589[8:0] );

									end
									else
									if((r_sys_run_step==7'h60)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp2571[8:0] );

									end
									else
									if((r_sys_run_step==7'h63)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp2601[8:0] );

									end
									else
									if((r_sys_run_step==7'h5f)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp2565[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h5f<=r_sys_run_step && r_sys_run_step<=7'h64)) begin
										r_sub17_T_datain <= w_sys_tmp2021;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h5f<=r_sys_run_step && r_sys_run_step<=7'h64)) begin
										r_sub17_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub17_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h62)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp1294[8:0] );

									end
									else
									if((r_sys_run_step==7'h63)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp1300[8:0] );

									end
									else
									if((r_sys_run_step==7'h61)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp1288[8:0] );

									end
									else
									if((r_sys_run_step==7'h60)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp1270[8:0] );

									end
									else
									if((r_sys_run_step==7'h64)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp1306[8:0] );

									end
									else
									if((r_sys_run_step==7'h5f)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp1264[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h5f<=r_sys_run_step && r_sys_run_step<=7'h64)) begin
										r_sub17_V_datain <= w_sys_tmp396;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h5f<=r_sys_run_step && r_sys_run_step<=7'h64)) begin
										r_sub17_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub17_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h62)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp1294[8:0] );

									end
									else
									if((r_sys_run_step==7'h63)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp1300[8:0] );

									end
									else
									if((r_sys_run_step==7'h61)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp1288[8:0] );

									end
									else
									if((r_sys_run_step==7'h60)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp1270[8:0] );

									end
									else
									if((r_sys_run_step==7'h64)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp1306[8:0] );

									end
									else
									if((r_sys_run_step==7'h5f)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp1264[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h5f<=r_sys_run_step && r_sys_run_step<=7'h64)) begin
										r_sub17_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h5f<=r_sys_run_step && r_sys_run_step<=7'h64)) begin
										r_sub17_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub17_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp3185[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp3170[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp3180[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp3175[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub17_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub10_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub10_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h38)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp2343[8:0] );

									end
									else
									if((r_sys_run_step==7'h3a)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp2355[8:0] );

									end
									else
									if((r_sys_run_step==7'h3b)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp2361[8:0] );

									end
									else
									if((r_sys_run_step==7'h3d)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp2373[8:0] );

									end
									else
									if((r_sys_run_step==7'h3c)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp2367[8:0] );

									end
									else
									if((r_sys_run_step==7'h39)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp2349[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h38<=r_sys_run_step && r_sys_run_step<=7'h3d)) begin
										r_sub10_T_datain <= w_sys_tmp2021;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h38<=r_sys_run_step && r_sys_run_step<=7'h3d)) begin
										r_sub10_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub10_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h38)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp880[8:0] );

									end
									else
									if((r_sys_run_step==7'h3c)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp904[8:0] );

									end
									else
									if((r_sys_run_step==7'h3a)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp892[8:0] );

									end
									else
									if((r_sys_run_step==7'h39)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp886[8:0] );

									end
									else
									if((r_sys_run_step==7'h3d)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp910[8:0] );

									end
									else
									if((r_sys_run_step==7'h3b)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp898[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h38<=r_sys_run_step && r_sys_run_step<=7'h3d)) begin
										r_sub10_V_datain <= w_sys_tmp396;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h38<=r_sys_run_step && r_sys_run_step<=7'h3d)) begin
										r_sub10_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub10_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h38)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp880[8:0] );

									end
									else
									if((r_sys_run_step==7'h3c)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp904[8:0] );

									end
									else
									if((r_sys_run_step==7'h3a)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp892[8:0] );

									end
									else
									if((r_sys_run_step==7'h39)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp886[8:0] );

									end
									else
									if((r_sys_run_step==7'h3d)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp910[8:0] );

									end
									else
									if((r_sys_run_step==7'h3b)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp898[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h38<=r_sys_run_step && r_sys_run_step<=7'h3d)) begin
										r_sub10_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h38<=r_sys_run_step && r_sys_run_step<=7'h3d)) begin
										r_sub10_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub10_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp3045[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp3050[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp3070[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp3035[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp3040[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h4)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub10_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub20_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub20_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp2697[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp2673[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp2703[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp2679[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp2691[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp2685[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sub20_T_datain <= w_sys_tmp2675;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sub20_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub20_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp1546[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp1564[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp1558[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp1552[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp1540[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp1534[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sub20_V_datain <= w_sys_tmp1698;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sub20_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub20_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp1546[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp1564[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp1558[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp1552[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp1540[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp1534[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sub20_U_datain <= w_sys_tmp1536;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sub20_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub20_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp3249[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp3231[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp3243[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp3237[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub20_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub21_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub21_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp2697[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp2703[8:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp2739[8:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp2733[8:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp2727[8:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp2721[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h8<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub21_T_datain <= w_sys_tmp2675;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h8<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub21_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub21_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp1582[8:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp1600[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp1564[8:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp1588[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp1558[8:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp1594[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h8<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub21_V_datain <= w_sys_tmp1698;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h8<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub21_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub21_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp1582[8:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp1600[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp1564[8:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp1588[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp1558[8:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp1594[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h8<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub21_U_datain <= w_sys_tmp1536;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h8<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub21_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub21_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp3265[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp3270[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp3260[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp3255[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4f: begin
							r_sub21_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h16)) begin
										r_sys_tmp0_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp0_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h16)) begin
										r_sys_tmp1_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp1_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h12) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h19)) begin
										r_sys_tmp2_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp2_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h11) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h17)) begin
										r_sys_tmp3_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp3_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hc) || (r_sys_run_step==7'hd)) begin
										r_sys_tmp4_float <= w_ip_FixedToFloat_floating_0;

									end
									else
									if((r_sys_run_step==7'hf) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h19)) begin
										r_sys_tmp4_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp4_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp5_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp5_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp6_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp6_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp7_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp7_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp8_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp8_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp9_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp9_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp10_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp10_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp11_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp11_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp12_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp12_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp13_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp13_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp14_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp14_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp15_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp15_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp16_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp16_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp17_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp17_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp18_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp18_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp19_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp19_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp20_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp21_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp21_float <= w_sys_tmp3330;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp22_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp23_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp24_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp25_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp26_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp27_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp28_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp29_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp30_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp31_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp32_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp33_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp34_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp35_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp36_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp37_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp38_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp39_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp40_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp41_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp42_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp43_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp44_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp45_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp46_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp47_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp48_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp49_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp50_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp51_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp52_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp53_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp54_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp55_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp56_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp57_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp58_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp59_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp60_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp61_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp62_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp63_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp64_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp65_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp66_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp67_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp68_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp69_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp70_float <= w_sub01_result_dataout;

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sys_tmp70_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
