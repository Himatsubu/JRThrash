/*
TimeStamp:	2016/9/15		17:35
*/


module c1(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy	
);

	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 5:0] r_sys_run_phase;
	reg         [ 4:0] r_sys_run_stage;
	reg         [ 8:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 4:0] w_sys_run_stage_p1;
	wire        [ 8:0] w_sys_run_step_p1;
	wire signed [14:0] w_fld_u_0_addr_0;
	wire        [31:0] w_fld_u_0_datain_0;
	wire        [31:0] w_fld_u_0_dataout_0;
	wire               w_fld_u_0_r_w_0;
	wire               w_fld_u_0_ce_0;
	reg  signed [14:0] r_fld_u_0_addr_1;
	reg         [31:0] r_fld_u_0_datain_1;
	wire        [31:0] w_fld_u_0_dataout_1;
	reg                r_fld_u_0_r_w_1;
	wire               w_fld_u_0_ce_1;
	reg  signed [31:0] r_run_k_17;
	reg  signed [31:0] r_run_j_18;
	reg  signed [31:0] r_run_n_19;
	reg  signed [31:0] r_run_mx_20;
	reg  signed [31:0] r_run_my_21;
	reg  signed [31:0] r_run_nlast_22;
	reg  signed [31:0] r_run_copy0_j_23;
	reg  signed [31:0] r_run_copy1_j_24;
	reg  signed [31:0] r_run_copy2_j_25;
	reg                r_sub09_run_req;
	wire               w_sub09_run_busy;
	wire signed [14:0] w_sub09_u_addr;
	reg  signed [14:0] r_sub09_u_addr;
	wire        [31:0] w_sub09_u_datain;
	reg         [31:0] r_sub09_u_datain;
	wire        [31:0] w_sub09_u_dataout;
	wire               w_sub09_u_r_w;
	reg                r_sub09_u_r_w;
	wire signed [14:0] w_sub09_result_addr;
	reg  signed [14:0] r_sub09_result_addr;
	wire        [31:0] w_sub09_result_datain;
	reg         [31:0] r_sub09_result_datain;
	wire        [31:0] w_sub09_result_dataout;
	wire               w_sub09_result_r_w;
	reg                r_sub09_result_r_w;
	reg                r_sub08_run_req;
	wire               w_sub08_run_busy;
	wire signed [14:0] w_sub08_u_addr;
	reg  signed [14:0] r_sub08_u_addr;
	wire        [31:0] w_sub08_u_datain;
	reg         [31:0] r_sub08_u_datain;
	wire        [31:0] w_sub08_u_dataout;
	wire               w_sub08_u_r_w;
	reg                r_sub08_u_r_w;
	wire signed [14:0] w_sub08_result_addr;
	reg  signed [14:0] r_sub08_result_addr;
	wire        [31:0] w_sub08_result_datain;
	reg         [31:0] r_sub08_result_datain;
	wire        [31:0] w_sub08_result_dataout;
	wire               w_sub08_result_r_w;
	reg                r_sub08_result_r_w;
	reg                r_sub12_run_req;
	wire               w_sub12_run_busy;
	wire signed [14:0] w_sub12_u_addr;
	reg  signed [14:0] r_sub12_u_addr;
	wire        [31:0] w_sub12_u_datain;
	reg         [31:0] r_sub12_u_datain;
	wire        [31:0] w_sub12_u_dataout;
	wire               w_sub12_u_r_w;
	reg                r_sub12_u_r_w;
	wire signed [14:0] w_sub12_result_addr;
	reg  signed [14:0] r_sub12_result_addr;
	wire        [31:0] w_sub12_result_datain;
	reg         [31:0] r_sub12_result_datain;
	wire        [31:0] w_sub12_result_dataout;
	wire               w_sub12_result_r_w;
	reg                r_sub12_result_r_w;
	reg                r_sub03_run_req;
	wire               w_sub03_run_busy;
	wire signed [14:0] w_sub03_u_addr;
	reg  signed [14:0] r_sub03_u_addr;
	wire        [31:0] w_sub03_u_datain;
	reg         [31:0] r_sub03_u_datain;
	wire        [31:0] w_sub03_u_dataout;
	wire               w_sub03_u_r_w;
	reg                r_sub03_u_r_w;
	wire signed [14:0] w_sub03_result_addr;
	reg  signed [14:0] r_sub03_result_addr;
	wire        [31:0] w_sub03_result_datain;
	reg         [31:0] r_sub03_result_datain;
	wire        [31:0] w_sub03_result_dataout;
	wire               w_sub03_result_r_w;
	reg                r_sub03_result_r_w;
	reg                r_sub02_run_req;
	wire               w_sub02_run_busy;
	wire signed [14:0] w_sub02_u_addr;
	reg  signed [14:0] r_sub02_u_addr;
	wire        [31:0] w_sub02_u_datain;
	reg         [31:0] r_sub02_u_datain;
	wire        [31:0] w_sub02_u_dataout;
	wire               w_sub02_u_r_w;
	reg                r_sub02_u_r_w;
	wire signed [14:0] w_sub02_result_addr;
	reg  signed [14:0] r_sub02_result_addr;
	wire        [31:0] w_sub02_result_datain;
	reg         [31:0] r_sub02_result_datain;
	wire        [31:0] w_sub02_result_dataout;
	wire               w_sub02_result_r_w;
	reg                r_sub02_result_r_w;
	reg                r_sub11_run_req;
	wire               w_sub11_run_busy;
	wire signed [14:0] w_sub11_u_addr;
	reg  signed [14:0] r_sub11_u_addr;
	wire        [31:0] w_sub11_u_datain;
	reg         [31:0] r_sub11_u_datain;
	wire        [31:0] w_sub11_u_dataout;
	wire               w_sub11_u_r_w;
	reg                r_sub11_u_r_w;
	wire signed [14:0] w_sub11_result_addr;
	reg  signed [14:0] r_sub11_result_addr;
	wire        [31:0] w_sub11_result_datain;
	reg         [31:0] r_sub11_result_datain;
	wire        [31:0] w_sub11_result_dataout;
	wire               w_sub11_result_r_w;
	reg                r_sub11_result_r_w;
	reg                r_sub14_run_req;
	wire               w_sub14_run_busy;
	wire signed [14:0] w_sub14_u_addr;
	reg  signed [14:0] r_sub14_u_addr;
	wire        [31:0] w_sub14_u_datain;
	reg         [31:0] r_sub14_u_datain;
	wire        [31:0] w_sub14_u_dataout;
	wire               w_sub14_u_r_w;
	reg                r_sub14_u_r_w;
	wire signed [14:0] w_sub14_result_addr;
	reg  signed [14:0] r_sub14_result_addr;
	wire        [31:0] w_sub14_result_datain;
	reg         [31:0] r_sub14_result_datain;
	wire        [31:0] w_sub14_result_dataout;
	wire               w_sub14_result_r_w;
	reg                r_sub14_result_r_w;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [14:0] w_sub01_u_addr;
	reg  signed [14:0] r_sub01_u_addr;
	wire        [31:0] w_sub01_u_datain;
	reg         [31:0] r_sub01_u_datain;
	wire        [31:0] w_sub01_u_dataout;
	wire               w_sub01_u_r_w;
	reg                r_sub01_u_r_w;
	wire signed [14:0] w_sub01_result_addr;
	reg  signed [14:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub13_run_req;
	wire               w_sub13_run_busy;
	wire signed [14:0] w_sub13_u_addr;
	reg  signed [14:0] r_sub13_u_addr;
	wire        [31:0] w_sub13_u_datain;
	reg         [31:0] r_sub13_u_datain;
	wire        [31:0] w_sub13_u_dataout;
	wire               w_sub13_u_r_w;
	reg                r_sub13_u_r_w;
	wire signed [14:0] w_sub13_result_addr;
	reg  signed [14:0] r_sub13_result_addr;
	wire        [31:0] w_sub13_result_datain;
	reg         [31:0] r_sub13_result_datain;
	wire        [31:0] w_sub13_result_dataout;
	wire               w_sub13_result_r_w;
	reg                r_sub13_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [14:0] w_sub00_u_addr;
	reg  signed [14:0] r_sub00_u_addr;
	wire        [31:0] w_sub00_u_datain;
	reg         [31:0] r_sub00_u_datain;
	wire        [31:0] w_sub00_u_dataout;
	wire               w_sub00_u_r_w;
	reg                r_sub00_u_r_w;
	wire signed [14:0] w_sub00_result_addr;
	reg  signed [14:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	reg                r_sub07_run_req;
	wire               w_sub07_run_busy;
	wire signed [14:0] w_sub07_u_addr;
	reg  signed [14:0] r_sub07_u_addr;
	wire        [31:0] w_sub07_u_datain;
	reg         [31:0] r_sub07_u_datain;
	wire        [31:0] w_sub07_u_dataout;
	wire               w_sub07_u_r_w;
	reg                r_sub07_u_r_w;
	wire signed [14:0] w_sub07_result_addr;
	reg  signed [14:0] r_sub07_result_addr;
	wire        [31:0] w_sub07_result_datain;
	reg         [31:0] r_sub07_result_datain;
	wire        [31:0] w_sub07_result_dataout;
	wire               w_sub07_result_r_w;
	reg                r_sub07_result_r_w;
	reg                r_sub06_run_req;
	wire               w_sub06_run_busy;
	wire signed [14:0] w_sub06_u_addr;
	reg  signed [14:0] r_sub06_u_addr;
	wire        [31:0] w_sub06_u_datain;
	reg         [31:0] r_sub06_u_datain;
	wire        [31:0] w_sub06_u_dataout;
	wire               w_sub06_u_r_w;
	reg                r_sub06_u_r_w;
	wire signed [14:0] w_sub06_result_addr;
	reg  signed [14:0] r_sub06_result_addr;
	wire        [31:0] w_sub06_result_datain;
	reg         [31:0] r_sub06_result_datain;
	wire        [31:0] w_sub06_result_dataout;
	wire               w_sub06_result_r_w;
	reg                r_sub06_result_r_w;
	reg                r_sub15_run_req;
	wire               w_sub15_run_busy;
	wire signed [14:0] w_sub15_u_addr;
	reg  signed [14:0] r_sub15_u_addr;
	wire        [31:0] w_sub15_u_datain;
	reg         [31:0] r_sub15_u_datain;
	wire        [31:0] w_sub15_u_dataout;
	wire               w_sub15_u_r_w;
	reg                r_sub15_u_r_w;
	wire signed [14:0] w_sub15_result_addr;
	reg  signed [14:0] r_sub15_result_addr;
	wire        [31:0] w_sub15_result_datain;
	reg         [31:0] r_sub15_result_datain;
	wire        [31:0] w_sub15_result_dataout;
	wire               w_sub15_result_r_w;
	reg                r_sub15_result_r_w;
	reg                r_sub05_run_req;
	wire               w_sub05_run_busy;
	wire signed [14:0] w_sub05_u_addr;
	reg  signed [14:0] r_sub05_u_addr;
	wire        [31:0] w_sub05_u_datain;
	reg         [31:0] r_sub05_u_datain;
	wire        [31:0] w_sub05_u_dataout;
	wire               w_sub05_u_r_w;
	reg                r_sub05_u_r_w;
	wire signed [14:0] w_sub05_result_addr;
	reg  signed [14:0] r_sub05_result_addr;
	wire        [31:0] w_sub05_result_datain;
	reg         [31:0] r_sub05_result_datain;
	wire        [31:0] w_sub05_result_dataout;
	wire               w_sub05_result_r_w;
	reg                r_sub05_result_r_w;
	reg                r_sub04_run_req;
	wire               w_sub04_run_busy;
	wire signed [14:0] w_sub04_u_addr;
	reg  signed [14:0] r_sub04_u_addr;
	wire        [31:0] w_sub04_u_datain;
	reg         [31:0] r_sub04_u_datain;
	wire        [31:0] w_sub04_u_dataout;
	wire               w_sub04_u_r_w;
	reg                r_sub04_u_r_w;
	wire signed [14:0] w_sub04_result_addr;
	reg  signed [14:0] r_sub04_result_addr;
	wire        [31:0] w_sub04_result_datain;
	reg         [31:0] r_sub04_result_datain;
	wire        [31:0] w_sub04_result_dataout;
	wire               w_sub04_result_r_w;
	reg                r_sub04_result_r_w;
	reg                r_sub10_run_req;
	wire               w_sub10_run_busy;
	wire signed [14:0] w_sub10_u_addr;
	reg  signed [14:0] r_sub10_u_addr;
	wire        [31:0] w_sub10_u_datain;
	reg         [31:0] r_sub10_u_datain;
	wire        [31:0] w_sub10_u_dataout;
	wire               w_sub10_u_r_w;
	reg                r_sub10_u_r_w;
	wire signed [14:0] w_sub10_result_addr;
	reg  signed [14:0] r_sub10_result_addr;
	wire        [31:0] w_sub10_result_datain;
	reg         [31:0] r_sub10_result_datain;
	wire        [31:0] w_sub10_result_dataout;
	wire               w_sub10_result_r_w;
	reg                r_sub10_result_r_w;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg         [31:0] r_sys_tmp4_float;
	reg         [31:0] r_sys_tmp5_float;
	reg         [31:0] r_sys_tmp6_float;
	reg         [31:0] r_sys_tmp7_float;
	reg         [31:0] r_sys_tmp8_float;
	reg         [31:0] r_sys_tmp9_float;
	reg         [31:0] r_sys_tmp10_float;
	reg         [31:0] r_sys_tmp11_float;
	reg         [31:0] r_sys_tmp12_float;
	reg         [31:0] r_sys_tmp13_float;
	reg         [31:0] r_sys_tmp14_float;
	reg         [31:0] r_sys_tmp15_float;
	reg         [31:0] r_sys_tmp16_float;
	reg         [31:0] r_sys_tmp17_float;
	reg         [31:0] r_sys_tmp18_float;
	reg         [31:0] r_sys_tmp19_float;
	reg         [31:0] r_sys_tmp20_float;
	reg         [31:0] r_sys_tmp21_float;
	reg         [31:0] r_sys_tmp22_float;
	reg         [31:0] r_sys_tmp23_float;
	reg         [31:0] r_sys_tmp24_float;
	reg         [31:0] r_sys_tmp25_float;
	reg         [31:0] r_sys_tmp26_float;
	reg         [31:0] r_sys_tmp27_float;
	reg         [31:0] r_sys_tmp28_float;
	reg         [31:0] r_sys_tmp29_float;
	reg         [31:0] r_sys_tmp30_float;
	reg         [31:0] r_sys_tmp31_float;
	reg         [31:0] r_sys_tmp32_float;
	reg         [31:0] r_sys_tmp33_float;
	reg         [31:0] r_sys_tmp34_float;
	reg         [31:0] r_sys_tmp35_float;
	reg         [31:0] r_sys_tmp36_float;
	reg         [31:0] r_sys_tmp37_float;
	reg         [31:0] r_sys_tmp38_float;
	reg         [31:0] r_sys_tmp39_float;
	reg         [31:0] r_sys_tmp40_float;
	reg         [31:0] r_sys_tmp41_float;
	reg         [31:0] r_sys_tmp42_float;
	reg         [31:0] r_sys_tmp43_float;
	reg         [31:0] r_sys_tmp44_float;
	reg         [31:0] r_sys_tmp45_float;
	reg         [31:0] r_sys_tmp46_float;
	reg         [31:0] r_sys_tmp47_float;
	reg         [31:0] r_sys_tmp48_float;
	reg         [31:0] r_sys_tmp49_float;
	reg         [31:0] r_sys_tmp50_float;
	reg         [31:0] r_sys_tmp51_float;
	reg         [31:0] r_sys_tmp52_float;
	reg         [31:0] r_sys_tmp53_float;
	reg         [31:0] r_sys_tmp54_float;
	reg         [31:0] r_sys_tmp55_float;
	reg         [31:0] r_sys_tmp56_float;
	reg         [31:0] r_sys_tmp57_float;
	reg         [31:0] r_sys_tmp58_float;
	reg         [31:0] r_sys_tmp59_float;
	reg         [31:0] r_sys_tmp60_float;
	reg         [31:0] r_sys_tmp61_float;
	reg         [31:0] r_sys_tmp62_float;
	reg         [31:0] r_sys_tmp63_float;
	reg         [31:0] r_sys_tmp64_float;
	reg         [31:0] r_sys_tmp65_float;
	reg         [31:0] r_sys_tmp66_float;
	reg         [31:0] r_sys_tmp67_float;
	reg         [31:0] r_sys_tmp68_float;
	reg         [31:0] r_sys_tmp69_float;
	reg         [31:0] r_sys_tmp70_float;
	reg         [31:0] r_sys_tmp71_float;
	reg         [31:0] r_sys_tmp72_float;
	reg         [31:0] r_sys_tmp73_float;
	reg         [31:0] r_sys_tmp74_float;
	reg         [31:0] r_sys_tmp75_float;
	reg         [31:0] r_sys_tmp76_float;
	reg         [31:0] r_sys_tmp77_float;
	reg         [31:0] r_sys_tmp78_float;
	reg         [31:0] r_sys_tmp79_float;
	reg         [31:0] r_sys_tmp80_float;
	reg         [31:0] r_sys_tmp81_float;
	reg         [31:0] r_sys_tmp82_float;
	reg         [31:0] r_sys_tmp83_float;
	reg         [31:0] r_sys_tmp84_float;
	reg         [31:0] r_sys_tmp85_float;
	reg         [31:0] r_sys_tmp86_float;
	reg         [31:0] r_sys_tmp87_float;
	reg         [31:0] r_sys_tmp88_float;
	reg         [31:0] r_sys_tmp89_float;
	reg         [31:0] r_sys_tmp90_float;
	reg         [31:0] r_sys_tmp91_float;
	reg         [31:0] r_sys_tmp92_float;
	reg         [31:0] r_sys_tmp93_float;
	reg         [31:0] r_sys_tmp94_float;
	reg         [31:0] r_sys_tmp95_float;
	reg         [31:0] r_sys_tmp96_float;
	reg         [31:0] r_sys_tmp97_float;
	reg         [31:0] r_sys_tmp98_float;
	reg         [31:0] r_sys_tmp99_float;
	reg         [31:0] r_sys_tmp100_float;
	reg         [31:0] r_sys_tmp101_float;
	reg         [31:0] r_sys_tmp102_float;
	reg         [31:0] r_sys_tmp103_float;
	reg         [31:0] r_sys_tmp104_float;
	reg         [31:0] r_sys_tmp105_float;
	reg         [31:0] r_sys_tmp106_float;
	reg         [31:0] r_sys_tmp107_float;
	reg         [31:0] r_sys_tmp108_float;
	reg         [31:0] r_sys_tmp109_float;
	reg         [31:0] r_sys_tmp110_float;
	reg         [31:0] r_sys_tmp111_float;
	reg         [31:0] r_sys_tmp112_float;
	reg         [31:0] r_sys_tmp113_float;
	reg         [31:0] r_sys_tmp114_float;
	reg         [31:0] r_sys_tmp115_float;
	reg         [31:0] r_sys_tmp116_float;
	reg         [31:0] r_sys_tmp117_float;
	reg         [31:0] r_sys_tmp118_float;
	reg         [31:0] r_sys_tmp119_float;
	reg         [31:0] r_sys_tmp120_float;
	reg         [31:0] r_sys_tmp121_float;
	reg         [31:0] r_sys_tmp122_float;
	reg         [31:0] r_sys_tmp123_float;
	reg         [31:0] r_sys_tmp124_float;
	reg         [31:0] r_sys_tmp125_float;
	reg         [31:0] r_sys_tmp126_float;
	reg         [31:0] r_sys_tmp127_float;
	reg         [31:0] r_sys_tmp128_float;
	reg         [31:0] r_sys_tmp129_float;
	reg         [31:0] r_sys_tmp130_float;
	reg         [31:0] r_sys_tmp131_float;
	reg         [31:0] r_sys_tmp132_float;
	reg         [31:0] r_sys_tmp133_float;
	reg         [31:0] r_sys_tmp134_float;
	reg         [31:0] r_sys_tmp135_float;
	reg         [31:0] r_sys_tmp136_float;
	reg         [31:0] r_sys_tmp137_float;
	reg         [31:0] r_sys_tmp138_float;
	reg         [31:0] r_sys_tmp139_float;
	reg         [31:0] r_sys_tmp140_float;
	reg         [31:0] r_sys_tmp141_float;
	reg         [31:0] r_sys_tmp142_float;
	reg         [31:0] r_sys_tmp143_float;
	reg         [31:0] r_sys_tmp144_float;
	reg         [31:0] r_sys_tmp145_float;
	reg         [31:0] r_sys_tmp146_float;
	reg         [31:0] r_sys_tmp147_float;
	reg         [31:0] r_sys_tmp148_float;
	reg         [31:0] r_sys_tmp149_float;
	reg         [31:0] r_sys_tmp150_float;
	reg         [31:0] r_sys_tmp151_float;
	reg         [31:0] r_sys_tmp152_float;
	reg         [31:0] r_sys_tmp153_float;
	reg         [31:0] r_sys_tmp154_float;
	reg         [31:0] r_sys_tmp155_float;
	reg         [31:0] r_sys_tmp156_float;
	reg         [31:0] r_sys_tmp157_float;
	reg         [31:0] r_sys_tmp158_float;
	reg         [31:0] r_sys_tmp159_float;
	reg         [31:0] r_sys_tmp160_float;
	reg         [31:0] r_sys_tmp161_float;
	reg         [31:0] r_sys_tmp162_float;
	reg         [31:0] r_sys_tmp163_float;
	reg         [31:0] r_sys_tmp164_float;
	reg         [31:0] r_sys_tmp165_float;
	reg         [31:0] r_sys_tmp166_float;
	reg         [31:0] r_sys_tmp167_float;
	reg         [31:0] r_sys_tmp168_float;
	reg         [31:0] r_sys_tmp169_float;
	reg         [31:0] r_sys_tmp170_float;
	reg         [31:0] r_sys_tmp171_float;
	reg         [31:0] r_sys_tmp172_float;
	reg         [31:0] r_sys_tmp173_float;
	reg         [31:0] r_sys_tmp174_float;
	reg         [31:0] r_sys_tmp175_float;
	reg         [31:0] r_sys_tmp176_float;
	reg         [31:0] r_sys_tmp177_float;
	reg         [31:0] r_sys_tmp178_float;
	reg         [31:0] r_sys_tmp179_float;
	reg         [31:0] r_sys_tmp180_float;
	reg         [31:0] r_sys_tmp181_float;
	reg         [31:0] r_sys_tmp182_float;
	reg         [31:0] r_sys_tmp183_float;
	reg         [31:0] r_sys_tmp184_float;
	reg         [31:0] r_sys_tmp185_float;
	reg         [31:0] r_sys_tmp186_float;
	reg         [31:0] r_sys_tmp187_float;
	reg         [31:0] r_sys_tmp188_float;
	reg         [31:0] r_sys_tmp189_float;
	reg         [31:0] r_sys_tmp190_float;
	reg         [31:0] r_sys_tmp191_float;
	reg         [31:0] r_sys_tmp192_float;
	reg         [31:0] r_sys_tmp193_float;
	reg         [31:0] r_sys_tmp194_float;
	reg         [31:0] r_sys_tmp195_float;
	reg         [31:0] r_sys_tmp196_float;
	reg         [31:0] r_sys_tmp197_float;
	reg         [31:0] r_sys_tmp198_float;
	reg         [31:0] r_sys_tmp199_float;
	reg         [31:0] r_sys_tmp200_float;
	reg         [31:0] r_sys_tmp201_float;
	reg         [31:0] r_sys_tmp202_float;
	reg         [31:0] r_sys_tmp203_float;
	reg         [31:0] r_sys_tmp204_float;
	reg         [31:0] r_sys_tmp205_float;
	reg         [31:0] r_sys_tmp206_float;
	reg         [31:0] r_sys_tmp207_float;
	reg         [31:0] r_sys_tmp208_float;
	reg         [31:0] r_sys_tmp209_float;
	reg         [31:0] r_sys_tmp210_float;
	reg         [31:0] r_sys_tmp211_float;
	reg         [31:0] r_sys_tmp212_float;
	reg         [31:0] r_sys_tmp213_float;
	reg         [31:0] r_sys_tmp214_float;
	reg         [31:0] r_sys_tmp215_float;
	reg         [31:0] r_sys_tmp216_float;
	reg         [31:0] r_sys_tmp217_float;
	reg         [31:0] r_sys_tmp218_float;
	reg         [31:0] r_sys_tmp219_float;
	reg         [31:0] r_sys_tmp220_float;
	reg         [31:0] r_sys_tmp221_float;
	reg         [31:0] r_sys_tmp222_float;
	reg         [31:0] r_sys_tmp223_float;
	reg         [31:0] r_sys_tmp224_float;
	reg         [31:0] r_sys_tmp225_float;
	reg         [31:0] r_sys_tmp226_float;
	reg         [31:0] r_sys_tmp227_float;
	reg         [31:0] r_sys_tmp228_float;
	reg         [31:0] r_sys_tmp229_float;
	reg         [31:0] r_sys_tmp230_float;
	reg         [31:0] r_sys_tmp231_float;
	reg         [31:0] r_sys_tmp232_float;
	reg         [31:0] r_sys_tmp233_float;
	reg         [31:0] r_sys_tmp234_float;
	reg         [31:0] r_sys_tmp235_float;
	reg         [31:0] r_sys_tmp236_float;
	reg         [31:0] r_sys_tmp237_float;
	reg         [31:0] r_sys_tmp238_float;
	reg         [31:0] r_sys_tmp239_float;
	reg         [31:0] r_sys_tmp240_float;
	reg         [31:0] r_sys_tmp241_float;
	reg         [31:0] r_sys_tmp242_float;
	reg         [31:0] r_sys_tmp243_float;
	reg         [31:0] r_sys_tmp244_float;
	reg         [31:0] r_sys_tmp245_float;
	reg         [31:0] r_sys_tmp246_float;
	reg         [31:0] r_sys_tmp247_float;
	reg         [31:0] r_sys_tmp248_float;
	reg         [31:0] r_sys_tmp249_float;
	reg         [31:0] r_sys_tmp250_float;
	reg         [31:0] r_sys_tmp251_float;
	reg         [31:0] r_sys_tmp252_float;
	reg         [31:0] r_sys_tmp253_float;
	reg         [31:0] r_sys_tmp254_float;
	reg         [31:0] r_sys_tmp255_float;
	reg         [31:0] r_sys_tmp256_float;
	reg         [31:0] r_sys_tmp257_float;
	reg         [31:0] r_sys_tmp258_float;
	reg         [31:0] r_sys_tmp259_float;
	reg         [31:0] r_sys_tmp260_float;
	reg         [31:0] r_sys_tmp261_float;
	reg         [31:0] r_sys_tmp262_float;
	reg         [31:0] r_sys_tmp263_float;
	reg         [31:0] r_sys_tmp264_float;
	reg         [31:0] r_sys_tmp265_float;
	reg         [31:0] r_sys_tmp266_float;
	reg         [31:0] r_sys_tmp267_float;
	reg         [31:0] r_sys_tmp268_float;
	reg         [31:0] r_sys_tmp269_float;
	reg         [31:0] r_sys_tmp270_float;
	reg         [31:0] r_sys_tmp271_float;
	reg         [31:0] r_sys_tmp272_float;
	reg         [31:0] r_sys_tmp273_float;
	reg         [31:0] r_sys_tmp274_float;
	reg         [31:0] r_sys_tmp275_float;
	reg         [31:0] r_sys_tmp276_float;
	reg         [31:0] r_sys_tmp277_float;
	reg         [31:0] r_sys_tmp278_float;
	reg         [31:0] r_sys_tmp279_float;
	reg         [31:0] r_sys_tmp280_float;
	reg         [31:0] r_sys_tmp281_float;
	reg         [31:0] r_sys_tmp282_float;
	reg         [31:0] r_sys_tmp283_float;
	reg         [31:0] r_sys_tmp284_float;
	reg         [31:0] r_sys_tmp285_float;
	reg         [31:0] r_sys_tmp286_float;
	reg         [31:0] r_sys_tmp287_float;
	reg         [31:0] r_sys_tmp288_float;
	reg         [31:0] r_sys_tmp289_float;
	reg         [31:0] r_sys_tmp290_float;
	reg         [31:0] r_sys_tmp291_float;
	reg         [31:0] r_sys_tmp292_float;
	reg         [31:0] r_sys_tmp293_float;
	reg         [31:0] r_sys_tmp294_float;
	reg         [31:0] r_sys_tmp295_float;
	reg         [31:0] r_sys_tmp296_float;
	reg         [31:0] r_sys_tmp297_float;
	reg         [31:0] r_sys_tmp298_float;
	reg         [31:0] r_sys_tmp299_float;
	reg         [31:0] r_sys_tmp300_float;
	reg         [31:0] r_sys_tmp301_float;
	reg         [31:0] r_sys_tmp302_float;
	reg         [31:0] r_sys_tmp303_float;
	reg         [31:0] r_sys_tmp304_float;
	reg         [31:0] r_sys_tmp305_float;
	reg         [31:0] r_sys_tmp306_float;
	reg         [31:0] r_sys_tmp307_float;
	reg         [31:0] r_sys_tmp308_float;
	reg         [31:0] r_sys_tmp309_float;
	reg         [31:0] r_sys_tmp310_float;
	reg         [31:0] r_sys_tmp311_float;
	reg         [31:0] r_sys_tmp312_float;
	reg         [31:0] r_sys_tmp313_float;
	reg         [31:0] r_sys_tmp314_float;
	reg         [31:0] r_sys_tmp315_float;
	reg         [31:0] r_sys_tmp316_float;
	reg         [31:0] r_sys_tmp317_float;
	reg         [31:0] r_sys_tmp318_float;
	reg         [31:0] r_sys_tmp319_float;
	reg         [31:0] r_sys_tmp320_float;
	reg         [31:0] r_sys_tmp321_float;
	reg         [31:0] r_sys_tmp322_float;
	reg         [31:0] r_sys_tmp323_float;
	reg         [31:0] r_sys_tmp324_float;
	reg         [31:0] r_sys_tmp325_float;
	reg         [31:0] r_sys_tmp326_float;
	reg         [31:0] r_sys_tmp327_float;
	reg         [31:0] r_sys_tmp328_float;
	reg         [31:0] r_sys_tmp329_float;
	reg         [31:0] r_sys_tmp330_float;
	reg         [31:0] r_sys_tmp331_float;
	reg         [31:0] r_sys_tmp332_float;
	reg         [31:0] r_sys_tmp333_float;
	reg         [31:0] r_sys_tmp334_float;
	reg         [31:0] r_sys_tmp335_float;
	reg         [31:0] r_sys_tmp336_float;
	reg         [31:0] r_sys_tmp337_float;
	reg         [31:0] r_sys_tmp338_float;
	reg         [31:0] r_sys_tmp339_float;
	reg         [31:0] r_sys_tmp340_float;
	reg         [31:0] r_sys_tmp341_float;
	reg         [31:0] r_sys_tmp342_float;
	reg         [31:0] r_sys_tmp343_float;
	reg         [31:0] r_sys_tmp344_float;
	reg         [31:0] r_sys_tmp345_float;
	reg         [31:0] r_sys_tmp346_float;
	reg         [31:0] r_sys_tmp347_float;
	reg         [31:0] r_sys_tmp348_float;
	wire signed [31:0] w_sys_tmp1;
	wire               w_sys_tmp3;
	wire               w_sys_tmp4;
	wire signed [31:0] w_sys_tmp5;
	wire               w_sys_tmp6;
	wire               w_sys_tmp7;
	wire signed [31:0] w_sys_tmp10;
	wire signed [31:0] w_sys_tmp11;
	wire signed [31:0] w_sys_tmp12;
	wire        [31:0] w_sys_tmp13;
	wire signed [31:0] w_sys_tmp14;
	wire               w_sys_tmp51;
	wire               w_sys_tmp52;
	wire signed [31:0] w_sys_tmp53;
	wire               w_sys_tmp54;
	wire               w_sys_tmp55;
	wire signed [31:0] w_sys_tmp58;
	wire signed [31:0] w_sys_tmp59;
	wire        [31:0] w_sys_tmp60;
	wire signed [31:0] w_sys_tmp62;
	wire signed [31:0] w_sys_tmp63;
	wire        [31:0] w_sys_tmp64;
	wire signed [31:0] w_sys_tmp66;
	wire signed [31:0] w_sys_tmp67;
	wire        [31:0] w_sys_tmp69;
	wire signed [31:0] w_sys_tmp71;
	wire signed [31:0] w_sys_tmp72;
	wire signed [31:0] w_sys_tmp75;
	wire signed [31:0] w_sys_tmp76;
	wire signed [31:0] w_sys_tmp77;
	wire signed [31:0] w_sys_tmp78;
	wire               w_sys_tmp211;
	wire               w_sys_tmp212;
	wire signed [31:0] w_sys_tmp213;
	wire signed [31:0] w_sys_tmp216;
	wire signed [31:0] w_sys_tmp217;
	wire        [31:0] w_sys_tmp218;
	wire signed [31:0] w_sys_tmp222;
	wire signed [31:0] w_sys_tmp223;
	wire signed [31:0] w_sys_tmp228;
	wire signed [31:0] w_sys_tmp229;
	wire signed [31:0] w_sys_tmp234;
	wire signed [31:0] w_sys_tmp235;
	wire signed [31:0] w_sys_tmp240;
	wire signed [31:0] w_sys_tmp241;
	wire signed [31:0] w_sys_tmp246;
	wire signed [31:0] w_sys_tmp247;
	wire signed [31:0] w_sys_tmp252;
	wire signed [31:0] w_sys_tmp253;
	wire signed [31:0] w_sys_tmp258;
	wire signed [31:0] w_sys_tmp259;
	wire signed [31:0] w_sys_tmp264;
	wire signed [31:0] w_sys_tmp265;
	wire signed [31:0] w_sys_tmp270;
	wire signed [31:0] w_sys_tmp271;
	wire signed [31:0] w_sys_tmp276;
	wire signed [31:0] w_sys_tmp277;
	wire signed [31:0] w_sys_tmp282;
	wire signed [31:0] w_sys_tmp283;
	wire signed [31:0] w_sys_tmp288;
	wire signed [31:0] w_sys_tmp289;
	wire signed [31:0] w_sys_tmp294;
	wire signed [31:0] w_sys_tmp295;
	wire signed [31:0] w_sys_tmp300;
	wire signed [31:0] w_sys_tmp301;
	wire signed [31:0] w_sys_tmp306;
	wire signed [31:0] w_sys_tmp307;
	wire signed [31:0] w_sys_tmp312;
	wire signed [31:0] w_sys_tmp313;
	wire signed [31:0] w_sys_tmp318;
	wire signed [31:0] w_sys_tmp319;
	wire signed [31:0] w_sys_tmp324;
	wire signed [31:0] w_sys_tmp325;
	wire signed [31:0] w_sys_tmp330;
	wire signed [31:0] w_sys_tmp331;
	wire signed [31:0] w_sys_tmp336;
	wire signed [31:0] w_sys_tmp337;
	wire signed [31:0] w_sys_tmp342;
	wire signed [31:0] w_sys_tmp343;
	wire signed [31:0] w_sys_tmp348;
	wire signed [31:0] w_sys_tmp349;
	wire signed [31:0] w_sys_tmp354;
	wire signed [31:0] w_sys_tmp355;
	wire signed [31:0] w_sys_tmp360;
	wire signed [31:0] w_sys_tmp361;
	wire signed [31:0] w_sys_tmp366;
	wire signed [31:0] w_sys_tmp367;
	wire signed [31:0] w_sys_tmp372;
	wire signed [31:0] w_sys_tmp373;
	wire signed [31:0] w_sys_tmp378;
	wire signed [31:0] w_sys_tmp379;
	wire signed [31:0] w_sys_tmp384;
	wire signed [31:0] w_sys_tmp385;
	wire signed [31:0] w_sys_tmp390;
	wire signed [31:0] w_sys_tmp391;
	wire signed [31:0] w_sys_tmp396;
	wire signed [31:0] w_sys_tmp397;
	wire signed [31:0] w_sys_tmp402;
	wire signed [31:0] w_sys_tmp403;
	wire signed [31:0] w_sys_tmp408;
	wire signed [31:0] w_sys_tmp409;
	wire signed [31:0] w_sys_tmp426;
	wire signed [31:0] w_sys_tmp427;
	wire signed [31:0] w_sys_tmp432;
	wire signed [31:0] w_sys_tmp433;
	wire signed [31:0] w_sys_tmp438;
	wire signed [31:0] w_sys_tmp439;
	wire signed [31:0] w_sys_tmp444;
	wire signed [31:0] w_sys_tmp445;
	wire signed [31:0] w_sys_tmp450;
	wire signed [31:0] w_sys_tmp451;
	wire signed [31:0] w_sys_tmp456;
	wire signed [31:0] w_sys_tmp457;
	wire signed [31:0] w_sys_tmp462;
	wire signed [31:0] w_sys_tmp463;
	wire signed [31:0] w_sys_tmp468;
	wire signed [31:0] w_sys_tmp469;
	wire signed [31:0] w_sys_tmp474;
	wire signed [31:0] w_sys_tmp475;
	wire signed [31:0] w_sys_tmp480;
	wire signed [31:0] w_sys_tmp481;
	wire signed [31:0] w_sys_tmp486;
	wire signed [31:0] w_sys_tmp487;
	wire signed [31:0] w_sys_tmp492;
	wire signed [31:0] w_sys_tmp493;
	wire signed [31:0] w_sys_tmp498;
	wire signed [31:0] w_sys_tmp499;
	wire signed [31:0] w_sys_tmp504;
	wire signed [31:0] w_sys_tmp505;
	wire signed [31:0] w_sys_tmp510;
	wire signed [31:0] w_sys_tmp511;
	wire signed [31:0] w_sys_tmp516;
	wire signed [31:0] w_sys_tmp517;
	wire signed [31:0] w_sys_tmp522;
	wire signed [31:0] w_sys_tmp523;
	wire signed [31:0] w_sys_tmp528;
	wire signed [31:0] w_sys_tmp529;
	wire signed [31:0] w_sys_tmp534;
	wire signed [31:0] w_sys_tmp535;
	wire signed [31:0] w_sys_tmp540;
	wire signed [31:0] w_sys_tmp541;
	wire signed [31:0] w_sys_tmp546;
	wire signed [31:0] w_sys_tmp547;
	wire signed [31:0] w_sys_tmp552;
	wire signed [31:0] w_sys_tmp553;
	wire signed [31:0] w_sys_tmp558;
	wire signed [31:0] w_sys_tmp559;
	wire signed [31:0] w_sys_tmp564;
	wire signed [31:0] w_sys_tmp565;
	wire signed [31:0] w_sys_tmp570;
	wire signed [31:0] w_sys_tmp571;
	wire signed [31:0] w_sys_tmp576;
	wire signed [31:0] w_sys_tmp577;
	wire signed [31:0] w_sys_tmp582;
	wire signed [31:0] w_sys_tmp583;
	wire signed [31:0] w_sys_tmp588;
	wire signed [31:0] w_sys_tmp589;
	wire signed [31:0] w_sys_tmp594;
	wire signed [31:0] w_sys_tmp595;
	wire signed [31:0] w_sys_tmp600;
	wire signed [31:0] w_sys_tmp601;
	wire signed [31:0] w_sys_tmp606;
	wire signed [31:0] w_sys_tmp607;
	wire signed [31:0] w_sys_tmp612;
	wire signed [31:0] w_sys_tmp613;
	wire signed [31:0] w_sys_tmp630;
	wire signed [31:0] w_sys_tmp631;
	wire signed [31:0] w_sys_tmp636;
	wire signed [31:0] w_sys_tmp637;
	wire signed [31:0] w_sys_tmp642;
	wire signed [31:0] w_sys_tmp643;
	wire signed [31:0] w_sys_tmp648;
	wire signed [31:0] w_sys_tmp649;
	wire signed [31:0] w_sys_tmp654;
	wire signed [31:0] w_sys_tmp655;
	wire signed [31:0] w_sys_tmp660;
	wire signed [31:0] w_sys_tmp661;
	wire signed [31:0] w_sys_tmp666;
	wire signed [31:0] w_sys_tmp667;
	wire signed [31:0] w_sys_tmp672;
	wire signed [31:0] w_sys_tmp673;
	wire signed [31:0] w_sys_tmp678;
	wire signed [31:0] w_sys_tmp679;
	wire signed [31:0] w_sys_tmp684;
	wire signed [31:0] w_sys_tmp685;
	wire signed [31:0] w_sys_tmp690;
	wire signed [31:0] w_sys_tmp691;
	wire signed [31:0] w_sys_tmp696;
	wire signed [31:0] w_sys_tmp697;
	wire signed [31:0] w_sys_tmp702;
	wire signed [31:0] w_sys_tmp703;
	wire signed [31:0] w_sys_tmp708;
	wire signed [31:0] w_sys_tmp709;
	wire signed [31:0] w_sys_tmp714;
	wire signed [31:0] w_sys_tmp715;
	wire signed [31:0] w_sys_tmp720;
	wire signed [31:0] w_sys_tmp721;
	wire signed [31:0] w_sys_tmp726;
	wire signed [31:0] w_sys_tmp727;
	wire signed [31:0] w_sys_tmp732;
	wire signed [31:0] w_sys_tmp733;
	wire signed [31:0] w_sys_tmp738;
	wire signed [31:0] w_sys_tmp739;
	wire signed [31:0] w_sys_tmp744;
	wire signed [31:0] w_sys_tmp745;
	wire signed [31:0] w_sys_tmp750;
	wire signed [31:0] w_sys_tmp751;
	wire signed [31:0] w_sys_tmp756;
	wire signed [31:0] w_sys_tmp757;
	wire signed [31:0] w_sys_tmp762;
	wire signed [31:0] w_sys_tmp763;
	wire signed [31:0] w_sys_tmp768;
	wire signed [31:0] w_sys_tmp769;
	wire signed [31:0] w_sys_tmp774;
	wire signed [31:0] w_sys_tmp775;
	wire signed [31:0] w_sys_tmp780;
	wire signed [31:0] w_sys_tmp781;
	wire signed [31:0] w_sys_tmp786;
	wire signed [31:0] w_sys_tmp787;
	wire signed [31:0] w_sys_tmp792;
	wire signed [31:0] w_sys_tmp793;
	wire signed [31:0] w_sys_tmp798;
	wire signed [31:0] w_sys_tmp799;
	wire signed [31:0] w_sys_tmp804;
	wire signed [31:0] w_sys_tmp805;
	wire signed [31:0] w_sys_tmp810;
	wire signed [31:0] w_sys_tmp811;
	wire signed [31:0] w_sys_tmp816;
	wire signed [31:0] w_sys_tmp817;
	wire signed [31:0] w_sys_tmp834;
	wire signed [31:0] w_sys_tmp835;
	wire signed [31:0] w_sys_tmp840;
	wire signed [31:0] w_sys_tmp841;
	wire signed [31:0] w_sys_tmp846;
	wire signed [31:0] w_sys_tmp847;
	wire signed [31:0] w_sys_tmp852;
	wire signed [31:0] w_sys_tmp853;
	wire signed [31:0] w_sys_tmp858;
	wire signed [31:0] w_sys_tmp859;
	wire signed [31:0] w_sys_tmp864;
	wire signed [31:0] w_sys_tmp865;
	wire signed [31:0] w_sys_tmp870;
	wire signed [31:0] w_sys_tmp871;
	wire signed [31:0] w_sys_tmp876;
	wire signed [31:0] w_sys_tmp877;
	wire signed [31:0] w_sys_tmp882;
	wire signed [31:0] w_sys_tmp883;
	wire signed [31:0] w_sys_tmp888;
	wire signed [31:0] w_sys_tmp889;
	wire signed [31:0] w_sys_tmp894;
	wire signed [31:0] w_sys_tmp895;
	wire signed [31:0] w_sys_tmp900;
	wire signed [31:0] w_sys_tmp901;
	wire signed [31:0] w_sys_tmp906;
	wire signed [31:0] w_sys_tmp907;
	wire signed [31:0] w_sys_tmp912;
	wire signed [31:0] w_sys_tmp913;
	wire signed [31:0] w_sys_tmp918;
	wire signed [31:0] w_sys_tmp919;
	wire signed [31:0] w_sys_tmp924;
	wire signed [31:0] w_sys_tmp925;
	wire signed [31:0] w_sys_tmp930;
	wire signed [31:0] w_sys_tmp931;
	wire signed [31:0] w_sys_tmp936;
	wire signed [31:0] w_sys_tmp937;
	wire signed [31:0] w_sys_tmp942;
	wire signed [31:0] w_sys_tmp943;
	wire signed [31:0] w_sys_tmp948;
	wire signed [31:0] w_sys_tmp949;
	wire signed [31:0] w_sys_tmp954;
	wire signed [31:0] w_sys_tmp955;
	wire signed [31:0] w_sys_tmp960;
	wire signed [31:0] w_sys_tmp961;
	wire signed [31:0] w_sys_tmp966;
	wire signed [31:0] w_sys_tmp967;
	wire signed [31:0] w_sys_tmp972;
	wire signed [31:0] w_sys_tmp973;
	wire signed [31:0] w_sys_tmp978;
	wire signed [31:0] w_sys_tmp979;
	wire signed [31:0] w_sys_tmp984;
	wire signed [31:0] w_sys_tmp985;
	wire signed [31:0] w_sys_tmp990;
	wire signed [31:0] w_sys_tmp991;
	wire signed [31:0] w_sys_tmp996;
	wire signed [31:0] w_sys_tmp997;
	wire signed [31:0] w_sys_tmp1002;
	wire signed [31:0] w_sys_tmp1003;
	wire signed [31:0] w_sys_tmp1008;
	wire signed [31:0] w_sys_tmp1009;
	wire signed [31:0] w_sys_tmp1014;
	wire signed [31:0] w_sys_tmp1015;
	wire signed [31:0] w_sys_tmp1020;
	wire signed [31:0] w_sys_tmp1021;
	wire signed [31:0] w_sys_tmp1025;
	wire signed [31:0] w_sys_tmp1026;
	wire               w_sys_tmp1027;
	wire               w_sys_tmp1028;
	wire signed [31:0] w_sys_tmp1029;
	wire signed [31:0] w_sys_tmp1032;
	wire signed [31:0] w_sys_tmp1033;
	wire        [31:0] w_sys_tmp1034;
	wire signed [31:0] w_sys_tmp1038;
	wire signed [31:0] w_sys_tmp1039;
	wire signed [31:0] w_sys_tmp1044;
	wire signed [31:0] w_sys_tmp1045;
	wire signed [31:0] w_sys_tmp1050;
	wire signed [31:0] w_sys_tmp1051;
	wire signed [31:0] w_sys_tmp1056;
	wire signed [31:0] w_sys_tmp1057;
	wire signed [31:0] w_sys_tmp1062;
	wire signed [31:0] w_sys_tmp1063;
	wire signed [31:0] w_sys_tmp1068;
	wire signed [31:0] w_sys_tmp1069;
	wire signed [31:0] w_sys_tmp1074;
	wire signed [31:0] w_sys_tmp1075;
	wire signed [31:0] w_sys_tmp1080;
	wire signed [31:0] w_sys_tmp1081;
	wire signed [31:0] w_sys_tmp1086;
	wire signed [31:0] w_sys_tmp1087;
	wire signed [31:0] w_sys_tmp1092;
	wire signed [31:0] w_sys_tmp1093;
	wire signed [31:0] w_sys_tmp1098;
	wire signed [31:0] w_sys_tmp1099;
	wire signed [31:0] w_sys_tmp1104;
	wire signed [31:0] w_sys_tmp1105;
	wire signed [31:0] w_sys_tmp1110;
	wire signed [31:0] w_sys_tmp1111;
	wire signed [31:0] w_sys_tmp1116;
	wire signed [31:0] w_sys_tmp1117;
	wire signed [31:0] w_sys_tmp1122;
	wire signed [31:0] w_sys_tmp1123;
	wire signed [31:0] w_sys_tmp1128;
	wire signed [31:0] w_sys_tmp1129;
	wire signed [31:0] w_sys_tmp1134;
	wire signed [31:0] w_sys_tmp1135;
	wire signed [31:0] w_sys_tmp1140;
	wire signed [31:0] w_sys_tmp1141;
	wire signed [31:0] w_sys_tmp1146;
	wire signed [31:0] w_sys_tmp1147;
	wire signed [31:0] w_sys_tmp1152;
	wire signed [31:0] w_sys_tmp1153;
	wire signed [31:0] w_sys_tmp1158;
	wire signed [31:0] w_sys_tmp1159;
	wire signed [31:0] w_sys_tmp1164;
	wire signed [31:0] w_sys_tmp1165;
	wire signed [31:0] w_sys_tmp1170;
	wire signed [31:0] w_sys_tmp1171;
	wire signed [31:0] w_sys_tmp1176;
	wire signed [31:0] w_sys_tmp1177;
	wire signed [31:0] w_sys_tmp1182;
	wire signed [31:0] w_sys_tmp1183;
	wire signed [31:0] w_sys_tmp1188;
	wire signed [31:0] w_sys_tmp1189;
	wire signed [31:0] w_sys_tmp1194;
	wire signed [31:0] w_sys_tmp1195;
	wire signed [31:0] w_sys_tmp1200;
	wire signed [31:0] w_sys_tmp1201;
	wire signed [31:0] w_sys_tmp1206;
	wire signed [31:0] w_sys_tmp1207;
	wire signed [31:0] w_sys_tmp1212;
	wire signed [31:0] w_sys_tmp1213;
	wire signed [31:0] w_sys_tmp1218;
	wire signed [31:0] w_sys_tmp1219;
	wire signed [31:0] w_sys_tmp1224;
	wire signed [31:0] w_sys_tmp1225;
	wire signed [31:0] w_sys_tmp1242;
	wire signed [31:0] w_sys_tmp1243;
	wire signed [31:0] w_sys_tmp1248;
	wire signed [31:0] w_sys_tmp1249;
	wire signed [31:0] w_sys_tmp1254;
	wire signed [31:0] w_sys_tmp1255;
	wire signed [31:0] w_sys_tmp1260;
	wire signed [31:0] w_sys_tmp1261;
	wire signed [31:0] w_sys_tmp1266;
	wire signed [31:0] w_sys_tmp1267;
	wire signed [31:0] w_sys_tmp1272;
	wire signed [31:0] w_sys_tmp1273;
	wire signed [31:0] w_sys_tmp1278;
	wire signed [31:0] w_sys_tmp1279;
	wire signed [31:0] w_sys_tmp1284;
	wire signed [31:0] w_sys_tmp1285;
	wire signed [31:0] w_sys_tmp1290;
	wire signed [31:0] w_sys_tmp1291;
	wire signed [31:0] w_sys_tmp1296;
	wire signed [31:0] w_sys_tmp1297;
	wire signed [31:0] w_sys_tmp1302;
	wire signed [31:0] w_sys_tmp1303;
	wire signed [31:0] w_sys_tmp1308;
	wire signed [31:0] w_sys_tmp1309;
	wire signed [31:0] w_sys_tmp1314;
	wire signed [31:0] w_sys_tmp1315;
	wire signed [31:0] w_sys_tmp1320;
	wire signed [31:0] w_sys_tmp1321;
	wire signed [31:0] w_sys_tmp1326;
	wire signed [31:0] w_sys_tmp1327;
	wire signed [31:0] w_sys_tmp1332;
	wire signed [31:0] w_sys_tmp1333;
	wire signed [31:0] w_sys_tmp1338;
	wire signed [31:0] w_sys_tmp1339;
	wire signed [31:0] w_sys_tmp1344;
	wire signed [31:0] w_sys_tmp1345;
	wire signed [31:0] w_sys_tmp1350;
	wire signed [31:0] w_sys_tmp1351;
	wire signed [31:0] w_sys_tmp1356;
	wire signed [31:0] w_sys_tmp1357;
	wire signed [31:0] w_sys_tmp1362;
	wire signed [31:0] w_sys_tmp1363;
	wire signed [31:0] w_sys_tmp1368;
	wire signed [31:0] w_sys_tmp1369;
	wire signed [31:0] w_sys_tmp1374;
	wire signed [31:0] w_sys_tmp1375;
	wire signed [31:0] w_sys_tmp1380;
	wire signed [31:0] w_sys_tmp1381;
	wire signed [31:0] w_sys_tmp1386;
	wire signed [31:0] w_sys_tmp1387;
	wire signed [31:0] w_sys_tmp1392;
	wire signed [31:0] w_sys_tmp1393;
	wire signed [31:0] w_sys_tmp1398;
	wire signed [31:0] w_sys_tmp1399;
	wire signed [31:0] w_sys_tmp1404;
	wire signed [31:0] w_sys_tmp1405;
	wire signed [31:0] w_sys_tmp1410;
	wire signed [31:0] w_sys_tmp1411;
	wire signed [31:0] w_sys_tmp1416;
	wire signed [31:0] w_sys_tmp1417;
	wire signed [31:0] w_sys_tmp1422;
	wire signed [31:0] w_sys_tmp1423;
	wire signed [31:0] w_sys_tmp1428;
	wire signed [31:0] w_sys_tmp1429;
	wire signed [31:0] w_sys_tmp1446;
	wire signed [31:0] w_sys_tmp1447;
	wire signed [31:0] w_sys_tmp1452;
	wire signed [31:0] w_sys_tmp1453;
	wire signed [31:0] w_sys_tmp1458;
	wire signed [31:0] w_sys_tmp1459;
	wire signed [31:0] w_sys_tmp1464;
	wire signed [31:0] w_sys_tmp1465;
	wire signed [31:0] w_sys_tmp1470;
	wire signed [31:0] w_sys_tmp1471;
	wire signed [31:0] w_sys_tmp1476;
	wire signed [31:0] w_sys_tmp1477;
	wire signed [31:0] w_sys_tmp1482;
	wire signed [31:0] w_sys_tmp1483;
	wire signed [31:0] w_sys_tmp1488;
	wire signed [31:0] w_sys_tmp1489;
	wire signed [31:0] w_sys_tmp1494;
	wire signed [31:0] w_sys_tmp1495;
	wire signed [31:0] w_sys_tmp1500;
	wire signed [31:0] w_sys_tmp1501;
	wire signed [31:0] w_sys_tmp1506;
	wire signed [31:0] w_sys_tmp1507;
	wire signed [31:0] w_sys_tmp1512;
	wire signed [31:0] w_sys_tmp1513;
	wire signed [31:0] w_sys_tmp1518;
	wire signed [31:0] w_sys_tmp1519;
	wire signed [31:0] w_sys_tmp1524;
	wire signed [31:0] w_sys_tmp1525;
	wire signed [31:0] w_sys_tmp1530;
	wire signed [31:0] w_sys_tmp1531;
	wire signed [31:0] w_sys_tmp1536;
	wire signed [31:0] w_sys_tmp1537;
	wire signed [31:0] w_sys_tmp1542;
	wire signed [31:0] w_sys_tmp1543;
	wire signed [31:0] w_sys_tmp1548;
	wire signed [31:0] w_sys_tmp1549;
	wire signed [31:0] w_sys_tmp1554;
	wire signed [31:0] w_sys_tmp1555;
	wire signed [31:0] w_sys_tmp1560;
	wire signed [31:0] w_sys_tmp1561;
	wire signed [31:0] w_sys_tmp1566;
	wire signed [31:0] w_sys_tmp1567;
	wire signed [31:0] w_sys_tmp1572;
	wire signed [31:0] w_sys_tmp1573;
	wire signed [31:0] w_sys_tmp1578;
	wire signed [31:0] w_sys_tmp1579;
	wire signed [31:0] w_sys_tmp1584;
	wire signed [31:0] w_sys_tmp1585;
	wire signed [31:0] w_sys_tmp1590;
	wire signed [31:0] w_sys_tmp1591;
	wire signed [31:0] w_sys_tmp1596;
	wire signed [31:0] w_sys_tmp1597;
	wire signed [31:0] w_sys_tmp1602;
	wire signed [31:0] w_sys_tmp1603;
	wire signed [31:0] w_sys_tmp1608;
	wire signed [31:0] w_sys_tmp1609;
	wire signed [31:0] w_sys_tmp1614;
	wire signed [31:0] w_sys_tmp1615;
	wire signed [31:0] w_sys_tmp1620;
	wire signed [31:0] w_sys_tmp1621;
	wire signed [31:0] w_sys_tmp1626;
	wire signed [31:0] w_sys_tmp1627;
	wire signed [31:0] w_sys_tmp1632;
	wire signed [31:0] w_sys_tmp1633;
	wire signed [31:0] w_sys_tmp1650;
	wire signed [31:0] w_sys_tmp1651;
	wire signed [31:0] w_sys_tmp1656;
	wire signed [31:0] w_sys_tmp1657;
	wire signed [31:0] w_sys_tmp1662;
	wire signed [31:0] w_sys_tmp1663;
	wire signed [31:0] w_sys_tmp1668;
	wire signed [31:0] w_sys_tmp1669;
	wire signed [31:0] w_sys_tmp1674;
	wire signed [31:0] w_sys_tmp1675;
	wire signed [31:0] w_sys_tmp1680;
	wire signed [31:0] w_sys_tmp1681;
	wire signed [31:0] w_sys_tmp1686;
	wire signed [31:0] w_sys_tmp1687;
	wire signed [31:0] w_sys_tmp1692;
	wire signed [31:0] w_sys_tmp1693;
	wire signed [31:0] w_sys_tmp1698;
	wire signed [31:0] w_sys_tmp1699;
	wire signed [31:0] w_sys_tmp1704;
	wire signed [31:0] w_sys_tmp1705;
	wire signed [31:0] w_sys_tmp1710;
	wire signed [31:0] w_sys_tmp1711;
	wire signed [31:0] w_sys_tmp1716;
	wire signed [31:0] w_sys_tmp1717;
	wire signed [31:0] w_sys_tmp1722;
	wire signed [31:0] w_sys_tmp1723;
	wire signed [31:0] w_sys_tmp1728;
	wire signed [31:0] w_sys_tmp1729;
	wire signed [31:0] w_sys_tmp1734;
	wire signed [31:0] w_sys_tmp1735;
	wire signed [31:0] w_sys_tmp1740;
	wire signed [31:0] w_sys_tmp1741;
	wire signed [31:0] w_sys_tmp1746;
	wire signed [31:0] w_sys_tmp1747;
	wire signed [31:0] w_sys_tmp1752;
	wire signed [31:0] w_sys_tmp1753;
	wire signed [31:0] w_sys_tmp1758;
	wire signed [31:0] w_sys_tmp1759;
	wire signed [31:0] w_sys_tmp1764;
	wire signed [31:0] w_sys_tmp1765;
	wire signed [31:0] w_sys_tmp1770;
	wire signed [31:0] w_sys_tmp1771;
	wire signed [31:0] w_sys_tmp1776;
	wire signed [31:0] w_sys_tmp1777;
	wire signed [31:0] w_sys_tmp1782;
	wire signed [31:0] w_sys_tmp1783;
	wire signed [31:0] w_sys_tmp1788;
	wire signed [31:0] w_sys_tmp1789;
	wire signed [31:0] w_sys_tmp1794;
	wire signed [31:0] w_sys_tmp1795;
	wire signed [31:0] w_sys_tmp1800;
	wire signed [31:0] w_sys_tmp1801;
	wire signed [31:0] w_sys_tmp1806;
	wire signed [31:0] w_sys_tmp1807;
	wire signed [31:0] w_sys_tmp1812;
	wire signed [31:0] w_sys_tmp1813;
	wire signed [31:0] w_sys_tmp1818;
	wire signed [31:0] w_sys_tmp1819;
	wire signed [31:0] w_sys_tmp1824;
	wire signed [31:0] w_sys_tmp1825;
	wire signed [31:0] w_sys_tmp1830;
	wire signed [31:0] w_sys_tmp1831;
	wire signed [31:0] w_sys_tmp1836;
	wire signed [31:0] w_sys_tmp1837;
	wire signed [31:0] w_sys_tmp1842;
	wire signed [31:0] w_sys_tmp1843;
	wire signed [31:0] w_sys_tmp1848;
	wire signed [31:0] w_sys_tmp1849;
	wire signed [31:0] w_sys_tmp1854;
	wire signed [31:0] w_sys_tmp1855;
	wire signed [31:0] w_sys_tmp1860;
	wire signed [31:0] w_sys_tmp1861;
	wire signed [31:0] w_sys_tmp1866;
	wire signed [31:0] w_sys_tmp1867;
	wire signed [31:0] w_sys_tmp1872;
	wire signed [31:0] w_sys_tmp1873;
	wire signed [31:0] w_sys_tmp1878;
	wire signed [31:0] w_sys_tmp1879;
	wire signed [31:0] w_sys_tmp1884;
	wire signed [31:0] w_sys_tmp1885;
	wire signed [31:0] w_sys_tmp1890;
	wire signed [31:0] w_sys_tmp1891;
	wire signed [31:0] w_sys_tmp1896;
	wire signed [31:0] w_sys_tmp1897;
	wire signed [31:0] w_sys_tmp1902;
	wire signed [31:0] w_sys_tmp1903;
	wire signed [31:0] w_sys_tmp1908;
	wire signed [31:0] w_sys_tmp1909;
	wire signed [31:0] w_sys_tmp1914;
	wire signed [31:0] w_sys_tmp1915;
	wire signed [31:0] w_sys_tmp1920;
	wire signed [31:0] w_sys_tmp1921;
	wire signed [31:0] w_sys_tmp1926;
	wire signed [31:0] w_sys_tmp1927;
	wire signed [31:0] w_sys_tmp1932;
	wire signed [31:0] w_sys_tmp1933;
	wire signed [31:0] w_sys_tmp1938;
	wire signed [31:0] w_sys_tmp1939;
	wire signed [31:0] w_sys_tmp1944;
	wire signed [31:0] w_sys_tmp1945;
	wire signed [31:0] w_sys_tmp1950;
	wire signed [31:0] w_sys_tmp1951;
	wire signed [31:0] w_sys_tmp1956;
	wire signed [31:0] w_sys_tmp1957;
	wire signed [31:0] w_sys_tmp1962;
	wire signed [31:0] w_sys_tmp1963;
	wire signed [31:0] w_sys_tmp1968;
	wire signed [31:0] w_sys_tmp1969;
	wire signed [31:0] w_sys_tmp1974;
	wire signed [31:0] w_sys_tmp1975;
	wire signed [31:0] w_sys_tmp1980;
	wire signed [31:0] w_sys_tmp1981;
	wire signed [31:0] w_sys_tmp1986;
	wire signed [31:0] w_sys_tmp1987;
	wire signed [31:0] w_sys_tmp1992;
	wire signed [31:0] w_sys_tmp1993;
	wire signed [31:0] w_sys_tmp1998;
	wire signed [31:0] w_sys_tmp1999;
	wire signed [31:0] w_sys_tmp2004;
	wire signed [31:0] w_sys_tmp2005;
	wire signed [31:0] w_sys_tmp2010;
	wire signed [31:0] w_sys_tmp2011;
	wire signed [31:0] w_sys_tmp2016;
	wire signed [31:0] w_sys_tmp2017;
	wire signed [31:0] w_sys_tmp2022;
	wire signed [31:0] w_sys_tmp2023;
	wire signed [31:0] w_sys_tmp2028;
	wire signed [31:0] w_sys_tmp2029;
	wire signed [31:0] w_sys_tmp2034;
	wire signed [31:0] w_sys_tmp2035;
	wire signed [31:0] w_sys_tmp2052;
	wire signed [31:0] w_sys_tmp2053;
	wire signed [31:0] w_sys_tmp2058;
	wire signed [31:0] w_sys_tmp2059;
	wire signed [31:0] w_sys_tmp2064;
	wire signed [31:0] w_sys_tmp2065;
	wire signed [31:0] w_sys_tmp2070;
	wire signed [31:0] w_sys_tmp2071;
	wire signed [31:0] w_sys_tmp2076;
	wire signed [31:0] w_sys_tmp2077;
	wire signed [31:0] w_sys_tmp2082;
	wire signed [31:0] w_sys_tmp2083;
	wire signed [31:0] w_sys_tmp2088;
	wire signed [31:0] w_sys_tmp2089;
	wire signed [31:0] w_sys_tmp2094;
	wire signed [31:0] w_sys_tmp2095;
	wire signed [31:0] w_sys_tmp2100;
	wire signed [31:0] w_sys_tmp2101;
	wire signed [31:0] w_sys_tmp2106;
	wire signed [31:0] w_sys_tmp2107;
	wire signed [31:0] w_sys_tmp2112;
	wire signed [31:0] w_sys_tmp2113;
	wire signed [31:0] w_sys_tmp2118;
	wire signed [31:0] w_sys_tmp2119;
	wire signed [31:0] w_sys_tmp2124;
	wire signed [31:0] w_sys_tmp2125;
	wire signed [31:0] w_sys_tmp2130;
	wire signed [31:0] w_sys_tmp2131;
	wire signed [31:0] w_sys_tmp2136;
	wire signed [31:0] w_sys_tmp2137;
	wire signed [31:0] w_sys_tmp2142;
	wire signed [31:0] w_sys_tmp2143;
	wire signed [31:0] w_sys_tmp2148;
	wire signed [31:0] w_sys_tmp2149;
	wire signed [31:0] w_sys_tmp2154;
	wire signed [31:0] w_sys_tmp2155;
	wire signed [31:0] w_sys_tmp2160;
	wire signed [31:0] w_sys_tmp2161;
	wire signed [31:0] w_sys_tmp2166;
	wire signed [31:0] w_sys_tmp2167;
	wire signed [31:0] w_sys_tmp2172;
	wire signed [31:0] w_sys_tmp2173;
	wire signed [31:0] w_sys_tmp2178;
	wire signed [31:0] w_sys_tmp2179;
	wire signed [31:0] w_sys_tmp2184;
	wire signed [31:0] w_sys_tmp2185;
	wire signed [31:0] w_sys_tmp2190;
	wire signed [31:0] w_sys_tmp2191;
	wire signed [31:0] w_sys_tmp2196;
	wire signed [31:0] w_sys_tmp2197;
	wire signed [31:0] w_sys_tmp2202;
	wire signed [31:0] w_sys_tmp2203;
	wire signed [31:0] w_sys_tmp2208;
	wire signed [31:0] w_sys_tmp2209;
	wire signed [31:0] w_sys_tmp2214;
	wire signed [31:0] w_sys_tmp2215;
	wire signed [31:0] w_sys_tmp2220;
	wire signed [31:0] w_sys_tmp2221;
	wire signed [31:0] w_sys_tmp2226;
	wire signed [31:0] w_sys_tmp2227;
	wire signed [31:0] w_sys_tmp2232;
	wire signed [31:0] w_sys_tmp2233;
	wire signed [31:0] w_sys_tmp2238;
	wire signed [31:0] w_sys_tmp2239;
	wire signed [31:0] w_sys_tmp2256;
	wire signed [31:0] w_sys_tmp2257;
	wire signed [31:0] w_sys_tmp2262;
	wire signed [31:0] w_sys_tmp2263;
	wire signed [31:0] w_sys_tmp2268;
	wire signed [31:0] w_sys_tmp2269;
	wire signed [31:0] w_sys_tmp2274;
	wire signed [31:0] w_sys_tmp2275;
	wire signed [31:0] w_sys_tmp2280;
	wire signed [31:0] w_sys_tmp2281;
	wire signed [31:0] w_sys_tmp2286;
	wire signed [31:0] w_sys_tmp2287;
	wire signed [31:0] w_sys_tmp2292;
	wire signed [31:0] w_sys_tmp2293;
	wire signed [31:0] w_sys_tmp2298;
	wire signed [31:0] w_sys_tmp2299;
	wire signed [31:0] w_sys_tmp2304;
	wire signed [31:0] w_sys_tmp2305;
	wire signed [31:0] w_sys_tmp2310;
	wire signed [31:0] w_sys_tmp2311;
	wire signed [31:0] w_sys_tmp2316;
	wire signed [31:0] w_sys_tmp2317;
	wire signed [31:0] w_sys_tmp2322;
	wire signed [31:0] w_sys_tmp2323;
	wire signed [31:0] w_sys_tmp2328;
	wire signed [31:0] w_sys_tmp2329;
	wire signed [31:0] w_sys_tmp2334;
	wire signed [31:0] w_sys_tmp2335;
	wire signed [31:0] w_sys_tmp2340;
	wire signed [31:0] w_sys_tmp2341;
	wire signed [31:0] w_sys_tmp2346;
	wire signed [31:0] w_sys_tmp2347;
	wire signed [31:0] w_sys_tmp2352;
	wire signed [31:0] w_sys_tmp2353;
	wire signed [31:0] w_sys_tmp2358;
	wire signed [31:0] w_sys_tmp2359;
	wire signed [31:0] w_sys_tmp2364;
	wire signed [31:0] w_sys_tmp2365;
	wire signed [31:0] w_sys_tmp2370;
	wire signed [31:0] w_sys_tmp2371;
	wire signed [31:0] w_sys_tmp2376;
	wire signed [31:0] w_sys_tmp2377;
	wire signed [31:0] w_sys_tmp2382;
	wire signed [31:0] w_sys_tmp2383;
	wire signed [31:0] w_sys_tmp2388;
	wire signed [31:0] w_sys_tmp2389;
	wire signed [31:0] w_sys_tmp2394;
	wire signed [31:0] w_sys_tmp2395;
	wire signed [31:0] w_sys_tmp2400;
	wire signed [31:0] w_sys_tmp2401;
	wire signed [31:0] w_sys_tmp2406;
	wire signed [31:0] w_sys_tmp2407;
	wire signed [31:0] w_sys_tmp2412;
	wire signed [31:0] w_sys_tmp2413;
	wire signed [31:0] w_sys_tmp2418;
	wire signed [31:0] w_sys_tmp2419;
	wire signed [31:0] w_sys_tmp2424;
	wire signed [31:0] w_sys_tmp2425;
	wire signed [31:0] w_sys_tmp2430;
	wire signed [31:0] w_sys_tmp2431;
	wire signed [31:0] w_sys_tmp2436;
	wire signed [31:0] w_sys_tmp2437;
	wire signed [31:0] w_sys_tmp2442;
	wire signed [31:0] w_sys_tmp2443;
	wire signed [31:0] w_sys_tmp2460;
	wire signed [31:0] w_sys_tmp2461;
	wire signed [31:0] w_sys_tmp2466;
	wire signed [31:0] w_sys_tmp2467;
	wire signed [31:0] w_sys_tmp2472;
	wire signed [31:0] w_sys_tmp2473;
	wire signed [31:0] w_sys_tmp2478;
	wire signed [31:0] w_sys_tmp2479;
	wire signed [31:0] w_sys_tmp2484;
	wire signed [31:0] w_sys_tmp2485;
	wire signed [31:0] w_sys_tmp2490;
	wire signed [31:0] w_sys_tmp2491;
	wire signed [31:0] w_sys_tmp2496;
	wire signed [31:0] w_sys_tmp2497;
	wire signed [31:0] w_sys_tmp2502;
	wire signed [31:0] w_sys_tmp2503;
	wire signed [31:0] w_sys_tmp2508;
	wire signed [31:0] w_sys_tmp2509;
	wire signed [31:0] w_sys_tmp2514;
	wire signed [31:0] w_sys_tmp2515;
	wire signed [31:0] w_sys_tmp2520;
	wire signed [31:0] w_sys_tmp2521;
	wire signed [31:0] w_sys_tmp2526;
	wire signed [31:0] w_sys_tmp2527;
	wire signed [31:0] w_sys_tmp2532;
	wire signed [31:0] w_sys_tmp2533;
	wire signed [31:0] w_sys_tmp2538;
	wire signed [31:0] w_sys_tmp2539;
	wire signed [31:0] w_sys_tmp2544;
	wire signed [31:0] w_sys_tmp2545;
	wire signed [31:0] w_sys_tmp2550;
	wire signed [31:0] w_sys_tmp2551;
	wire signed [31:0] w_sys_tmp2556;
	wire signed [31:0] w_sys_tmp2557;
	wire signed [31:0] w_sys_tmp2562;
	wire signed [31:0] w_sys_tmp2563;
	wire signed [31:0] w_sys_tmp2568;
	wire signed [31:0] w_sys_tmp2569;
	wire signed [31:0] w_sys_tmp2574;
	wire signed [31:0] w_sys_tmp2575;
	wire signed [31:0] w_sys_tmp2580;
	wire signed [31:0] w_sys_tmp2581;
	wire signed [31:0] w_sys_tmp2586;
	wire signed [31:0] w_sys_tmp2587;
	wire signed [31:0] w_sys_tmp2592;
	wire signed [31:0] w_sys_tmp2593;
	wire signed [31:0] w_sys_tmp2598;
	wire signed [31:0] w_sys_tmp2599;
	wire signed [31:0] w_sys_tmp2604;
	wire signed [31:0] w_sys_tmp2605;
	wire signed [31:0] w_sys_tmp2610;
	wire signed [31:0] w_sys_tmp2611;
	wire signed [31:0] w_sys_tmp2616;
	wire signed [31:0] w_sys_tmp2617;
	wire signed [31:0] w_sys_tmp2622;
	wire signed [31:0] w_sys_tmp2623;
	wire signed [31:0] w_sys_tmp2628;
	wire signed [31:0] w_sys_tmp2629;
	wire signed [31:0] w_sys_tmp2634;
	wire signed [31:0] w_sys_tmp2635;
	wire signed [31:0] w_sys_tmp2640;
	wire signed [31:0] w_sys_tmp2641;
	wire signed [31:0] w_sys_tmp2646;
	wire signed [31:0] w_sys_tmp2647;
	wire signed [31:0] w_sys_tmp2652;
	wire signed [31:0] w_sys_tmp2653;
	wire signed [31:0] w_sys_tmp2658;
	wire signed [31:0] w_sys_tmp2659;
	wire signed [31:0] w_sys_tmp2664;
	wire signed [31:0] w_sys_tmp2665;
	wire signed [31:0] w_sys_tmp2670;
	wire signed [31:0] w_sys_tmp2671;
	wire signed [31:0] w_sys_tmp2676;
	wire signed [31:0] w_sys_tmp2677;
	wire signed [31:0] w_sys_tmp2682;
	wire signed [31:0] w_sys_tmp2683;
	wire signed [31:0] w_sys_tmp2688;
	wire signed [31:0] w_sys_tmp2689;
	wire signed [31:0] w_sys_tmp2694;
	wire signed [31:0] w_sys_tmp2695;
	wire signed [31:0] w_sys_tmp2700;
	wire signed [31:0] w_sys_tmp2701;
	wire signed [31:0] w_sys_tmp2706;
	wire signed [31:0] w_sys_tmp2707;
	wire signed [31:0] w_sys_tmp2712;
	wire signed [31:0] w_sys_tmp2713;
	wire signed [31:0] w_sys_tmp2718;
	wire signed [31:0] w_sys_tmp2719;
	wire signed [31:0] w_sys_tmp2724;
	wire signed [31:0] w_sys_tmp2725;
	wire signed [31:0] w_sys_tmp2730;
	wire signed [31:0] w_sys_tmp2731;
	wire signed [31:0] w_sys_tmp2736;
	wire signed [31:0] w_sys_tmp2737;
	wire signed [31:0] w_sys_tmp2742;
	wire signed [31:0] w_sys_tmp2743;
	wire signed [31:0] w_sys_tmp2748;
	wire signed [31:0] w_sys_tmp2749;
	wire signed [31:0] w_sys_tmp2754;
	wire signed [31:0] w_sys_tmp2755;
	wire signed [31:0] w_sys_tmp2760;
	wire signed [31:0] w_sys_tmp2761;
	wire signed [31:0] w_sys_tmp2766;
	wire signed [31:0] w_sys_tmp2767;
	wire signed [31:0] w_sys_tmp2772;
	wire signed [31:0] w_sys_tmp2773;
	wire signed [31:0] w_sys_tmp2778;
	wire signed [31:0] w_sys_tmp2779;
	wire signed [31:0] w_sys_tmp2784;
	wire signed [31:0] w_sys_tmp2785;
	wire signed [31:0] w_sys_tmp2790;
	wire signed [31:0] w_sys_tmp2791;
	wire signed [31:0] w_sys_tmp2796;
	wire signed [31:0] w_sys_tmp2797;
	wire signed [31:0] w_sys_tmp2802;
	wire signed [31:0] w_sys_tmp2803;
	wire signed [31:0] w_sys_tmp2808;
	wire signed [31:0] w_sys_tmp2809;
	wire signed [31:0] w_sys_tmp2814;
	wire signed [31:0] w_sys_tmp2815;
	wire signed [31:0] w_sys_tmp2820;
	wire signed [31:0] w_sys_tmp2821;
	wire signed [31:0] w_sys_tmp2826;
	wire signed [31:0] w_sys_tmp2827;
	wire signed [31:0] w_sys_tmp2832;
	wire signed [31:0] w_sys_tmp2833;
	wire signed [31:0] w_sys_tmp2838;
	wire signed [31:0] w_sys_tmp2839;
	wire signed [31:0] w_sys_tmp2844;
	wire signed [31:0] w_sys_tmp2845;
	wire signed [31:0] w_sys_tmp2862;
	wire signed [31:0] w_sys_tmp2863;
	wire signed [31:0] w_sys_tmp2868;
	wire signed [31:0] w_sys_tmp2869;
	wire signed [31:0] w_sys_tmp2874;
	wire signed [31:0] w_sys_tmp2875;
	wire signed [31:0] w_sys_tmp2880;
	wire signed [31:0] w_sys_tmp2881;
	wire signed [31:0] w_sys_tmp2886;
	wire signed [31:0] w_sys_tmp2887;
	wire signed [31:0] w_sys_tmp2892;
	wire signed [31:0] w_sys_tmp2893;
	wire signed [31:0] w_sys_tmp2898;
	wire signed [31:0] w_sys_tmp2899;
	wire signed [31:0] w_sys_tmp2904;
	wire signed [31:0] w_sys_tmp2905;
	wire signed [31:0] w_sys_tmp2910;
	wire signed [31:0] w_sys_tmp2911;
	wire signed [31:0] w_sys_tmp2916;
	wire signed [31:0] w_sys_tmp2917;
	wire signed [31:0] w_sys_tmp2922;
	wire signed [31:0] w_sys_tmp2923;
	wire signed [31:0] w_sys_tmp2928;
	wire signed [31:0] w_sys_tmp2929;
	wire signed [31:0] w_sys_tmp2934;
	wire signed [31:0] w_sys_tmp2935;
	wire signed [31:0] w_sys_tmp2940;
	wire signed [31:0] w_sys_tmp2941;
	wire signed [31:0] w_sys_tmp2946;
	wire signed [31:0] w_sys_tmp2947;
	wire signed [31:0] w_sys_tmp2952;
	wire signed [31:0] w_sys_tmp2953;
	wire signed [31:0] w_sys_tmp2958;
	wire signed [31:0] w_sys_tmp2959;
	wire signed [31:0] w_sys_tmp2964;
	wire signed [31:0] w_sys_tmp2965;
	wire signed [31:0] w_sys_tmp2970;
	wire signed [31:0] w_sys_tmp2971;
	wire signed [31:0] w_sys_tmp2976;
	wire signed [31:0] w_sys_tmp2977;
	wire signed [31:0] w_sys_tmp2982;
	wire signed [31:0] w_sys_tmp2983;
	wire signed [31:0] w_sys_tmp2988;
	wire signed [31:0] w_sys_tmp2989;
	wire signed [31:0] w_sys_tmp2994;
	wire signed [31:0] w_sys_tmp2995;
	wire signed [31:0] w_sys_tmp3000;
	wire signed [31:0] w_sys_tmp3001;
	wire signed [31:0] w_sys_tmp3006;
	wire signed [31:0] w_sys_tmp3007;
	wire signed [31:0] w_sys_tmp3012;
	wire signed [31:0] w_sys_tmp3013;
	wire signed [31:0] w_sys_tmp3018;
	wire signed [31:0] w_sys_tmp3019;
	wire signed [31:0] w_sys_tmp3024;
	wire signed [31:0] w_sys_tmp3025;
	wire signed [31:0] w_sys_tmp3030;
	wire signed [31:0] w_sys_tmp3031;
	wire signed [31:0] w_sys_tmp3036;
	wire signed [31:0] w_sys_tmp3037;
	wire signed [31:0] w_sys_tmp3042;
	wire signed [31:0] w_sys_tmp3043;
	wire signed [31:0] w_sys_tmp3048;
	wire signed [31:0] w_sys_tmp3049;
	wire signed [31:0] w_sys_tmp3066;
	wire signed [31:0] w_sys_tmp3067;
	wire signed [31:0] w_sys_tmp3072;
	wire signed [31:0] w_sys_tmp3073;
	wire signed [31:0] w_sys_tmp3078;
	wire signed [31:0] w_sys_tmp3079;
	wire signed [31:0] w_sys_tmp3084;
	wire signed [31:0] w_sys_tmp3085;
	wire signed [31:0] w_sys_tmp3090;
	wire signed [31:0] w_sys_tmp3091;
	wire signed [31:0] w_sys_tmp3096;
	wire signed [31:0] w_sys_tmp3097;
	wire signed [31:0] w_sys_tmp3102;
	wire signed [31:0] w_sys_tmp3103;
	wire signed [31:0] w_sys_tmp3108;
	wire signed [31:0] w_sys_tmp3109;
	wire signed [31:0] w_sys_tmp3114;
	wire signed [31:0] w_sys_tmp3115;
	wire signed [31:0] w_sys_tmp3120;
	wire signed [31:0] w_sys_tmp3121;
	wire signed [31:0] w_sys_tmp3126;
	wire signed [31:0] w_sys_tmp3127;
	wire signed [31:0] w_sys_tmp3132;
	wire signed [31:0] w_sys_tmp3133;
	wire signed [31:0] w_sys_tmp3138;
	wire signed [31:0] w_sys_tmp3139;
	wire signed [31:0] w_sys_tmp3144;
	wire signed [31:0] w_sys_tmp3145;
	wire signed [31:0] w_sys_tmp3150;
	wire signed [31:0] w_sys_tmp3151;
	wire signed [31:0] w_sys_tmp3156;
	wire signed [31:0] w_sys_tmp3157;
	wire signed [31:0] w_sys_tmp3162;
	wire signed [31:0] w_sys_tmp3163;
	wire signed [31:0] w_sys_tmp3168;
	wire signed [31:0] w_sys_tmp3169;
	wire signed [31:0] w_sys_tmp3174;
	wire signed [31:0] w_sys_tmp3175;
	wire signed [31:0] w_sys_tmp3180;
	wire signed [31:0] w_sys_tmp3181;
	wire signed [31:0] w_sys_tmp3186;
	wire signed [31:0] w_sys_tmp3187;
	wire signed [31:0] w_sys_tmp3192;
	wire signed [31:0] w_sys_tmp3193;
	wire signed [31:0] w_sys_tmp3198;
	wire signed [31:0] w_sys_tmp3199;
	wire signed [31:0] w_sys_tmp3204;
	wire signed [31:0] w_sys_tmp3205;
	wire signed [31:0] w_sys_tmp3210;
	wire signed [31:0] w_sys_tmp3211;
	wire signed [31:0] w_sys_tmp3216;
	wire signed [31:0] w_sys_tmp3217;
	wire signed [31:0] w_sys_tmp3222;
	wire signed [31:0] w_sys_tmp3223;
	wire signed [31:0] w_sys_tmp3228;
	wire signed [31:0] w_sys_tmp3229;
	wire signed [31:0] w_sys_tmp3234;
	wire signed [31:0] w_sys_tmp3235;
	wire signed [31:0] w_sys_tmp3240;
	wire signed [31:0] w_sys_tmp3241;
	wire signed [31:0] w_sys_tmp3246;
	wire signed [31:0] w_sys_tmp3247;
	wire signed [31:0] w_sys_tmp3252;
	wire signed [31:0] w_sys_tmp3253;
	wire signed [31:0] w_sys_tmp3270;
	wire signed [31:0] w_sys_tmp3271;
	wire signed [31:0] w_sys_tmp3276;
	wire signed [31:0] w_sys_tmp3277;
	wire signed [31:0] w_sys_tmp3282;
	wire signed [31:0] w_sys_tmp3283;
	wire signed [31:0] w_sys_tmp3288;
	wire signed [31:0] w_sys_tmp3289;
	wire signed [31:0] w_sys_tmp3294;
	wire signed [31:0] w_sys_tmp3295;
	wire signed [31:0] w_sys_tmp3300;
	wire signed [31:0] w_sys_tmp3301;
	wire signed [31:0] w_sys_tmp3306;
	wire signed [31:0] w_sys_tmp3307;
	wire signed [31:0] w_sys_tmp3312;
	wire signed [31:0] w_sys_tmp3313;
	wire signed [31:0] w_sys_tmp3318;
	wire signed [31:0] w_sys_tmp3319;
	wire signed [31:0] w_sys_tmp3324;
	wire signed [31:0] w_sys_tmp3325;
	wire signed [31:0] w_sys_tmp3330;
	wire signed [31:0] w_sys_tmp3331;
	wire signed [31:0] w_sys_tmp3336;
	wire signed [31:0] w_sys_tmp3337;
	wire signed [31:0] w_sys_tmp3342;
	wire signed [31:0] w_sys_tmp3343;
	wire signed [31:0] w_sys_tmp3348;
	wire signed [31:0] w_sys_tmp3349;
	wire signed [31:0] w_sys_tmp3354;
	wire signed [31:0] w_sys_tmp3355;
	wire signed [31:0] w_sys_tmp3360;
	wire signed [31:0] w_sys_tmp3361;
	wire signed [31:0] w_sys_tmp3366;
	wire signed [31:0] w_sys_tmp3367;
	wire signed [31:0] w_sys_tmp3372;
	wire signed [31:0] w_sys_tmp3373;
	wire signed [31:0] w_sys_tmp3378;
	wire signed [31:0] w_sys_tmp3379;
	wire signed [31:0] w_sys_tmp3384;
	wire signed [31:0] w_sys_tmp3385;
	wire signed [31:0] w_sys_tmp3390;
	wire signed [31:0] w_sys_tmp3391;
	wire signed [31:0] w_sys_tmp3396;
	wire signed [31:0] w_sys_tmp3397;
	wire signed [31:0] w_sys_tmp3402;
	wire signed [31:0] w_sys_tmp3403;
	wire signed [31:0] w_sys_tmp3408;
	wire signed [31:0] w_sys_tmp3409;
	wire signed [31:0] w_sys_tmp3414;
	wire signed [31:0] w_sys_tmp3415;
	wire signed [31:0] w_sys_tmp3420;
	wire signed [31:0] w_sys_tmp3421;
	wire signed [31:0] w_sys_tmp3426;
	wire signed [31:0] w_sys_tmp3427;
	wire signed [31:0] w_sys_tmp3432;
	wire signed [31:0] w_sys_tmp3433;
	wire signed [31:0] w_sys_tmp3438;
	wire signed [31:0] w_sys_tmp3439;
	wire signed [31:0] w_sys_tmp3444;
	wire signed [31:0] w_sys_tmp3445;
	wire signed [31:0] w_sys_tmp3450;
	wire signed [31:0] w_sys_tmp3451;
	wire signed [31:0] w_sys_tmp3456;
	wire signed [31:0] w_sys_tmp3457;
	wire signed [31:0] w_sys_tmp3461;
	wire signed [31:0] w_sys_tmp3462;
	wire               w_sys_tmp3463;
	wire               w_sys_tmp3464;
	wire signed [31:0] w_sys_tmp3465;
	wire signed [31:0] w_sys_tmp3468;
	wire signed [31:0] w_sys_tmp3469;
	wire        [31:0] w_sys_tmp3470;
	wire signed [31:0] w_sys_tmp3474;
	wire signed [31:0] w_sys_tmp3475;
	wire signed [31:0] w_sys_tmp3480;
	wire signed [31:0] w_sys_tmp3481;
	wire signed [31:0] w_sys_tmp3486;
	wire signed [31:0] w_sys_tmp3487;
	wire signed [31:0] w_sys_tmp3492;
	wire signed [31:0] w_sys_tmp3493;
	wire signed [31:0] w_sys_tmp3498;
	wire signed [31:0] w_sys_tmp3499;
	wire signed [31:0] w_sys_tmp3504;
	wire signed [31:0] w_sys_tmp3505;
	wire signed [31:0] w_sys_tmp3510;
	wire signed [31:0] w_sys_tmp3511;
	wire signed [31:0] w_sys_tmp3516;
	wire signed [31:0] w_sys_tmp3517;
	wire signed [31:0] w_sys_tmp3522;
	wire signed [31:0] w_sys_tmp3523;
	wire signed [31:0] w_sys_tmp3528;
	wire signed [31:0] w_sys_tmp3529;
	wire signed [31:0] w_sys_tmp3534;
	wire signed [31:0] w_sys_tmp3535;
	wire signed [31:0] w_sys_tmp3540;
	wire signed [31:0] w_sys_tmp3541;
	wire signed [31:0] w_sys_tmp3546;
	wire signed [31:0] w_sys_tmp3547;
	wire signed [31:0] w_sys_tmp3552;
	wire signed [31:0] w_sys_tmp3553;
	wire signed [31:0] w_sys_tmp3558;
	wire signed [31:0] w_sys_tmp3559;
	wire signed [31:0] w_sys_tmp3564;
	wire signed [31:0] w_sys_tmp3565;
	wire signed [31:0] w_sys_tmp3570;
	wire signed [31:0] w_sys_tmp3571;
	wire signed [31:0] w_sys_tmp3576;
	wire signed [31:0] w_sys_tmp3577;
	wire signed [31:0] w_sys_tmp3582;
	wire signed [31:0] w_sys_tmp3583;
	wire signed [31:0] w_sys_tmp3588;
	wire signed [31:0] w_sys_tmp3589;
	wire signed [31:0] w_sys_tmp3594;
	wire signed [31:0] w_sys_tmp3595;
	wire signed [31:0] w_sys_tmp3600;
	wire signed [31:0] w_sys_tmp3601;
	wire signed [31:0] w_sys_tmp3606;
	wire signed [31:0] w_sys_tmp3607;
	wire signed [31:0] w_sys_tmp3612;
	wire signed [31:0] w_sys_tmp3613;
	wire signed [31:0] w_sys_tmp3618;
	wire signed [31:0] w_sys_tmp3619;
	wire signed [31:0] w_sys_tmp3624;
	wire signed [31:0] w_sys_tmp3625;
	wire signed [31:0] w_sys_tmp3630;
	wire signed [31:0] w_sys_tmp3631;
	wire signed [31:0] w_sys_tmp3636;
	wire signed [31:0] w_sys_tmp3637;
	wire signed [31:0] w_sys_tmp3642;
	wire signed [31:0] w_sys_tmp3643;
	wire signed [31:0] w_sys_tmp3648;
	wire signed [31:0] w_sys_tmp3649;
	wire signed [31:0] w_sys_tmp3654;
	wire signed [31:0] w_sys_tmp3655;
	wire signed [31:0] w_sys_tmp3659;
	wire signed [31:0] w_sys_tmp3660;
	wire signed [31:0] w_sys_tmp3664;
	wire signed [31:0] w_sys_tmp3665;
	wire signed [31:0] w_sys_tmp3669;
	wire signed [31:0] w_sys_tmp3670;
	wire signed [31:0] w_sys_tmp3674;
	wire signed [31:0] w_sys_tmp3675;
	wire signed [31:0] w_sys_tmp3679;
	wire signed [31:0] w_sys_tmp3680;
	wire signed [31:0] w_sys_tmp3684;
	wire signed [31:0] w_sys_tmp3685;
	wire signed [31:0] w_sys_tmp3689;
	wire signed [31:0] w_sys_tmp3690;
	wire signed [31:0] w_sys_tmp3694;
	wire signed [31:0] w_sys_tmp3695;
	wire signed [31:0] w_sys_tmp3699;
	wire signed [31:0] w_sys_tmp3700;
	wire signed [31:0] w_sys_tmp3704;
	wire signed [31:0] w_sys_tmp3705;
	wire signed [31:0] w_sys_tmp3709;
	wire signed [31:0] w_sys_tmp3710;
	wire signed [31:0] w_sys_tmp3714;
	wire signed [31:0] w_sys_tmp3715;
	wire signed [31:0] w_sys_tmp3719;
	wire signed [31:0] w_sys_tmp3720;
	wire signed [31:0] w_sys_tmp3724;
	wire signed [31:0] w_sys_tmp3725;
	wire signed [31:0] w_sys_tmp3729;
	wire signed [31:0] w_sys_tmp3730;
	wire signed [31:0] w_sys_tmp3734;
	wire signed [31:0] w_sys_tmp3735;
	wire signed [31:0] w_sys_tmp3739;
	wire signed [31:0] w_sys_tmp3740;
	wire signed [31:0] w_sys_tmp3744;
	wire signed [31:0] w_sys_tmp3745;
	wire signed [31:0] w_sys_tmp3749;
	wire signed [31:0] w_sys_tmp3750;
	wire signed [31:0] w_sys_tmp3754;
	wire signed [31:0] w_sys_tmp3755;
	wire signed [31:0] w_sys_tmp3759;
	wire signed [31:0] w_sys_tmp3760;
	wire signed [31:0] w_sys_tmp3764;
	wire signed [31:0] w_sys_tmp3765;
	wire signed [31:0] w_sys_tmp3769;
	wire signed [31:0] w_sys_tmp3770;
	wire signed [31:0] w_sys_tmp3774;
	wire signed [31:0] w_sys_tmp3775;
	wire signed [31:0] w_sys_tmp3779;
	wire signed [31:0] w_sys_tmp3780;
	wire signed [31:0] w_sys_tmp3784;
	wire signed [31:0] w_sys_tmp3785;
	wire signed [31:0] w_sys_tmp3789;
	wire signed [31:0] w_sys_tmp3790;
	wire signed [31:0] w_sys_tmp3794;
	wire signed [31:0] w_sys_tmp3795;
	wire signed [31:0] w_sys_tmp3799;
	wire signed [31:0] w_sys_tmp3800;
	wire signed [31:0] w_sys_tmp3804;
	wire signed [31:0] w_sys_tmp3805;
	wire signed [31:0] w_sys_tmp3809;
	wire signed [31:0] w_sys_tmp3810;
	wire signed [31:0] w_sys_tmp3814;
	wire signed [31:0] w_sys_tmp3815;
	wire signed [31:0] w_sys_tmp3819;
	wire signed [31:0] w_sys_tmp3820;
	wire signed [31:0] w_sys_tmp3824;
	wire signed [31:0] w_sys_tmp3825;
	wire signed [31:0] w_sys_tmp3829;
	wire signed [31:0] w_sys_tmp3830;
	wire signed [31:0] w_sys_tmp3834;
	wire signed [31:0] w_sys_tmp3835;
	wire signed [31:0] w_sys_tmp3839;
	wire signed [31:0] w_sys_tmp3840;
	wire signed [31:0] w_sys_tmp3844;
	wire signed [31:0] w_sys_tmp3845;
	wire signed [31:0] w_sys_tmp3849;
	wire signed [31:0] w_sys_tmp3850;
	wire signed [31:0] w_sys_tmp3854;
	wire signed [31:0] w_sys_tmp3855;
	wire signed [31:0] w_sys_tmp3859;
	wire signed [31:0] w_sys_tmp3860;
	wire signed [31:0] w_sys_tmp3864;
	wire signed [31:0] w_sys_tmp3865;
	wire signed [31:0] w_sys_tmp3869;
	wire signed [31:0] w_sys_tmp3870;
	wire signed [31:0] w_sys_tmp3874;
	wire signed [31:0] w_sys_tmp3875;
	wire signed [31:0] w_sys_tmp3879;
	wire signed [31:0] w_sys_tmp3880;
	wire signed [31:0] w_sys_tmp3884;
	wire signed [31:0] w_sys_tmp3885;
	wire signed [31:0] w_sys_tmp3889;
	wire signed [31:0] w_sys_tmp3890;
	wire signed [31:0] w_sys_tmp3894;
	wire signed [31:0] w_sys_tmp3895;
	wire signed [31:0] w_sys_tmp3899;
	wire signed [31:0] w_sys_tmp3900;
	wire signed [31:0] w_sys_tmp3904;
	wire signed [31:0] w_sys_tmp3905;
	wire signed [31:0] w_sys_tmp3909;
	wire signed [31:0] w_sys_tmp3910;
	wire signed [31:0] w_sys_tmp3914;
	wire signed [31:0] w_sys_tmp3915;
	wire signed [31:0] w_sys_tmp3919;
	wire signed [31:0] w_sys_tmp3920;
	wire signed [31:0] w_sys_tmp3924;
	wire signed [31:0] w_sys_tmp3925;
	wire signed [31:0] w_sys_tmp3929;
	wire signed [31:0] w_sys_tmp3930;
	wire signed [31:0] w_sys_tmp3934;
	wire signed [31:0] w_sys_tmp3935;
	wire signed [31:0] w_sys_tmp3939;
	wire signed [31:0] w_sys_tmp3940;
	wire signed [31:0] w_sys_tmp3944;
	wire signed [31:0] w_sys_tmp3945;
	wire signed [31:0] w_sys_tmp3949;
	wire signed [31:0] w_sys_tmp3950;
	wire signed [31:0] w_sys_tmp3954;
	wire signed [31:0] w_sys_tmp3955;
	wire signed [31:0] w_sys_tmp3959;
	wire signed [31:0] w_sys_tmp3960;
	wire signed [31:0] w_sys_tmp3964;
	wire signed [31:0] w_sys_tmp3965;
	wire signed [31:0] w_sys_tmp3969;
	wire signed [31:0] w_sys_tmp3970;
	wire signed [31:0] w_sys_tmp3974;
	wire signed [31:0] w_sys_tmp3975;
	wire signed [31:0] w_sys_tmp3979;
	wire signed [31:0] w_sys_tmp3980;
	wire signed [31:0] w_sys_tmp3984;
	wire signed [31:0] w_sys_tmp3985;
	wire signed [31:0] w_sys_tmp3989;
	wire signed [31:0] w_sys_tmp3990;
	wire signed [31:0] w_sys_tmp3994;
	wire signed [31:0] w_sys_tmp3995;
	wire signed [31:0] w_sys_tmp3999;
	wire signed [31:0] w_sys_tmp4000;
	wire signed [31:0] w_sys_tmp4004;
	wire signed [31:0] w_sys_tmp4005;
	wire signed [31:0] w_sys_tmp4009;
	wire signed [31:0] w_sys_tmp4010;
	wire signed [31:0] w_sys_tmp4014;
	wire signed [31:0] w_sys_tmp4015;
	wire signed [31:0] w_sys_tmp4019;
	wire signed [31:0] w_sys_tmp4020;
	wire signed [31:0] w_sys_tmp4024;
	wire signed [31:0] w_sys_tmp4025;
	wire signed [31:0] w_sys_tmp4029;
	wire signed [31:0] w_sys_tmp4030;
	wire signed [31:0] w_sys_tmp4034;
	wire signed [31:0] w_sys_tmp4035;
	wire signed [31:0] w_sys_tmp4039;
	wire signed [31:0] w_sys_tmp4040;
	wire signed [31:0] w_sys_tmp4044;
	wire signed [31:0] w_sys_tmp4045;
	wire signed [31:0] w_sys_tmp4049;
	wire signed [31:0] w_sys_tmp4050;
	wire signed [31:0] w_sys_tmp4054;
	wire signed [31:0] w_sys_tmp4055;
	wire signed [31:0] w_sys_tmp4059;
	wire signed [31:0] w_sys_tmp4060;
	wire signed [31:0] w_sys_tmp4064;
	wire signed [31:0] w_sys_tmp4065;
	wire signed [31:0] w_sys_tmp4069;
	wire signed [31:0] w_sys_tmp4070;
	wire signed [31:0] w_sys_tmp4074;
	wire signed [31:0] w_sys_tmp4075;
	wire signed [31:0] w_sys_tmp4079;
	wire signed [31:0] w_sys_tmp4080;
	wire signed [31:0] w_sys_tmp4084;
	wire signed [31:0] w_sys_tmp4085;
	wire signed [31:0] w_sys_tmp4089;
	wire signed [31:0] w_sys_tmp4090;
	wire signed [31:0] w_sys_tmp4094;
	wire signed [31:0] w_sys_tmp4095;
	wire signed [31:0] w_sys_tmp4099;
	wire signed [31:0] w_sys_tmp4100;
	wire signed [31:0] w_sys_tmp4104;
	wire signed [31:0] w_sys_tmp4105;
	wire signed [31:0] w_sys_tmp4109;
	wire signed [31:0] w_sys_tmp4110;
	wire signed [31:0] w_sys_tmp4114;
	wire signed [31:0] w_sys_tmp4115;
	wire signed [31:0] w_sys_tmp4119;
	wire signed [31:0] w_sys_tmp4120;
	wire signed [31:0] w_sys_tmp4124;
	wire signed [31:0] w_sys_tmp4125;
	wire signed [31:0] w_sys_tmp4129;
	wire signed [31:0] w_sys_tmp4130;
	wire signed [31:0] w_sys_tmp4133;
	wire signed [31:0] w_sys_tmp4134;
	wire               w_sys_tmp4135;
	wire               w_sys_tmp4136;
	wire signed [31:0] w_sys_tmp4137;
	wire signed [31:0] w_sys_tmp4140;
	wire signed [31:0] w_sys_tmp4141;
	wire        [31:0] w_sys_tmp4142;
	wire signed [31:0] w_sys_tmp4146;
	wire signed [31:0] w_sys_tmp4147;
	wire signed [31:0] w_sys_tmp4152;
	wire signed [31:0] w_sys_tmp4153;
	wire signed [31:0] w_sys_tmp4158;
	wire signed [31:0] w_sys_tmp4159;
	wire signed [31:0] w_sys_tmp4164;
	wire signed [31:0] w_sys_tmp4165;
	wire signed [31:0] w_sys_tmp4170;
	wire signed [31:0] w_sys_tmp4171;
	wire signed [31:0] w_sys_tmp4176;
	wire signed [31:0] w_sys_tmp4177;
	wire signed [31:0] w_sys_tmp4182;
	wire signed [31:0] w_sys_tmp4183;
	wire signed [31:0] w_sys_tmp4188;
	wire signed [31:0] w_sys_tmp4189;
	wire signed [31:0] w_sys_tmp4194;
	wire signed [31:0] w_sys_tmp4195;
	wire signed [31:0] w_sys_tmp4200;
	wire signed [31:0] w_sys_tmp4201;
	wire signed [31:0] w_sys_tmp4206;
	wire signed [31:0] w_sys_tmp4207;
	wire signed [31:0] w_sys_tmp4212;
	wire signed [31:0] w_sys_tmp4213;
	wire signed [31:0] w_sys_tmp4218;
	wire signed [31:0] w_sys_tmp4219;
	wire signed [31:0] w_sys_tmp4224;
	wire signed [31:0] w_sys_tmp4225;
	wire signed [31:0] w_sys_tmp4230;
	wire signed [31:0] w_sys_tmp4231;
	wire signed [31:0] w_sys_tmp4236;
	wire signed [31:0] w_sys_tmp4237;
	wire signed [31:0] w_sys_tmp4242;
	wire signed [31:0] w_sys_tmp4243;
	wire signed [31:0] w_sys_tmp4248;
	wire signed [31:0] w_sys_tmp4249;
	wire signed [31:0] w_sys_tmp4254;
	wire signed [31:0] w_sys_tmp4255;
	wire signed [31:0] w_sys_tmp4260;
	wire signed [31:0] w_sys_tmp4261;
	wire signed [31:0] w_sys_tmp4266;
	wire signed [31:0] w_sys_tmp4267;
	wire signed [31:0] w_sys_tmp4272;
	wire signed [31:0] w_sys_tmp4273;
	wire signed [31:0] w_sys_tmp4278;
	wire signed [31:0] w_sys_tmp4279;
	wire signed [31:0] w_sys_tmp4284;
	wire signed [31:0] w_sys_tmp4285;
	wire signed [31:0] w_sys_tmp4290;
	wire signed [31:0] w_sys_tmp4291;
	wire signed [31:0] w_sys_tmp4296;
	wire signed [31:0] w_sys_tmp4297;
	wire signed [31:0] w_sys_tmp4302;
	wire signed [31:0] w_sys_tmp4303;
	wire signed [31:0] w_sys_tmp4308;
	wire signed [31:0] w_sys_tmp4309;
	wire signed [31:0] w_sys_tmp4314;
	wire signed [31:0] w_sys_tmp4315;
	wire signed [31:0] w_sys_tmp4320;
	wire signed [31:0] w_sys_tmp4321;
	wire signed [31:0] w_sys_tmp4326;
	wire signed [31:0] w_sys_tmp4327;
	wire signed [31:0] w_sys_tmp4331;
	wire signed [31:0] w_sys_tmp4332;
	wire signed [31:0] w_sys_tmp4336;
	wire signed [31:0] w_sys_tmp4337;
	wire signed [31:0] w_sys_tmp4341;
	wire signed [31:0] w_sys_tmp4342;
	wire signed [31:0] w_sys_tmp4346;
	wire signed [31:0] w_sys_tmp4347;
	wire signed [31:0] w_sys_tmp4351;
	wire signed [31:0] w_sys_tmp4352;
	wire signed [31:0] w_sys_tmp4356;
	wire signed [31:0] w_sys_tmp4357;
	wire signed [31:0] w_sys_tmp4361;
	wire signed [31:0] w_sys_tmp4362;
	wire signed [31:0] w_sys_tmp4366;
	wire signed [31:0] w_sys_tmp4367;
	wire signed [31:0] w_sys_tmp4371;
	wire signed [31:0] w_sys_tmp4372;
	wire signed [31:0] w_sys_tmp4376;
	wire signed [31:0] w_sys_tmp4377;
	wire signed [31:0] w_sys_tmp4381;
	wire signed [31:0] w_sys_tmp4382;
	wire signed [31:0] w_sys_tmp4386;
	wire signed [31:0] w_sys_tmp4387;
	wire signed [31:0] w_sys_tmp4391;
	wire signed [31:0] w_sys_tmp4392;
	wire signed [31:0] w_sys_tmp4396;
	wire signed [31:0] w_sys_tmp4397;
	wire signed [31:0] w_sys_tmp4401;
	wire signed [31:0] w_sys_tmp4402;
	wire signed [31:0] w_sys_tmp4406;
	wire signed [31:0] w_sys_tmp4407;
	wire signed [31:0] w_sys_tmp4411;
	wire signed [31:0] w_sys_tmp4412;
	wire signed [31:0] w_sys_tmp4416;
	wire signed [31:0] w_sys_tmp4417;
	wire signed [31:0] w_sys_tmp4421;
	wire signed [31:0] w_sys_tmp4422;
	wire signed [31:0] w_sys_tmp4426;
	wire signed [31:0] w_sys_tmp4427;
	wire signed [31:0] w_sys_tmp4431;
	wire signed [31:0] w_sys_tmp4432;
	wire signed [31:0] w_sys_tmp4436;
	wire signed [31:0] w_sys_tmp4437;
	wire signed [31:0] w_sys_tmp4441;
	wire signed [31:0] w_sys_tmp4442;
	wire signed [31:0] w_sys_tmp4446;
	wire signed [31:0] w_sys_tmp4447;
	wire signed [31:0] w_sys_tmp4451;
	wire signed [31:0] w_sys_tmp4452;
	wire signed [31:0] w_sys_tmp4456;
	wire signed [31:0] w_sys_tmp4457;
	wire signed [31:0] w_sys_tmp4461;
	wire signed [31:0] w_sys_tmp4462;
	wire signed [31:0] w_sys_tmp4466;
	wire signed [31:0] w_sys_tmp4467;
	wire signed [31:0] w_sys_tmp4471;
	wire signed [31:0] w_sys_tmp4472;
	wire signed [31:0] w_sys_tmp4476;
	wire signed [31:0] w_sys_tmp4477;
	wire signed [31:0] w_sys_tmp4481;
	wire signed [31:0] w_sys_tmp4482;
	wire signed [31:0] w_sys_tmp4486;
	wire signed [31:0] w_sys_tmp4487;
	wire signed [31:0] w_sys_tmp4491;
	wire signed [31:0] w_sys_tmp4492;
	wire signed [31:0] w_sys_tmp4496;
	wire signed [31:0] w_sys_tmp4497;
	wire signed [31:0] w_sys_tmp4501;
	wire signed [31:0] w_sys_tmp4502;
	wire signed [31:0] w_sys_tmp4506;
	wire signed [31:0] w_sys_tmp4507;
	wire signed [31:0] w_sys_tmp4511;
	wire signed [31:0] w_sys_tmp4512;
	wire signed [31:0] w_sys_tmp4516;
	wire signed [31:0] w_sys_tmp4517;
	wire signed [31:0] w_sys_tmp4521;
	wire signed [31:0] w_sys_tmp4522;
	wire signed [31:0] w_sys_tmp4526;
	wire signed [31:0] w_sys_tmp4527;
	wire signed [31:0] w_sys_tmp4531;
	wire signed [31:0] w_sys_tmp4532;
	wire signed [31:0] w_sys_tmp4536;
	wire signed [31:0] w_sys_tmp4537;
	wire signed [31:0] w_sys_tmp4541;
	wire signed [31:0] w_sys_tmp4542;
	wire signed [31:0] w_sys_tmp4546;
	wire signed [31:0] w_sys_tmp4547;
	wire signed [31:0] w_sys_tmp4551;
	wire signed [31:0] w_sys_tmp4552;
	wire signed [31:0] w_sys_tmp4556;
	wire signed [31:0] w_sys_tmp4557;
	wire signed [31:0] w_sys_tmp4561;
	wire signed [31:0] w_sys_tmp4562;
	wire signed [31:0] w_sys_tmp4566;
	wire signed [31:0] w_sys_tmp4567;
	wire signed [31:0] w_sys_tmp4571;
	wire signed [31:0] w_sys_tmp4572;
	wire signed [31:0] w_sys_tmp4576;
	wire signed [31:0] w_sys_tmp4577;
	wire signed [31:0] w_sys_tmp4581;
	wire signed [31:0] w_sys_tmp4582;
	wire signed [31:0] w_sys_tmp4586;
	wire signed [31:0] w_sys_tmp4587;
	wire signed [31:0] w_sys_tmp4591;
	wire signed [31:0] w_sys_tmp4592;
	wire signed [31:0] w_sys_tmp4596;
	wire signed [31:0] w_sys_tmp4597;
	wire signed [31:0] w_sys_tmp4601;
	wire signed [31:0] w_sys_tmp4602;
	wire signed [31:0] w_sys_tmp4606;
	wire signed [31:0] w_sys_tmp4607;
	wire signed [31:0] w_sys_tmp4611;
	wire signed [31:0] w_sys_tmp4612;
	wire signed [31:0] w_sys_tmp4616;
	wire signed [31:0] w_sys_tmp4617;
	wire signed [31:0] w_sys_tmp4621;
	wire signed [31:0] w_sys_tmp4622;
	wire signed [31:0] w_sys_tmp4626;
	wire signed [31:0] w_sys_tmp4627;
	wire signed [31:0] w_sys_tmp4631;
	wire signed [31:0] w_sys_tmp4632;
	wire signed [31:0] w_sys_tmp4636;
	wire signed [31:0] w_sys_tmp4637;
	wire signed [31:0] w_sys_tmp4641;
	wire signed [31:0] w_sys_tmp4642;
	wire signed [31:0] w_sys_tmp4646;
	wire signed [31:0] w_sys_tmp4647;
	wire signed [31:0] w_sys_tmp4651;
	wire signed [31:0] w_sys_tmp4652;
	wire signed [31:0] w_sys_tmp4656;
	wire signed [31:0] w_sys_tmp4657;
	wire signed [31:0] w_sys_tmp4661;
	wire signed [31:0] w_sys_tmp4662;
	wire signed [31:0] w_sys_tmp4666;
	wire signed [31:0] w_sys_tmp4667;
	wire signed [31:0] w_sys_tmp4671;
	wire signed [31:0] w_sys_tmp4672;
	wire signed [31:0] w_sys_tmp4676;
	wire signed [31:0] w_sys_tmp4677;
	wire signed [31:0] w_sys_tmp4681;
	wire signed [31:0] w_sys_tmp4682;
	wire signed [31:0] w_sys_tmp4686;
	wire signed [31:0] w_sys_tmp4687;
	wire signed [31:0] w_sys_tmp4691;
	wire signed [31:0] w_sys_tmp4692;
	wire signed [31:0] w_sys_tmp4696;
	wire signed [31:0] w_sys_tmp4697;
	wire signed [31:0] w_sys_tmp4701;
	wire signed [31:0] w_sys_tmp4702;
	wire signed [31:0] w_sys_tmp4706;
	wire signed [31:0] w_sys_tmp4707;
	wire signed [31:0] w_sys_tmp4711;
	wire signed [31:0] w_sys_tmp4712;
	wire signed [31:0] w_sys_tmp4716;
	wire signed [31:0] w_sys_tmp4717;
	wire signed [31:0] w_sys_tmp4721;
	wire signed [31:0] w_sys_tmp4722;
	wire signed [31:0] w_sys_tmp4726;
	wire signed [31:0] w_sys_tmp4727;
	wire signed [31:0] w_sys_tmp4731;
	wire signed [31:0] w_sys_tmp4732;
	wire signed [31:0] w_sys_tmp4736;
	wire signed [31:0] w_sys_tmp4737;
	wire signed [31:0] w_sys_tmp4741;
	wire signed [31:0] w_sys_tmp4742;
	wire signed [31:0] w_sys_tmp4746;
	wire signed [31:0] w_sys_tmp4747;
	wire signed [31:0] w_sys_tmp4751;
	wire signed [31:0] w_sys_tmp4752;
	wire signed [31:0] w_sys_tmp4756;
	wire signed [31:0] w_sys_tmp4757;
	wire signed [31:0] w_sys_tmp4761;
	wire signed [31:0] w_sys_tmp4762;
	wire signed [31:0] w_sys_tmp4766;
	wire signed [31:0] w_sys_tmp4767;
	wire signed [31:0] w_sys_tmp4771;
	wire signed [31:0] w_sys_tmp4772;
	wire signed [31:0] w_sys_tmp4776;
	wire signed [31:0] w_sys_tmp4777;
	wire signed [31:0] w_sys_tmp4781;
	wire signed [31:0] w_sys_tmp4782;
	wire signed [31:0] w_sys_tmp4786;
	wire signed [31:0] w_sys_tmp4787;
	wire signed [31:0] w_sys_tmp4791;
	wire signed [31:0] w_sys_tmp4792;
	wire signed [31:0] w_sys_tmp4796;
	wire signed [31:0] w_sys_tmp4797;
	wire signed [31:0] w_sys_tmp4801;
	wire signed [31:0] w_sys_tmp4802;
	wire signed [31:0] w_sys_tmp4806;
	wire signed [31:0] w_sys_tmp4807;
	wire signed [31:0] w_sys_tmp4811;
	wire signed [31:0] w_sys_tmp4812;
	wire signed [31:0] w_sys_tmp4816;
	wire signed [31:0] w_sys_tmp4817;
	wire signed [31:0] w_sys_tmp4821;
	wire signed [31:0] w_sys_tmp4822;
	wire signed [31:0] w_sys_tmp4826;
	wire signed [31:0] w_sys_tmp4827;
	wire signed [31:0] w_sys_tmp4831;
	wire signed [31:0] w_sys_tmp4832;
	wire signed [31:0] w_sys_tmp4836;
	wire signed [31:0] w_sys_tmp4837;
	wire signed [31:0] w_sys_tmp4841;
	wire signed [31:0] w_sys_tmp4842;
	wire signed [31:0] w_sys_tmp4846;
	wire signed [31:0] w_sys_tmp4847;
	wire signed [31:0] w_sys_tmp4851;
	wire signed [31:0] w_sys_tmp4852;
	wire signed [31:0] w_sys_tmp4856;
	wire signed [31:0] w_sys_tmp4857;
	wire signed [31:0] w_sys_tmp4861;
	wire signed [31:0] w_sys_tmp4862;
	wire signed [31:0] w_sys_tmp4866;
	wire signed [31:0] w_sys_tmp4867;
	wire signed [31:0] w_sys_tmp4871;
	wire signed [31:0] w_sys_tmp4872;
	wire signed [31:0] w_sys_tmp4876;
	wire signed [31:0] w_sys_tmp4877;
	wire signed [31:0] w_sys_tmp4881;
	wire signed [31:0] w_sys_tmp4882;
	wire signed [31:0] w_sys_tmp4886;
	wire signed [31:0] w_sys_tmp4887;
	wire signed [31:0] w_sys_tmp4891;
	wire signed [31:0] w_sys_tmp4892;
	wire signed [31:0] w_sys_tmp4896;
	wire signed [31:0] w_sys_tmp4897;
	wire signed [31:0] w_sys_tmp4901;
	wire signed [31:0] w_sys_tmp4902;
	wire signed [31:0] w_sys_tmp4906;
	wire signed [31:0] w_sys_tmp4907;
	wire signed [31:0] w_sys_tmp4911;
	wire signed [31:0] w_sys_tmp4912;
	wire signed [31:0] w_sys_tmp4916;
	wire signed [31:0] w_sys_tmp4917;
	wire signed [31:0] w_sys_tmp4921;
	wire signed [31:0] w_sys_tmp4922;
	wire signed [31:0] w_sys_tmp4926;
	wire signed [31:0] w_sys_tmp4927;
	wire signed [31:0] w_sys_tmp4931;
	wire signed [31:0] w_sys_tmp4932;
	wire signed [31:0] w_sys_tmp4936;
	wire signed [31:0] w_sys_tmp4937;
	wire signed [31:0] w_sys_tmp4941;
	wire signed [31:0] w_sys_tmp4942;
	wire signed [31:0] w_sys_tmp4946;
	wire signed [31:0] w_sys_tmp4947;
	wire signed [31:0] w_sys_tmp4951;
	wire signed [31:0] w_sys_tmp4952;
	wire signed [31:0] w_sys_tmp4956;
	wire signed [31:0] w_sys_tmp4957;
	wire signed [31:0] w_sys_tmp4961;
	wire signed [31:0] w_sys_tmp4962;
	wire signed [31:0] w_sys_tmp4966;
	wire signed [31:0] w_sys_tmp4967;
	wire signed [31:0] w_sys_tmp4971;
	wire signed [31:0] w_sys_tmp4972;
	wire signed [31:0] w_sys_tmp4976;
	wire signed [31:0] w_sys_tmp4977;
	wire signed [31:0] w_sys_tmp4981;
	wire signed [31:0] w_sys_tmp4982;
	wire signed [31:0] w_sys_tmp4986;
	wire signed [31:0] w_sys_tmp4987;
	wire signed [31:0] w_sys_tmp4991;
	wire signed [31:0] w_sys_tmp4992;
	wire signed [31:0] w_sys_tmp4996;
	wire signed [31:0] w_sys_tmp4997;
	wire signed [31:0] w_sys_tmp5001;
	wire signed [31:0] w_sys_tmp5002;
	wire signed [31:0] w_sys_tmp5006;
	wire signed [31:0] w_sys_tmp5007;
	wire signed [31:0] w_sys_tmp5011;
	wire signed [31:0] w_sys_tmp5012;
	wire signed [31:0] w_sys_tmp5016;
	wire signed [31:0] w_sys_tmp5017;
	wire signed [31:0] w_sys_tmp5021;
	wire signed [31:0] w_sys_tmp5022;
	wire signed [31:0] w_sys_tmp5026;
	wire signed [31:0] w_sys_tmp5027;
	wire signed [31:0] w_sys_tmp5031;
	wire signed [31:0] w_sys_tmp5032;
	wire signed [31:0] w_sys_tmp5036;
	wire signed [31:0] w_sys_tmp5037;
	wire signed [31:0] w_sys_tmp5041;
	wire signed [31:0] w_sys_tmp5042;
	wire signed [31:0] w_sys_tmp5046;
	wire signed [31:0] w_sys_tmp5047;
	wire signed [31:0] w_sys_tmp5051;
	wire signed [31:0] w_sys_tmp5052;
	wire signed [31:0] w_sys_tmp5056;
	wire signed [31:0] w_sys_tmp5057;
	wire signed [31:0] w_sys_tmp5061;
	wire signed [31:0] w_sys_tmp5062;
	wire signed [31:0] w_sys_tmp5066;
	wire signed [31:0] w_sys_tmp5067;
	wire signed [31:0] w_sys_tmp5071;
	wire signed [31:0] w_sys_tmp5072;
	wire signed [31:0] w_sys_tmp5076;
	wire signed [31:0] w_sys_tmp5077;
	wire signed [31:0] w_sys_tmp5081;
	wire signed [31:0] w_sys_tmp5082;
	wire signed [31:0] w_sys_tmp5086;
	wire signed [31:0] w_sys_tmp5087;
	wire signed [31:0] w_sys_tmp5091;
	wire signed [31:0] w_sys_tmp5092;
	wire signed [31:0] w_sys_tmp5096;
	wire signed [31:0] w_sys_tmp5097;
	wire signed [31:0] w_sys_tmp5101;
	wire signed [31:0] w_sys_tmp5102;
	wire signed [31:0] w_sys_tmp5106;
	wire signed [31:0] w_sys_tmp5107;
	wire signed [31:0] w_sys_tmp5111;
	wire signed [31:0] w_sys_tmp5112;
	wire signed [31:0] w_sys_tmp5116;
	wire signed [31:0] w_sys_tmp5117;
	wire signed [31:0] w_sys_tmp5121;
	wire signed [31:0] w_sys_tmp5122;
	wire signed [31:0] w_sys_tmp5126;
	wire signed [31:0] w_sys_tmp5127;
	wire signed [31:0] w_sys_tmp5131;
	wire signed [31:0] w_sys_tmp5132;
	wire signed [31:0] w_sys_tmp5136;
	wire signed [31:0] w_sys_tmp5137;
	wire signed [31:0] w_sys_tmp5141;
	wire signed [31:0] w_sys_tmp5142;
	wire signed [31:0] w_sys_tmp5146;
	wire signed [31:0] w_sys_tmp5147;
	wire signed [31:0] w_sys_tmp5151;
	wire signed [31:0] w_sys_tmp5152;
	wire signed [31:0] w_sys_tmp5156;
	wire signed [31:0] w_sys_tmp5157;
	wire signed [31:0] w_sys_tmp5161;
	wire signed [31:0] w_sys_tmp5162;
	wire signed [31:0] w_sys_tmp5166;
	wire signed [31:0] w_sys_tmp5167;
	wire signed [31:0] w_sys_tmp5171;
	wire signed [31:0] w_sys_tmp5172;
	wire signed [31:0] w_sys_tmp5176;
	wire signed [31:0] w_sys_tmp5177;
	wire signed [31:0] w_sys_tmp5181;
	wire signed [31:0] w_sys_tmp5182;
	wire signed [31:0] w_sys_tmp5186;
	wire signed [31:0] w_sys_tmp5187;
	wire signed [31:0] w_sys_tmp5191;
	wire signed [31:0] w_sys_tmp5192;
	wire signed [31:0] w_sys_tmp5196;
	wire signed [31:0] w_sys_tmp5197;
	wire signed [31:0] w_sys_tmp5201;
	wire signed [31:0] w_sys_tmp5202;
	wire signed [31:0] w_sys_tmp5206;
	wire signed [31:0] w_sys_tmp5207;
	wire signed [31:0] w_sys_tmp5211;
	wire signed [31:0] w_sys_tmp5212;
	wire signed [31:0] w_sys_tmp5216;
	wire signed [31:0] w_sys_tmp5217;
	wire signed [31:0] w_sys_tmp5221;
	wire signed [31:0] w_sys_tmp5222;
	wire signed [31:0] w_sys_tmp5226;
	wire signed [31:0] w_sys_tmp5227;
	wire signed [31:0] w_sys_tmp5231;
	wire signed [31:0] w_sys_tmp5232;
	wire signed [31:0] w_sys_tmp5236;
	wire signed [31:0] w_sys_tmp5237;
	wire signed [31:0] w_sys_tmp5241;
	wire signed [31:0] w_sys_tmp5242;
	wire signed [31:0] w_sys_tmp5246;
	wire signed [31:0] w_sys_tmp5247;
	wire signed [31:0] w_sys_tmp5251;
	wire signed [31:0] w_sys_tmp5252;
	wire signed [31:0] w_sys_tmp5256;
	wire signed [31:0] w_sys_tmp5257;
	wire signed [31:0] w_sys_tmp5261;
	wire signed [31:0] w_sys_tmp5262;
	wire signed [31:0] w_sys_tmp5266;
	wire signed [31:0] w_sys_tmp5267;
	wire signed [31:0] w_sys_tmp5271;
	wire signed [31:0] w_sys_tmp5272;
	wire signed [31:0] w_sys_tmp5276;
	wire signed [31:0] w_sys_tmp5277;
	wire signed [31:0] w_sys_tmp5281;
	wire signed [31:0] w_sys_tmp5282;
	wire signed [31:0] w_sys_tmp5286;
	wire signed [31:0] w_sys_tmp5287;
	wire signed [31:0] w_sys_tmp5291;
	wire signed [31:0] w_sys_tmp5292;
	wire signed [31:0] w_sys_tmp5296;
	wire signed [31:0] w_sys_tmp5297;
	wire signed [31:0] w_sys_tmp5301;
	wire signed [31:0] w_sys_tmp5302;
	wire signed [31:0] w_sys_tmp5306;
	wire signed [31:0] w_sys_tmp5307;
	wire signed [31:0] w_sys_tmp5311;
	wire signed [31:0] w_sys_tmp5312;
	wire signed [31:0] w_sys_tmp5316;
	wire signed [31:0] w_sys_tmp5317;
	wire signed [31:0] w_sys_tmp5321;
	wire signed [31:0] w_sys_tmp5322;
	wire signed [31:0] w_sys_tmp5326;
	wire signed [31:0] w_sys_tmp5327;
	wire signed [31:0] w_sys_tmp5331;
	wire signed [31:0] w_sys_tmp5332;
	wire signed [31:0] w_sys_tmp5336;
	wire signed [31:0] w_sys_tmp5337;
	wire signed [31:0] w_sys_tmp5341;
	wire signed [31:0] w_sys_tmp5342;
	wire signed [31:0] w_sys_tmp5346;
	wire signed [31:0] w_sys_tmp5347;
	wire signed [31:0] w_sys_tmp5351;
	wire signed [31:0] w_sys_tmp5352;
	wire signed [31:0] w_sys_tmp5356;
	wire signed [31:0] w_sys_tmp5357;
	wire signed [31:0] w_sys_tmp5361;
	wire signed [31:0] w_sys_tmp5362;
	wire signed [31:0] w_sys_tmp5366;
	wire signed [31:0] w_sys_tmp5367;
	wire signed [31:0] w_sys_tmp5371;
	wire signed [31:0] w_sys_tmp5372;
	wire signed [31:0] w_sys_tmp5376;
	wire signed [31:0] w_sys_tmp5377;
	wire signed [31:0] w_sys_tmp5381;
	wire signed [31:0] w_sys_tmp5382;
	wire signed [31:0] w_sys_tmp5386;
	wire signed [31:0] w_sys_tmp5387;
	wire signed [31:0] w_sys_tmp5391;
	wire signed [31:0] w_sys_tmp5392;
	wire signed [31:0] w_sys_tmp5396;
	wire signed [31:0] w_sys_tmp5397;
	wire signed [31:0] w_sys_tmp5401;
	wire signed [31:0] w_sys_tmp5402;
	wire signed [31:0] w_sys_tmp5406;
	wire signed [31:0] w_sys_tmp5407;
	wire signed [31:0] w_sys_tmp5411;
	wire signed [31:0] w_sys_tmp5412;
	wire signed [31:0] w_sys_tmp5416;
	wire signed [31:0] w_sys_tmp5417;
	wire signed [31:0] w_sys_tmp5421;
	wire signed [31:0] w_sys_tmp5422;
	wire signed [31:0] w_sys_tmp5426;
	wire signed [31:0] w_sys_tmp5427;
	wire signed [31:0] w_sys_tmp5431;
	wire signed [31:0] w_sys_tmp5432;
	wire signed [31:0] w_sys_tmp5436;
	wire signed [31:0] w_sys_tmp5437;
	wire signed [31:0] w_sys_tmp5441;
	wire signed [31:0] w_sys_tmp5442;
	wire signed [31:0] w_sys_tmp5446;
	wire signed [31:0] w_sys_tmp5447;
	wire signed [31:0] w_sys_tmp5451;
	wire signed [31:0] w_sys_tmp5452;
	wire signed [31:0] w_sys_tmp5456;
	wire signed [31:0] w_sys_tmp5457;
	wire signed [31:0] w_sys_tmp5461;
	wire signed [31:0] w_sys_tmp5462;
	wire signed [31:0] w_sys_tmp5466;
	wire signed [31:0] w_sys_tmp5467;
	wire signed [31:0] w_sys_tmp5471;
	wire signed [31:0] w_sys_tmp5472;
	wire signed [31:0] w_sys_tmp5476;
	wire signed [31:0] w_sys_tmp5477;
	wire signed [31:0] w_sys_tmp5481;
	wire signed [31:0] w_sys_tmp5482;
	wire signed [31:0] w_sys_tmp5486;
	wire signed [31:0] w_sys_tmp5487;
	wire signed [31:0] w_sys_tmp5491;
	wire signed [31:0] w_sys_tmp5492;
	wire signed [31:0] w_sys_tmp5496;
	wire signed [31:0] w_sys_tmp5497;
	wire signed [31:0] w_sys_tmp5501;
	wire signed [31:0] w_sys_tmp5502;
	wire signed [31:0] w_sys_tmp5506;
	wire signed [31:0] w_sys_tmp5507;
	wire signed [31:0] w_sys_tmp5511;
	wire signed [31:0] w_sys_tmp5512;
	wire signed [31:0] w_sys_tmp5516;
	wire signed [31:0] w_sys_tmp5517;
	wire signed [31:0] w_sys_tmp5521;
	wire signed [31:0] w_sys_tmp5522;
	wire signed [31:0] w_sys_tmp5526;
	wire signed [31:0] w_sys_tmp5527;
	wire signed [31:0] w_sys_tmp5531;
	wire signed [31:0] w_sys_tmp5532;
	wire signed [31:0] w_sys_tmp5536;
	wire signed [31:0] w_sys_tmp5537;
	wire signed [31:0] w_sys_tmp5541;
	wire signed [31:0] w_sys_tmp5542;
	wire signed [31:0] w_sys_tmp5546;
	wire signed [31:0] w_sys_tmp5547;
	wire signed [31:0] w_sys_tmp5551;
	wire signed [31:0] w_sys_tmp5552;
	wire signed [31:0] w_sys_tmp5556;
	wire signed [31:0] w_sys_tmp5557;
	wire signed [31:0] w_sys_tmp5561;
	wire signed [31:0] w_sys_tmp5562;
	wire signed [31:0] w_sys_tmp5566;
	wire signed [31:0] w_sys_tmp5567;
	wire signed [31:0] w_sys_tmp5571;
	wire signed [31:0] w_sys_tmp5572;
	wire signed [31:0] w_sys_tmp5576;
	wire signed [31:0] w_sys_tmp5577;
	wire signed [31:0] w_sys_tmp5581;
	wire signed [31:0] w_sys_tmp5582;
	wire signed [31:0] w_sys_tmp5586;
	wire signed [31:0] w_sys_tmp5587;
	wire signed [31:0] w_sys_tmp5591;
	wire signed [31:0] w_sys_tmp5592;
	wire signed [31:0] w_sys_tmp5596;
	wire signed [31:0] w_sys_tmp5597;
	wire signed [31:0] w_sys_tmp5601;
	wire signed [31:0] w_sys_tmp5602;
	wire signed [31:0] w_sys_tmp5606;
	wire signed [31:0] w_sys_tmp5607;
	wire signed [31:0] w_sys_tmp5611;
	wire signed [31:0] w_sys_tmp5612;
	wire signed [31:0] w_sys_tmp5616;
	wire signed [31:0] w_sys_tmp5617;
	wire signed [31:0] w_sys_tmp5621;
	wire signed [31:0] w_sys_tmp5622;
	wire signed [31:0] w_sys_tmp5626;
	wire signed [31:0] w_sys_tmp5627;
	wire signed [31:0] w_sys_tmp5631;
	wire signed [31:0] w_sys_tmp5632;
	wire signed [31:0] w_sys_tmp5636;
	wire signed [31:0] w_sys_tmp5637;
	wire signed [31:0] w_sys_tmp5641;
	wire signed [31:0] w_sys_tmp5642;
	wire signed [31:0] w_sys_tmp5646;
	wire signed [31:0] w_sys_tmp5647;
	wire signed [31:0] w_sys_tmp5651;
	wire signed [31:0] w_sys_tmp5652;
	wire signed [31:0] w_sys_tmp5656;
	wire signed [31:0] w_sys_tmp5657;
	wire signed [31:0] w_sys_tmp5661;
	wire signed [31:0] w_sys_tmp5662;
	wire signed [31:0] w_sys_tmp5666;
	wire signed [31:0] w_sys_tmp5667;
	wire signed [31:0] w_sys_tmp5671;
	wire signed [31:0] w_sys_tmp5672;
	wire signed [31:0] w_sys_tmp5676;
	wire signed [31:0] w_sys_tmp5677;
	wire signed [31:0] w_sys_tmp5681;
	wire signed [31:0] w_sys_tmp5682;
	wire signed [31:0] w_sys_tmp5686;
	wire signed [31:0] w_sys_tmp5687;
	wire signed [31:0] w_sys_tmp5691;
	wire signed [31:0] w_sys_tmp5692;
	wire signed [31:0] w_sys_tmp5696;
	wire signed [31:0] w_sys_tmp5697;
	wire signed [31:0] w_sys_tmp5701;
	wire signed [31:0] w_sys_tmp5702;
	wire signed [31:0] w_sys_tmp5706;
	wire signed [31:0] w_sys_tmp5707;
	wire signed [31:0] w_sys_tmp5711;
	wire signed [31:0] w_sys_tmp5712;
	wire signed [31:0] w_sys_tmp5716;
	wire signed [31:0] w_sys_tmp5717;
	wire signed [31:0] w_sys_tmp5721;
	wire signed [31:0] w_sys_tmp5722;
	wire signed [31:0] w_sys_tmp5726;
	wire signed [31:0] w_sys_tmp5727;
	wire signed [31:0] w_sys_tmp5731;
	wire signed [31:0] w_sys_tmp5732;
	wire signed [31:0] w_sys_tmp5736;
	wire signed [31:0] w_sys_tmp5737;
	wire signed [31:0] w_sys_tmp5741;
	wire signed [31:0] w_sys_tmp5742;
	wire signed [31:0] w_sys_tmp5746;
	wire signed [31:0] w_sys_tmp5747;
	wire signed [31:0] w_sys_tmp5751;
	wire signed [31:0] w_sys_tmp5752;
	wire signed [31:0] w_sys_tmp5756;
	wire signed [31:0] w_sys_tmp5757;
	wire signed [31:0] w_sys_tmp5761;
	wire signed [31:0] w_sys_tmp5762;
	wire signed [31:0] w_sys_tmp5766;
	wire signed [31:0] w_sys_tmp5767;
	wire signed [31:0] w_sys_tmp5771;
	wire signed [31:0] w_sys_tmp5772;
	wire signed [31:0] w_sys_tmp5776;
	wire signed [31:0] w_sys_tmp5777;
	wire signed [31:0] w_sys_tmp5781;
	wire signed [31:0] w_sys_tmp5782;
	wire signed [31:0] w_sys_tmp5786;
	wire signed [31:0] w_sys_tmp5787;
	wire signed [31:0] w_sys_tmp5791;
	wire signed [31:0] w_sys_tmp5792;
	wire signed [31:0] w_sys_tmp5796;
	wire signed [31:0] w_sys_tmp5797;
	wire signed [31:0] w_sys_tmp5801;
	wire signed [31:0] w_sys_tmp5802;
	wire signed [31:0] w_sys_tmp5806;
	wire signed [31:0] w_sys_tmp5807;
	wire signed [31:0] w_sys_tmp5811;
	wire signed [31:0] w_sys_tmp5812;
	wire signed [31:0] w_sys_tmp5816;
	wire signed [31:0] w_sys_tmp5817;
	wire signed [31:0] w_sys_tmp5821;
	wire signed [31:0] w_sys_tmp5822;
	wire signed [31:0] w_sys_tmp5826;
	wire signed [31:0] w_sys_tmp5827;
	wire signed [31:0] w_sys_tmp5831;
	wire signed [31:0] w_sys_tmp5832;
	wire signed [31:0] w_sys_tmp5836;
	wire signed [31:0] w_sys_tmp5837;
	wire signed [31:0] w_sys_tmp5841;
	wire signed [31:0] w_sys_tmp5842;
	wire signed [31:0] w_sys_tmp5846;
	wire signed [31:0] w_sys_tmp5847;
	wire signed [31:0] w_sys_tmp5851;
	wire signed [31:0] w_sys_tmp5852;
	wire signed [31:0] w_sys_tmp5856;
	wire signed [31:0] w_sys_tmp5857;
	wire signed [31:0] w_sys_tmp5861;
	wire signed [31:0] w_sys_tmp5862;
	wire signed [31:0] w_sys_tmp5866;
	wire signed [31:0] w_sys_tmp5867;
	wire signed [31:0] w_sys_tmp5871;
	wire signed [31:0] w_sys_tmp5872;
	wire signed [31:0] w_sys_tmp5876;
	wire signed [31:0] w_sys_tmp5877;
	wire signed [31:0] w_sys_tmp5881;
	wire signed [31:0] w_sys_tmp5882;
	wire signed [31:0] w_sys_tmp5886;
	wire signed [31:0] w_sys_tmp5887;
	wire signed [31:0] w_sys_tmp5891;
	wire signed [31:0] w_sys_tmp5892;
	wire signed [31:0] w_sys_tmp5896;
	wire signed [31:0] w_sys_tmp5897;
	wire signed [31:0] w_sys_tmp5901;
	wire signed [31:0] w_sys_tmp5902;
	wire signed [31:0] w_sys_tmp5906;
	wire signed [31:0] w_sys_tmp5907;
	wire signed [31:0] w_sys_tmp5911;
	wire signed [31:0] w_sys_tmp5912;
	wire signed [31:0] w_sys_tmp5916;
	wire signed [31:0] w_sys_tmp5917;
	wire signed [31:0] w_sys_tmp5921;
	wire signed [31:0] w_sys_tmp5922;
	wire signed [31:0] w_sys_tmp5926;
	wire signed [31:0] w_sys_tmp5927;
	wire signed [31:0] w_sys_tmp5931;
	wire signed [31:0] w_sys_tmp5932;
	wire signed [31:0] w_sys_tmp5936;
	wire signed [31:0] w_sys_tmp5937;
	wire signed [31:0] w_sys_tmp5941;
	wire signed [31:0] w_sys_tmp5942;
	wire signed [31:0] w_sys_tmp5946;
	wire signed [31:0] w_sys_tmp5947;
	wire signed [31:0] w_sys_tmp5951;
	wire signed [31:0] w_sys_tmp5952;
	wire signed [31:0] w_sys_tmp5956;
	wire signed [31:0] w_sys_tmp5957;
	wire signed [31:0] w_sys_tmp5961;
	wire signed [31:0] w_sys_tmp5962;
	wire signed [31:0] w_sys_tmp5966;
	wire signed [31:0] w_sys_tmp5967;
	wire signed [31:0] w_sys_tmp5971;
	wire signed [31:0] w_sys_tmp5972;
	wire signed [31:0] w_sys_tmp5976;
	wire signed [31:0] w_sys_tmp5977;
	wire signed [31:0] w_sys_tmp5981;
	wire signed [31:0] w_sys_tmp5982;
	wire signed [31:0] w_sys_tmp5986;
	wire signed [31:0] w_sys_tmp5987;
	wire signed [31:0] w_sys_tmp5991;
	wire signed [31:0] w_sys_tmp5992;
	wire signed [31:0] w_sys_tmp5996;
	wire signed [31:0] w_sys_tmp5997;
	wire signed [31:0] w_sys_tmp6001;
	wire signed [31:0] w_sys_tmp6002;
	wire signed [31:0] w_sys_tmp6006;
	wire signed [31:0] w_sys_tmp6007;
	wire signed [31:0] w_sys_tmp6011;
	wire signed [31:0] w_sys_tmp6012;
	wire signed [31:0] w_sys_tmp6016;
	wire signed [31:0] w_sys_tmp6017;
	wire signed [31:0] w_sys_tmp6021;
	wire signed [31:0] w_sys_tmp6022;
	wire signed [31:0] w_sys_tmp6026;
	wire signed [31:0] w_sys_tmp6027;
	wire signed [31:0] w_sys_tmp6031;
	wire signed [31:0] w_sys_tmp6032;
	wire signed [31:0] w_sys_tmp6036;
	wire signed [31:0] w_sys_tmp6037;
	wire signed [31:0] w_sys_tmp6041;
	wire signed [31:0] w_sys_tmp6042;
	wire signed [31:0] w_sys_tmp6046;
	wire signed [31:0] w_sys_tmp6047;
	wire signed [31:0] w_sys_tmp6051;
	wire signed [31:0] w_sys_tmp6052;
	wire signed [31:0] w_sys_tmp6056;
	wire signed [31:0] w_sys_tmp6057;
	wire signed [31:0] w_sys_tmp6061;
	wire signed [31:0] w_sys_tmp6062;
	wire signed [31:0] w_sys_tmp6066;
	wire signed [31:0] w_sys_tmp6067;
	wire signed [31:0] w_sys_tmp6071;
	wire signed [31:0] w_sys_tmp6072;
	wire signed [31:0] w_sys_tmp6075;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 5'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 9'h1);
	assign w_fld_u_0_addr_0 = 15'sh0;
	assign w_fld_u_0_datain_0 = 32'h0;
	assign w_fld_u_0_r_w_0 = 1'h0;
	assign w_fld_u_0_ce_0 = w_sys_ce;
	assign w_fld_u_0_ce_1 = w_sys_ce;
	assign w_sub09_u_addr = ( (|r_sys_processing_methodID) ? r_sub09_u_addr : 15'sh0 ) ;
	assign w_sub09_u_datain = ( (|r_sys_processing_methodID) ? r_sub09_u_datain : 32'h0 ) ;
	assign w_sub09_u_r_w = ( (|r_sys_processing_methodID) ? r_sub09_u_r_w : 1'h0 ) ;
	assign w_sub09_result_addr = ( (|r_sys_processing_methodID) ? r_sub09_result_addr : 15'sh0 ) ;
	assign w_sub09_result_datain = ( (|r_sys_processing_methodID) ? r_sub09_result_datain : 32'h0 ) ;
	assign w_sub09_result_r_w = ( (|r_sys_processing_methodID) ? r_sub09_result_r_w : 1'h0 ) ;
	assign w_sub08_u_addr = ( (|r_sys_processing_methodID) ? r_sub08_u_addr : 15'sh0 ) ;
	assign w_sub08_u_datain = ( (|r_sys_processing_methodID) ? r_sub08_u_datain : 32'h0 ) ;
	assign w_sub08_u_r_w = ( (|r_sys_processing_methodID) ? r_sub08_u_r_w : 1'h0 ) ;
	assign w_sub08_result_addr = ( (|r_sys_processing_methodID) ? r_sub08_result_addr : 15'sh0 ) ;
	assign w_sub08_result_datain = ( (|r_sys_processing_methodID) ? r_sub08_result_datain : 32'h0 ) ;
	assign w_sub08_result_r_w = ( (|r_sys_processing_methodID) ? r_sub08_result_r_w : 1'h0 ) ;
	assign w_sub12_u_addr = ( (|r_sys_processing_methodID) ? r_sub12_u_addr : 15'sh0 ) ;
	assign w_sub12_u_datain = ( (|r_sys_processing_methodID) ? r_sub12_u_datain : 32'h0 ) ;
	assign w_sub12_u_r_w = ( (|r_sys_processing_methodID) ? r_sub12_u_r_w : 1'h0 ) ;
	assign w_sub12_result_addr = ( (|r_sys_processing_methodID) ? r_sub12_result_addr : 15'sh0 ) ;
	assign w_sub12_result_datain = ( (|r_sys_processing_methodID) ? r_sub12_result_datain : 32'h0 ) ;
	assign w_sub12_result_r_w = ( (|r_sys_processing_methodID) ? r_sub12_result_r_w : 1'h0 ) ;
	assign w_sub03_u_addr = ( (|r_sys_processing_methodID) ? r_sub03_u_addr : 15'sh0 ) ;
	assign w_sub03_u_datain = ( (|r_sys_processing_methodID) ? r_sub03_u_datain : 32'h0 ) ;
	assign w_sub03_u_r_w = ( (|r_sys_processing_methodID) ? r_sub03_u_r_w : 1'h0 ) ;
	assign w_sub03_result_addr = ( (|r_sys_processing_methodID) ? r_sub03_result_addr : 15'sh0 ) ;
	assign w_sub03_result_datain = ( (|r_sys_processing_methodID) ? r_sub03_result_datain : 32'h0 ) ;
	assign w_sub03_result_r_w = ( (|r_sys_processing_methodID) ? r_sub03_result_r_w : 1'h0 ) ;
	assign w_sub02_u_addr = ( (|r_sys_processing_methodID) ? r_sub02_u_addr : 15'sh0 ) ;
	assign w_sub02_u_datain = ( (|r_sys_processing_methodID) ? r_sub02_u_datain : 32'h0 ) ;
	assign w_sub02_u_r_w = ( (|r_sys_processing_methodID) ? r_sub02_u_r_w : 1'h0 ) ;
	assign w_sub02_result_addr = ( (|r_sys_processing_methodID) ? r_sub02_result_addr : 15'sh0 ) ;
	assign w_sub02_result_datain = ( (|r_sys_processing_methodID) ? r_sub02_result_datain : 32'h0 ) ;
	assign w_sub02_result_r_w = ( (|r_sys_processing_methodID) ? r_sub02_result_r_w : 1'h0 ) ;
	assign w_sub11_u_addr = ( (|r_sys_processing_methodID) ? r_sub11_u_addr : 15'sh0 ) ;
	assign w_sub11_u_datain = ( (|r_sys_processing_methodID) ? r_sub11_u_datain : 32'h0 ) ;
	assign w_sub11_u_r_w = ( (|r_sys_processing_methodID) ? r_sub11_u_r_w : 1'h0 ) ;
	assign w_sub11_result_addr = ( (|r_sys_processing_methodID) ? r_sub11_result_addr : 15'sh0 ) ;
	assign w_sub11_result_datain = ( (|r_sys_processing_methodID) ? r_sub11_result_datain : 32'h0 ) ;
	assign w_sub11_result_r_w = ( (|r_sys_processing_methodID) ? r_sub11_result_r_w : 1'h0 ) ;
	assign w_sub14_u_addr = ( (|r_sys_processing_methodID) ? r_sub14_u_addr : 15'sh0 ) ;
	assign w_sub14_u_datain = ( (|r_sys_processing_methodID) ? r_sub14_u_datain : 32'h0 ) ;
	assign w_sub14_u_r_w = ( (|r_sys_processing_methodID) ? r_sub14_u_r_w : 1'h0 ) ;
	assign w_sub14_result_addr = ( (|r_sys_processing_methodID) ? r_sub14_result_addr : 15'sh0 ) ;
	assign w_sub14_result_datain = ( (|r_sys_processing_methodID) ? r_sub14_result_datain : 32'h0 ) ;
	assign w_sub14_result_r_w = ( (|r_sys_processing_methodID) ? r_sub14_result_r_w : 1'h0 ) ;
	assign w_sub01_u_addr = ( (|r_sys_processing_methodID) ? r_sub01_u_addr : 15'sh0 ) ;
	assign w_sub01_u_datain = ( (|r_sys_processing_methodID) ? r_sub01_u_datain : 32'h0 ) ;
	assign w_sub01_u_r_w = ( (|r_sys_processing_methodID) ? r_sub01_u_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 15'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub13_u_addr = ( (|r_sys_processing_methodID) ? r_sub13_u_addr : 15'sh0 ) ;
	assign w_sub13_u_datain = ( (|r_sys_processing_methodID) ? r_sub13_u_datain : 32'h0 ) ;
	assign w_sub13_u_r_w = ( (|r_sys_processing_methodID) ? r_sub13_u_r_w : 1'h0 ) ;
	assign w_sub13_result_addr = ( (|r_sys_processing_methodID) ? r_sub13_result_addr : 15'sh0 ) ;
	assign w_sub13_result_datain = ( (|r_sys_processing_methodID) ? r_sub13_result_datain : 32'h0 ) ;
	assign w_sub13_result_r_w = ( (|r_sys_processing_methodID) ? r_sub13_result_r_w : 1'h0 ) ;
	assign w_sub00_u_addr = ( (|r_sys_processing_methodID) ? r_sub00_u_addr : 15'sh0 ) ;
	assign w_sub00_u_datain = ( (|r_sys_processing_methodID) ? r_sub00_u_datain : 32'h0 ) ;
	assign w_sub00_u_r_w = ( (|r_sys_processing_methodID) ? r_sub00_u_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 15'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sub07_u_addr = ( (|r_sys_processing_methodID) ? r_sub07_u_addr : 15'sh0 ) ;
	assign w_sub07_u_datain = ( (|r_sys_processing_methodID) ? r_sub07_u_datain : 32'h0 ) ;
	assign w_sub07_u_r_w = ( (|r_sys_processing_methodID) ? r_sub07_u_r_w : 1'h0 ) ;
	assign w_sub07_result_addr = ( (|r_sys_processing_methodID) ? r_sub07_result_addr : 15'sh0 ) ;
	assign w_sub07_result_datain = ( (|r_sys_processing_methodID) ? r_sub07_result_datain : 32'h0 ) ;
	assign w_sub07_result_r_w = ( (|r_sys_processing_methodID) ? r_sub07_result_r_w : 1'h0 ) ;
	assign w_sub06_u_addr = ( (|r_sys_processing_methodID) ? r_sub06_u_addr : 15'sh0 ) ;
	assign w_sub06_u_datain = ( (|r_sys_processing_methodID) ? r_sub06_u_datain : 32'h0 ) ;
	assign w_sub06_u_r_w = ( (|r_sys_processing_methodID) ? r_sub06_u_r_w : 1'h0 ) ;
	assign w_sub06_result_addr = ( (|r_sys_processing_methodID) ? r_sub06_result_addr : 15'sh0 ) ;
	assign w_sub06_result_datain = ( (|r_sys_processing_methodID) ? r_sub06_result_datain : 32'h0 ) ;
	assign w_sub06_result_r_w = ( (|r_sys_processing_methodID) ? r_sub06_result_r_w : 1'h0 ) ;
	assign w_sub15_u_addr = ( (|r_sys_processing_methodID) ? r_sub15_u_addr : 15'sh0 ) ;
	assign w_sub15_u_datain = ( (|r_sys_processing_methodID) ? r_sub15_u_datain : 32'h0 ) ;
	assign w_sub15_u_r_w = ( (|r_sys_processing_methodID) ? r_sub15_u_r_w : 1'h0 ) ;
	assign w_sub15_result_addr = ( (|r_sys_processing_methodID) ? r_sub15_result_addr : 15'sh0 ) ;
	assign w_sub15_result_datain = ( (|r_sys_processing_methodID) ? r_sub15_result_datain : 32'h0 ) ;
	assign w_sub15_result_r_w = ( (|r_sys_processing_methodID) ? r_sub15_result_r_w : 1'h0 ) ;
	assign w_sub05_u_addr = ( (|r_sys_processing_methodID) ? r_sub05_u_addr : 15'sh0 ) ;
	assign w_sub05_u_datain = ( (|r_sys_processing_methodID) ? r_sub05_u_datain : 32'h0 ) ;
	assign w_sub05_u_r_w = ( (|r_sys_processing_methodID) ? r_sub05_u_r_w : 1'h0 ) ;
	assign w_sub05_result_addr = ( (|r_sys_processing_methodID) ? r_sub05_result_addr : 15'sh0 ) ;
	assign w_sub05_result_datain = ( (|r_sys_processing_methodID) ? r_sub05_result_datain : 32'h0 ) ;
	assign w_sub05_result_r_w = ( (|r_sys_processing_methodID) ? r_sub05_result_r_w : 1'h0 ) ;
	assign w_sub04_u_addr = ( (|r_sys_processing_methodID) ? r_sub04_u_addr : 15'sh0 ) ;
	assign w_sub04_u_datain = ( (|r_sys_processing_methodID) ? r_sub04_u_datain : 32'h0 ) ;
	assign w_sub04_u_r_w = ( (|r_sys_processing_methodID) ? r_sub04_u_r_w : 1'h0 ) ;
	assign w_sub04_result_addr = ( (|r_sys_processing_methodID) ? r_sub04_result_addr : 15'sh0 ) ;
	assign w_sub04_result_datain = ( (|r_sys_processing_methodID) ? r_sub04_result_datain : 32'h0 ) ;
	assign w_sub04_result_r_w = ( (|r_sys_processing_methodID) ? r_sub04_result_r_w : 1'h0 ) ;
	assign w_sub10_u_addr = ( (|r_sys_processing_methodID) ? r_sub10_u_addr : 15'sh0 ) ;
	assign w_sub10_u_datain = ( (|r_sys_processing_methodID) ? r_sub10_u_datain : 32'h0 ) ;
	assign w_sub10_u_r_w = ( (|r_sys_processing_methodID) ? r_sub10_u_r_w : 1'h0 ) ;
	assign w_sub10_result_addr = ( (|r_sys_processing_methodID) ? r_sub10_result_addr : 15'sh0 ) ;
	assign w_sub10_result_datain = ( (|r_sys_processing_methodID) ? r_sub10_result_datain : 32'h0 ) ;
	assign w_sub10_result_r_w = ( (|r_sys_processing_methodID) ? r_sub10_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh00000081;
	assign w_sys_tmp3 = ( !w_sys_tmp4 );
	assign w_sys_tmp4 = (r_run_my_21 < r_run_k_17);
	assign w_sys_tmp5 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp6 = ( !w_sys_tmp7 );
	assign w_sys_tmp7 = (r_run_mx_20 < r_run_j_18);
	assign w_sys_tmp10 = (w_sys_tmp11 + r_run_k_17);
	assign w_sys_tmp11 = (r_run_j_18 * w_sys_tmp12);
	assign w_sys_tmp12 = 32'sh00000081;
	assign w_sys_tmp13 = 32'h0;
	assign w_sys_tmp14 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp51 = ( !w_sys_tmp52 );
	assign w_sys_tmp52 = (r_run_nlast_22 < r_run_n_19);
	assign w_sys_tmp53 = (r_run_n_19 + w_sys_intOne);
	assign w_sys_tmp54 = ( !w_sys_tmp55 );
	assign w_sys_tmp55 = (r_run_my_21 < r_run_j_18);
	assign w_sys_tmp58 = (w_sys_tmp59 + r_run_j_18);
	assign w_sys_tmp59 = 32'sh00000081;
	assign w_sys_tmp60 = 32'h3f000000;
	assign w_sys_tmp62 = (w_sys_tmp63 + r_run_copy2_j_25);
	assign w_sys_tmp63 = 32'sh00004101;
	assign w_sys_tmp64 = 32'h0;
	assign w_sys_tmp66 = (w_sys_tmp67 + w_sys_intOne);
	assign w_sys_tmp67 = (r_run_copy1_j_24 * w_sys_tmp59);
	assign w_sys_tmp69 = 32'h3f800000;
	assign w_sys_tmp71 = (w_sys_tmp72 + r_run_my_21);
	assign w_sys_tmp72 = (r_run_copy0_j_23 * w_sys_tmp59);
	assign w_sys_tmp75 = (r_run_copy0_j_23 + w_sys_intOne);
	assign w_sys_tmp76 = (r_run_copy1_j_24 + w_sys_intOne);
	assign w_sys_tmp77 = (r_run_copy2_j_25 + w_sys_intOne);
	assign w_sys_tmp78 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp211 = ( !w_sys_tmp212 );
	assign w_sys_tmp212 = (w_sys_tmp213 < r_run_k_17);
	assign w_sys_tmp213 = 32'sh00000021;
	assign w_sys_tmp216 = (w_sys_tmp217 + r_run_k_17);
	assign w_sys_tmp217 = 32'sh00000081;
	assign w_sys_tmp218 = w_fld_u_0_dataout_1;
	assign w_sys_tmp222 = (w_sys_tmp223 + r_run_k_17);
	assign w_sys_tmp223 = 32'sh00000102;
	assign w_sys_tmp228 = (w_sys_tmp229 + r_run_k_17);
	assign w_sys_tmp229 = 32'sh00000183;
	assign w_sys_tmp234 = (w_sys_tmp235 + r_run_k_17);
	assign w_sys_tmp235 = 32'sh00000204;
	assign w_sys_tmp240 = (w_sys_tmp241 + r_run_k_17);
	assign w_sys_tmp241 = 32'sh00000285;
	assign w_sys_tmp246 = (w_sys_tmp247 + r_run_k_17);
	assign w_sys_tmp247 = 32'sh00000306;
	assign w_sys_tmp252 = (w_sys_tmp253 + r_run_k_17);
	assign w_sys_tmp253 = 32'sh00000387;
	assign w_sys_tmp258 = (w_sys_tmp259 + r_run_k_17);
	assign w_sys_tmp259 = 32'sh00000408;
	assign w_sys_tmp264 = (w_sys_tmp265 + r_run_k_17);
	assign w_sys_tmp265 = 32'sh00000489;
	assign w_sys_tmp270 = (w_sys_tmp271 + r_run_k_17);
	assign w_sys_tmp271 = 32'sh0000050a;
	assign w_sys_tmp276 = (w_sys_tmp277 + r_run_k_17);
	assign w_sys_tmp277 = 32'sh0000058b;
	assign w_sys_tmp282 = (w_sys_tmp283 + r_run_k_17);
	assign w_sys_tmp283 = 32'sh0000060c;
	assign w_sys_tmp288 = (w_sys_tmp289 + r_run_k_17);
	assign w_sys_tmp289 = 32'sh0000068d;
	assign w_sys_tmp294 = (w_sys_tmp295 + r_run_k_17);
	assign w_sys_tmp295 = 32'sh0000070e;
	assign w_sys_tmp300 = (w_sys_tmp301 + r_run_k_17);
	assign w_sys_tmp301 = 32'sh0000078f;
	assign w_sys_tmp306 = (w_sys_tmp307 + r_run_k_17);
	assign w_sys_tmp307 = 32'sh00000810;
	assign w_sys_tmp312 = (w_sys_tmp313 + r_run_k_17);
	assign w_sys_tmp313 = 32'sh00000891;
	assign w_sys_tmp318 = (w_sys_tmp319 + r_run_k_17);
	assign w_sys_tmp319 = 32'sh00000912;
	assign w_sys_tmp324 = (w_sys_tmp325 + r_run_k_17);
	assign w_sys_tmp325 = 32'sh00000993;
	assign w_sys_tmp330 = (w_sys_tmp331 + r_run_k_17);
	assign w_sys_tmp331 = 32'sh00000a14;
	assign w_sys_tmp336 = (w_sys_tmp337 + r_run_k_17);
	assign w_sys_tmp337 = 32'sh00000a95;
	assign w_sys_tmp342 = (w_sys_tmp343 + r_run_k_17);
	assign w_sys_tmp343 = 32'sh00000b16;
	assign w_sys_tmp348 = (w_sys_tmp349 + r_run_k_17);
	assign w_sys_tmp349 = 32'sh00000b97;
	assign w_sys_tmp354 = (w_sys_tmp355 + r_run_k_17);
	assign w_sys_tmp355 = 32'sh00000c18;
	assign w_sys_tmp360 = (w_sys_tmp361 + r_run_k_17);
	assign w_sys_tmp361 = 32'sh00000c99;
	assign w_sys_tmp366 = (w_sys_tmp367 + r_run_k_17);
	assign w_sys_tmp367 = 32'sh00000d1a;
	assign w_sys_tmp372 = (w_sys_tmp373 + r_run_k_17);
	assign w_sys_tmp373 = 32'sh00000d9b;
	assign w_sys_tmp378 = (w_sys_tmp379 + r_run_k_17);
	assign w_sys_tmp379 = 32'sh00000e1c;
	assign w_sys_tmp384 = (w_sys_tmp385 + r_run_k_17);
	assign w_sys_tmp385 = 32'sh00000e9d;
	assign w_sys_tmp390 = (w_sys_tmp391 + r_run_k_17);
	assign w_sys_tmp391 = 32'sh00000f1e;
	assign w_sys_tmp396 = (w_sys_tmp397 + r_run_k_17);
	assign w_sys_tmp397 = 32'sh00000f9f;
	assign w_sys_tmp402 = (w_sys_tmp403 + r_run_k_17);
	assign w_sys_tmp403 = 32'sh00001020;
	assign w_sys_tmp408 = (w_sys_tmp409 + r_run_k_17);
	assign w_sys_tmp409 = 32'sh000010a1;
	assign w_sys_tmp426 = (w_sys_tmp427 + r_run_k_17);
	assign w_sys_tmp427 = 32'sh00001122;
	assign w_sys_tmp432 = (w_sys_tmp433 + r_run_k_17);
	assign w_sys_tmp433 = 32'sh000011a3;
	assign w_sys_tmp438 = (w_sys_tmp439 + r_run_k_17);
	assign w_sys_tmp439 = 32'sh00001224;
	assign w_sys_tmp444 = (w_sys_tmp445 + r_run_k_17);
	assign w_sys_tmp445 = 32'sh000012a5;
	assign w_sys_tmp450 = (w_sys_tmp451 + r_run_k_17);
	assign w_sys_tmp451 = 32'sh00001326;
	assign w_sys_tmp456 = (w_sys_tmp457 + r_run_k_17);
	assign w_sys_tmp457 = 32'sh000013a7;
	assign w_sys_tmp462 = (w_sys_tmp463 + r_run_k_17);
	assign w_sys_tmp463 = 32'sh00001428;
	assign w_sys_tmp468 = (w_sys_tmp469 + r_run_k_17);
	assign w_sys_tmp469 = 32'sh000014a9;
	assign w_sys_tmp474 = (w_sys_tmp475 + r_run_k_17);
	assign w_sys_tmp475 = 32'sh0000152a;
	assign w_sys_tmp480 = (w_sys_tmp481 + r_run_k_17);
	assign w_sys_tmp481 = 32'sh000015ab;
	assign w_sys_tmp486 = (w_sys_tmp487 + r_run_k_17);
	assign w_sys_tmp487 = 32'sh0000162c;
	assign w_sys_tmp492 = (w_sys_tmp493 + r_run_k_17);
	assign w_sys_tmp493 = 32'sh000016ad;
	assign w_sys_tmp498 = (w_sys_tmp499 + r_run_k_17);
	assign w_sys_tmp499 = 32'sh0000172e;
	assign w_sys_tmp504 = (w_sys_tmp505 + r_run_k_17);
	assign w_sys_tmp505 = 32'sh000017af;
	assign w_sys_tmp510 = (w_sys_tmp511 + r_run_k_17);
	assign w_sys_tmp511 = 32'sh00001830;
	assign w_sys_tmp516 = (w_sys_tmp517 + r_run_k_17);
	assign w_sys_tmp517 = 32'sh000018b1;
	assign w_sys_tmp522 = (w_sys_tmp523 + r_run_k_17);
	assign w_sys_tmp523 = 32'sh00001932;
	assign w_sys_tmp528 = (w_sys_tmp529 + r_run_k_17);
	assign w_sys_tmp529 = 32'sh000019b3;
	assign w_sys_tmp534 = (w_sys_tmp535 + r_run_k_17);
	assign w_sys_tmp535 = 32'sh00001a34;
	assign w_sys_tmp540 = (w_sys_tmp541 + r_run_k_17);
	assign w_sys_tmp541 = 32'sh00001ab5;
	assign w_sys_tmp546 = (w_sys_tmp547 + r_run_k_17);
	assign w_sys_tmp547 = 32'sh00001b36;
	assign w_sys_tmp552 = (w_sys_tmp553 + r_run_k_17);
	assign w_sys_tmp553 = 32'sh00001bb7;
	assign w_sys_tmp558 = (w_sys_tmp559 + r_run_k_17);
	assign w_sys_tmp559 = 32'sh00001c38;
	assign w_sys_tmp564 = (w_sys_tmp565 + r_run_k_17);
	assign w_sys_tmp565 = 32'sh00001cb9;
	assign w_sys_tmp570 = (w_sys_tmp571 + r_run_k_17);
	assign w_sys_tmp571 = 32'sh00001d3a;
	assign w_sys_tmp576 = (w_sys_tmp577 + r_run_k_17);
	assign w_sys_tmp577 = 32'sh00001dbb;
	assign w_sys_tmp582 = (w_sys_tmp583 + r_run_k_17);
	assign w_sys_tmp583 = 32'sh00001e3c;
	assign w_sys_tmp588 = (w_sys_tmp589 + r_run_k_17);
	assign w_sys_tmp589 = 32'sh00001ebd;
	assign w_sys_tmp594 = (w_sys_tmp595 + r_run_k_17);
	assign w_sys_tmp595 = 32'sh00001f3e;
	assign w_sys_tmp600 = (w_sys_tmp601 + r_run_k_17);
	assign w_sys_tmp601 = 32'sh00001fbf;
	assign w_sys_tmp606 = (w_sys_tmp607 + r_run_k_17);
	assign w_sys_tmp607 = 32'sh00002040;
	assign w_sys_tmp612 = (w_sys_tmp613 + r_run_k_17);
	assign w_sys_tmp613 = 32'sh000020c1;
	assign w_sys_tmp630 = (w_sys_tmp631 + r_run_k_17);
	assign w_sys_tmp631 = 32'sh00002142;
	assign w_sys_tmp636 = (w_sys_tmp637 + r_run_k_17);
	assign w_sys_tmp637 = 32'sh000021c3;
	assign w_sys_tmp642 = (w_sys_tmp643 + r_run_k_17);
	assign w_sys_tmp643 = 32'sh00002244;
	assign w_sys_tmp648 = (w_sys_tmp649 + r_run_k_17);
	assign w_sys_tmp649 = 32'sh000022c5;
	assign w_sys_tmp654 = (w_sys_tmp655 + r_run_k_17);
	assign w_sys_tmp655 = 32'sh00002346;
	assign w_sys_tmp660 = (w_sys_tmp661 + r_run_k_17);
	assign w_sys_tmp661 = 32'sh000023c7;
	assign w_sys_tmp666 = (w_sys_tmp667 + r_run_k_17);
	assign w_sys_tmp667 = 32'sh00002448;
	assign w_sys_tmp672 = (w_sys_tmp673 + r_run_k_17);
	assign w_sys_tmp673 = 32'sh000024c9;
	assign w_sys_tmp678 = (w_sys_tmp679 + r_run_k_17);
	assign w_sys_tmp679 = 32'sh0000254a;
	assign w_sys_tmp684 = (w_sys_tmp685 + r_run_k_17);
	assign w_sys_tmp685 = 32'sh000025cb;
	assign w_sys_tmp690 = (w_sys_tmp691 + r_run_k_17);
	assign w_sys_tmp691 = 32'sh0000264c;
	assign w_sys_tmp696 = (w_sys_tmp697 + r_run_k_17);
	assign w_sys_tmp697 = 32'sh000026cd;
	assign w_sys_tmp702 = (w_sys_tmp703 + r_run_k_17);
	assign w_sys_tmp703 = 32'sh0000274e;
	assign w_sys_tmp708 = (w_sys_tmp709 + r_run_k_17);
	assign w_sys_tmp709 = 32'sh000027cf;
	assign w_sys_tmp714 = (w_sys_tmp715 + r_run_k_17);
	assign w_sys_tmp715 = 32'sh00002850;
	assign w_sys_tmp720 = (w_sys_tmp721 + r_run_k_17);
	assign w_sys_tmp721 = 32'sh000028d1;
	assign w_sys_tmp726 = (w_sys_tmp727 + r_run_k_17);
	assign w_sys_tmp727 = 32'sh00002952;
	assign w_sys_tmp732 = (w_sys_tmp733 + r_run_k_17);
	assign w_sys_tmp733 = 32'sh000029d3;
	assign w_sys_tmp738 = (w_sys_tmp739 + r_run_k_17);
	assign w_sys_tmp739 = 32'sh00002a54;
	assign w_sys_tmp744 = (w_sys_tmp745 + r_run_k_17);
	assign w_sys_tmp745 = 32'sh00002ad5;
	assign w_sys_tmp750 = (w_sys_tmp751 + r_run_k_17);
	assign w_sys_tmp751 = 32'sh00002b56;
	assign w_sys_tmp756 = (w_sys_tmp757 + r_run_k_17);
	assign w_sys_tmp757 = 32'sh00002bd7;
	assign w_sys_tmp762 = (w_sys_tmp763 + r_run_k_17);
	assign w_sys_tmp763 = 32'sh00002c58;
	assign w_sys_tmp768 = (w_sys_tmp769 + r_run_k_17);
	assign w_sys_tmp769 = 32'sh00002cd9;
	assign w_sys_tmp774 = (w_sys_tmp775 + r_run_k_17);
	assign w_sys_tmp775 = 32'sh00002d5a;
	assign w_sys_tmp780 = (w_sys_tmp781 + r_run_k_17);
	assign w_sys_tmp781 = 32'sh00002ddb;
	assign w_sys_tmp786 = (w_sys_tmp787 + r_run_k_17);
	assign w_sys_tmp787 = 32'sh00002e5c;
	assign w_sys_tmp792 = (w_sys_tmp793 + r_run_k_17);
	assign w_sys_tmp793 = 32'sh00002edd;
	assign w_sys_tmp798 = (w_sys_tmp799 + r_run_k_17);
	assign w_sys_tmp799 = 32'sh00002f5e;
	assign w_sys_tmp804 = (w_sys_tmp805 + r_run_k_17);
	assign w_sys_tmp805 = 32'sh00002fdf;
	assign w_sys_tmp810 = (w_sys_tmp811 + r_run_k_17);
	assign w_sys_tmp811 = 32'sh00003060;
	assign w_sys_tmp816 = (w_sys_tmp817 + r_run_k_17);
	assign w_sys_tmp817 = 32'sh000030e1;
	assign w_sys_tmp834 = (w_sys_tmp835 + r_run_k_17);
	assign w_sys_tmp835 = 32'sh00003162;
	assign w_sys_tmp840 = (w_sys_tmp841 + r_run_k_17);
	assign w_sys_tmp841 = 32'sh000031e3;
	assign w_sys_tmp846 = (w_sys_tmp847 + r_run_k_17);
	assign w_sys_tmp847 = 32'sh00003264;
	assign w_sys_tmp852 = (w_sys_tmp853 + r_run_k_17);
	assign w_sys_tmp853 = 32'sh000032e5;
	assign w_sys_tmp858 = (w_sys_tmp859 + r_run_k_17);
	assign w_sys_tmp859 = 32'sh00003366;
	assign w_sys_tmp864 = (w_sys_tmp865 + r_run_k_17);
	assign w_sys_tmp865 = 32'sh000033e7;
	assign w_sys_tmp870 = (w_sys_tmp871 + r_run_k_17);
	assign w_sys_tmp871 = 32'sh00003468;
	assign w_sys_tmp876 = (w_sys_tmp877 + r_run_k_17);
	assign w_sys_tmp877 = 32'sh000034e9;
	assign w_sys_tmp882 = (w_sys_tmp883 + r_run_k_17);
	assign w_sys_tmp883 = 32'sh0000356a;
	assign w_sys_tmp888 = (w_sys_tmp889 + r_run_k_17);
	assign w_sys_tmp889 = 32'sh000035eb;
	assign w_sys_tmp894 = (w_sys_tmp895 + r_run_k_17);
	assign w_sys_tmp895 = 32'sh0000366c;
	assign w_sys_tmp900 = (w_sys_tmp901 + r_run_k_17);
	assign w_sys_tmp901 = 32'sh000036ed;
	assign w_sys_tmp906 = (w_sys_tmp907 + r_run_k_17);
	assign w_sys_tmp907 = 32'sh0000376e;
	assign w_sys_tmp912 = (w_sys_tmp913 + r_run_k_17);
	assign w_sys_tmp913 = 32'sh000037ef;
	assign w_sys_tmp918 = (w_sys_tmp919 + r_run_k_17);
	assign w_sys_tmp919 = 32'sh00003870;
	assign w_sys_tmp924 = (w_sys_tmp925 + r_run_k_17);
	assign w_sys_tmp925 = 32'sh000038f1;
	assign w_sys_tmp930 = (w_sys_tmp931 + r_run_k_17);
	assign w_sys_tmp931 = 32'sh00003972;
	assign w_sys_tmp936 = (w_sys_tmp937 + r_run_k_17);
	assign w_sys_tmp937 = 32'sh000039f3;
	assign w_sys_tmp942 = (w_sys_tmp943 + r_run_k_17);
	assign w_sys_tmp943 = 32'sh00003a74;
	assign w_sys_tmp948 = (w_sys_tmp949 + r_run_k_17);
	assign w_sys_tmp949 = 32'sh00003af5;
	assign w_sys_tmp954 = (w_sys_tmp955 + r_run_k_17);
	assign w_sys_tmp955 = 32'sh00003b76;
	assign w_sys_tmp960 = (w_sys_tmp961 + r_run_k_17);
	assign w_sys_tmp961 = 32'sh00003bf7;
	assign w_sys_tmp966 = (w_sys_tmp967 + r_run_k_17);
	assign w_sys_tmp967 = 32'sh00003c78;
	assign w_sys_tmp972 = (w_sys_tmp973 + r_run_k_17);
	assign w_sys_tmp973 = 32'sh00003cf9;
	assign w_sys_tmp978 = (w_sys_tmp979 + r_run_k_17);
	assign w_sys_tmp979 = 32'sh00003d7a;
	assign w_sys_tmp984 = (w_sys_tmp985 + r_run_k_17);
	assign w_sys_tmp985 = 32'sh00003dfb;
	assign w_sys_tmp990 = (w_sys_tmp991 + r_run_k_17);
	assign w_sys_tmp991 = 32'sh00003e7c;
	assign w_sys_tmp996 = (w_sys_tmp997 + r_run_k_17);
	assign w_sys_tmp997 = 32'sh00003efd;
	assign w_sys_tmp1002 = (w_sys_tmp1003 + r_run_k_17);
	assign w_sys_tmp1003 = 32'sh00003f7e;
	assign w_sys_tmp1008 = (w_sys_tmp1009 + r_run_k_17);
	assign w_sys_tmp1009 = 32'sh00003fff;
	assign w_sys_tmp1014 = (w_sys_tmp1015 + r_run_k_17);
	assign w_sys_tmp1015 = 32'sh00004080;
	assign w_sys_tmp1020 = (w_sys_tmp1021 + r_run_k_17);
	assign w_sys_tmp1021 = 32'sh00004101;
	assign w_sys_tmp1025 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp1026 = 32'sh00000020;
	assign w_sys_tmp1027 = ( !w_sys_tmp1028 );
	assign w_sys_tmp1028 = (w_sys_tmp1029 < r_run_k_17);
	assign w_sys_tmp1029 = 32'sh00000041;
	assign w_sys_tmp1032 = (w_sys_tmp1033 + r_run_k_17);
	assign w_sys_tmp1033 = 32'sh00000081;
	assign w_sys_tmp1034 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1038 = (w_sys_tmp1039 + r_run_k_17);
	assign w_sys_tmp1039 = 32'sh00000102;
	assign w_sys_tmp1044 = (w_sys_tmp1045 + r_run_k_17);
	assign w_sys_tmp1045 = 32'sh00000183;
	assign w_sys_tmp1050 = (w_sys_tmp1051 + r_run_k_17);
	assign w_sys_tmp1051 = 32'sh00000204;
	assign w_sys_tmp1056 = (w_sys_tmp1057 + r_run_k_17);
	assign w_sys_tmp1057 = 32'sh00000285;
	assign w_sys_tmp1062 = (w_sys_tmp1063 + r_run_k_17);
	assign w_sys_tmp1063 = 32'sh00000306;
	assign w_sys_tmp1068 = (w_sys_tmp1069 + r_run_k_17);
	assign w_sys_tmp1069 = 32'sh00000387;
	assign w_sys_tmp1074 = (w_sys_tmp1075 + r_run_k_17);
	assign w_sys_tmp1075 = 32'sh00000408;
	assign w_sys_tmp1080 = (w_sys_tmp1081 + r_run_k_17);
	assign w_sys_tmp1081 = 32'sh00000489;
	assign w_sys_tmp1086 = (w_sys_tmp1087 + r_run_k_17);
	assign w_sys_tmp1087 = 32'sh0000050a;
	assign w_sys_tmp1092 = (w_sys_tmp1093 + r_run_k_17);
	assign w_sys_tmp1093 = 32'sh0000058b;
	assign w_sys_tmp1098 = (w_sys_tmp1099 + r_run_k_17);
	assign w_sys_tmp1099 = 32'sh0000060c;
	assign w_sys_tmp1104 = (w_sys_tmp1105 + r_run_k_17);
	assign w_sys_tmp1105 = 32'sh0000068d;
	assign w_sys_tmp1110 = (w_sys_tmp1111 + r_run_k_17);
	assign w_sys_tmp1111 = 32'sh0000070e;
	assign w_sys_tmp1116 = (w_sys_tmp1117 + r_run_k_17);
	assign w_sys_tmp1117 = 32'sh0000078f;
	assign w_sys_tmp1122 = (w_sys_tmp1123 + r_run_k_17);
	assign w_sys_tmp1123 = 32'sh00000810;
	assign w_sys_tmp1128 = (w_sys_tmp1129 + r_run_k_17);
	assign w_sys_tmp1129 = 32'sh00000891;
	assign w_sys_tmp1134 = (w_sys_tmp1135 + r_run_k_17);
	assign w_sys_tmp1135 = 32'sh00000912;
	assign w_sys_tmp1140 = (w_sys_tmp1141 + r_run_k_17);
	assign w_sys_tmp1141 = 32'sh00000993;
	assign w_sys_tmp1146 = (w_sys_tmp1147 + r_run_k_17);
	assign w_sys_tmp1147 = 32'sh00000a14;
	assign w_sys_tmp1152 = (w_sys_tmp1153 + r_run_k_17);
	assign w_sys_tmp1153 = 32'sh00000a95;
	assign w_sys_tmp1158 = (w_sys_tmp1159 + r_run_k_17);
	assign w_sys_tmp1159 = 32'sh00000b16;
	assign w_sys_tmp1164 = (w_sys_tmp1165 + r_run_k_17);
	assign w_sys_tmp1165 = 32'sh00000b97;
	assign w_sys_tmp1170 = (w_sys_tmp1171 + r_run_k_17);
	assign w_sys_tmp1171 = 32'sh00000c18;
	assign w_sys_tmp1176 = (w_sys_tmp1177 + r_run_k_17);
	assign w_sys_tmp1177 = 32'sh00000c99;
	assign w_sys_tmp1182 = (w_sys_tmp1183 + r_run_k_17);
	assign w_sys_tmp1183 = 32'sh00000d1a;
	assign w_sys_tmp1188 = (w_sys_tmp1189 + r_run_k_17);
	assign w_sys_tmp1189 = 32'sh00000d9b;
	assign w_sys_tmp1194 = (w_sys_tmp1195 + r_run_k_17);
	assign w_sys_tmp1195 = 32'sh00000e1c;
	assign w_sys_tmp1200 = (w_sys_tmp1201 + r_run_k_17);
	assign w_sys_tmp1201 = 32'sh00000e9d;
	assign w_sys_tmp1206 = (w_sys_tmp1207 + r_run_k_17);
	assign w_sys_tmp1207 = 32'sh00000f1e;
	assign w_sys_tmp1212 = (w_sys_tmp1213 + r_run_k_17);
	assign w_sys_tmp1213 = 32'sh00000f9f;
	assign w_sys_tmp1218 = (w_sys_tmp1219 + r_run_k_17);
	assign w_sys_tmp1219 = 32'sh00001020;
	assign w_sys_tmp1224 = (w_sys_tmp1225 + r_run_k_17);
	assign w_sys_tmp1225 = 32'sh000010a1;
	assign w_sys_tmp1242 = (w_sys_tmp1243 + r_run_k_17);
	assign w_sys_tmp1243 = 32'sh00001122;
	assign w_sys_tmp1248 = (w_sys_tmp1249 + r_run_k_17);
	assign w_sys_tmp1249 = 32'sh000011a3;
	assign w_sys_tmp1254 = (w_sys_tmp1255 + r_run_k_17);
	assign w_sys_tmp1255 = 32'sh00001224;
	assign w_sys_tmp1260 = (w_sys_tmp1261 + r_run_k_17);
	assign w_sys_tmp1261 = 32'sh000012a5;
	assign w_sys_tmp1266 = (w_sys_tmp1267 + r_run_k_17);
	assign w_sys_tmp1267 = 32'sh00001326;
	assign w_sys_tmp1272 = (w_sys_tmp1273 + r_run_k_17);
	assign w_sys_tmp1273 = 32'sh000013a7;
	assign w_sys_tmp1278 = (w_sys_tmp1279 + r_run_k_17);
	assign w_sys_tmp1279 = 32'sh00001428;
	assign w_sys_tmp1284 = (w_sys_tmp1285 + r_run_k_17);
	assign w_sys_tmp1285 = 32'sh000014a9;
	assign w_sys_tmp1290 = (w_sys_tmp1291 + r_run_k_17);
	assign w_sys_tmp1291 = 32'sh0000152a;
	assign w_sys_tmp1296 = (w_sys_tmp1297 + r_run_k_17);
	assign w_sys_tmp1297 = 32'sh000015ab;
	assign w_sys_tmp1302 = (w_sys_tmp1303 + r_run_k_17);
	assign w_sys_tmp1303 = 32'sh0000162c;
	assign w_sys_tmp1308 = (w_sys_tmp1309 + r_run_k_17);
	assign w_sys_tmp1309 = 32'sh000016ad;
	assign w_sys_tmp1314 = (w_sys_tmp1315 + r_run_k_17);
	assign w_sys_tmp1315 = 32'sh0000172e;
	assign w_sys_tmp1320 = (w_sys_tmp1321 + r_run_k_17);
	assign w_sys_tmp1321 = 32'sh000017af;
	assign w_sys_tmp1326 = (w_sys_tmp1327 + r_run_k_17);
	assign w_sys_tmp1327 = 32'sh00001830;
	assign w_sys_tmp1332 = (w_sys_tmp1333 + r_run_k_17);
	assign w_sys_tmp1333 = 32'sh000018b1;
	assign w_sys_tmp1338 = (w_sys_tmp1339 + r_run_k_17);
	assign w_sys_tmp1339 = 32'sh00001932;
	assign w_sys_tmp1344 = (w_sys_tmp1345 + r_run_k_17);
	assign w_sys_tmp1345 = 32'sh000019b3;
	assign w_sys_tmp1350 = (w_sys_tmp1351 + r_run_k_17);
	assign w_sys_tmp1351 = 32'sh00001a34;
	assign w_sys_tmp1356 = (w_sys_tmp1357 + r_run_k_17);
	assign w_sys_tmp1357 = 32'sh00001ab5;
	assign w_sys_tmp1362 = (w_sys_tmp1363 + r_run_k_17);
	assign w_sys_tmp1363 = 32'sh00001b36;
	assign w_sys_tmp1368 = (w_sys_tmp1369 + r_run_k_17);
	assign w_sys_tmp1369 = 32'sh00001bb7;
	assign w_sys_tmp1374 = (w_sys_tmp1375 + r_run_k_17);
	assign w_sys_tmp1375 = 32'sh00001c38;
	assign w_sys_tmp1380 = (w_sys_tmp1381 + r_run_k_17);
	assign w_sys_tmp1381 = 32'sh00001cb9;
	assign w_sys_tmp1386 = (w_sys_tmp1387 + r_run_k_17);
	assign w_sys_tmp1387 = 32'sh00001d3a;
	assign w_sys_tmp1392 = (w_sys_tmp1393 + r_run_k_17);
	assign w_sys_tmp1393 = 32'sh00001dbb;
	assign w_sys_tmp1398 = (w_sys_tmp1399 + r_run_k_17);
	assign w_sys_tmp1399 = 32'sh00001e3c;
	assign w_sys_tmp1404 = (w_sys_tmp1405 + r_run_k_17);
	assign w_sys_tmp1405 = 32'sh00001ebd;
	assign w_sys_tmp1410 = (w_sys_tmp1411 + r_run_k_17);
	assign w_sys_tmp1411 = 32'sh00001f3e;
	assign w_sys_tmp1416 = (w_sys_tmp1417 + r_run_k_17);
	assign w_sys_tmp1417 = 32'sh00001fbf;
	assign w_sys_tmp1422 = (w_sys_tmp1423 + r_run_k_17);
	assign w_sys_tmp1423 = 32'sh00002040;
	assign w_sys_tmp1428 = (w_sys_tmp1429 + r_run_k_17);
	assign w_sys_tmp1429 = 32'sh000020c1;
	assign w_sys_tmp1446 = (w_sys_tmp1447 + r_run_k_17);
	assign w_sys_tmp1447 = 32'sh00002142;
	assign w_sys_tmp1452 = (w_sys_tmp1453 + r_run_k_17);
	assign w_sys_tmp1453 = 32'sh000021c3;
	assign w_sys_tmp1458 = (w_sys_tmp1459 + r_run_k_17);
	assign w_sys_tmp1459 = 32'sh00002244;
	assign w_sys_tmp1464 = (w_sys_tmp1465 + r_run_k_17);
	assign w_sys_tmp1465 = 32'sh000022c5;
	assign w_sys_tmp1470 = (w_sys_tmp1471 + r_run_k_17);
	assign w_sys_tmp1471 = 32'sh00002346;
	assign w_sys_tmp1476 = (w_sys_tmp1477 + r_run_k_17);
	assign w_sys_tmp1477 = 32'sh000023c7;
	assign w_sys_tmp1482 = (w_sys_tmp1483 + r_run_k_17);
	assign w_sys_tmp1483 = 32'sh00002448;
	assign w_sys_tmp1488 = (w_sys_tmp1489 + r_run_k_17);
	assign w_sys_tmp1489 = 32'sh000024c9;
	assign w_sys_tmp1494 = (w_sys_tmp1495 + r_run_k_17);
	assign w_sys_tmp1495 = 32'sh0000254a;
	assign w_sys_tmp1500 = (w_sys_tmp1501 + r_run_k_17);
	assign w_sys_tmp1501 = 32'sh000025cb;
	assign w_sys_tmp1506 = (w_sys_tmp1507 + r_run_k_17);
	assign w_sys_tmp1507 = 32'sh0000264c;
	assign w_sys_tmp1512 = (w_sys_tmp1513 + r_run_k_17);
	assign w_sys_tmp1513 = 32'sh000026cd;
	assign w_sys_tmp1518 = (w_sys_tmp1519 + r_run_k_17);
	assign w_sys_tmp1519 = 32'sh0000274e;
	assign w_sys_tmp1524 = (w_sys_tmp1525 + r_run_k_17);
	assign w_sys_tmp1525 = 32'sh000027cf;
	assign w_sys_tmp1530 = (w_sys_tmp1531 + r_run_k_17);
	assign w_sys_tmp1531 = 32'sh00002850;
	assign w_sys_tmp1536 = (w_sys_tmp1537 + r_run_k_17);
	assign w_sys_tmp1537 = 32'sh000028d1;
	assign w_sys_tmp1542 = (w_sys_tmp1543 + r_run_k_17);
	assign w_sys_tmp1543 = 32'sh00002952;
	assign w_sys_tmp1548 = (w_sys_tmp1549 + r_run_k_17);
	assign w_sys_tmp1549 = 32'sh000029d3;
	assign w_sys_tmp1554 = (w_sys_tmp1555 + r_run_k_17);
	assign w_sys_tmp1555 = 32'sh00002a54;
	assign w_sys_tmp1560 = (w_sys_tmp1561 + r_run_k_17);
	assign w_sys_tmp1561 = 32'sh00002ad5;
	assign w_sys_tmp1566 = (w_sys_tmp1567 + r_run_k_17);
	assign w_sys_tmp1567 = 32'sh00002b56;
	assign w_sys_tmp1572 = (w_sys_tmp1573 + r_run_k_17);
	assign w_sys_tmp1573 = 32'sh00002bd7;
	assign w_sys_tmp1578 = (w_sys_tmp1579 + r_run_k_17);
	assign w_sys_tmp1579 = 32'sh00002c58;
	assign w_sys_tmp1584 = (w_sys_tmp1585 + r_run_k_17);
	assign w_sys_tmp1585 = 32'sh00002cd9;
	assign w_sys_tmp1590 = (w_sys_tmp1591 + r_run_k_17);
	assign w_sys_tmp1591 = 32'sh00002d5a;
	assign w_sys_tmp1596 = (w_sys_tmp1597 + r_run_k_17);
	assign w_sys_tmp1597 = 32'sh00002ddb;
	assign w_sys_tmp1602 = (w_sys_tmp1603 + r_run_k_17);
	assign w_sys_tmp1603 = 32'sh00002e5c;
	assign w_sys_tmp1608 = (w_sys_tmp1609 + r_run_k_17);
	assign w_sys_tmp1609 = 32'sh00002edd;
	assign w_sys_tmp1614 = (w_sys_tmp1615 + r_run_k_17);
	assign w_sys_tmp1615 = 32'sh00002f5e;
	assign w_sys_tmp1620 = (w_sys_tmp1621 + r_run_k_17);
	assign w_sys_tmp1621 = 32'sh00002fdf;
	assign w_sys_tmp1626 = (w_sys_tmp1627 + r_run_k_17);
	assign w_sys_tmp1627 = 32'sh00003060;
	assign w_sys_tmp1632 = (w_sys_tmp1633 + r_run_k_17);
	assign w_sys_tmp1633 = 32'sh000030e1;
	assign w_sys_tmp1650 = (w_sys_tmp1651 + r_run_k_17);
	assign w_sys_tmp1651 = 32'sh00003162;
	assign w_sys_tmp1656 = (w_sys_tmp1657 + r_run_k_17);
	assign w_sys_tmp1657 = 32'sh000031e3;
	assign w_sys_tmp1662 = (w_sys_tmp1663 + r_run_k_17);
	assign w_sys_tmp1663 = 32'sh00003264;
	assign w_sys_tmp1668 = (w_sys_tmp1669 + r_run_k_17);
	assign w_sys_tmp1669 = 32'sh000032e5;
	assign w_sys_tmp1674 = (w_sys_tmp1675 + r_run_k_17);
	assign w_sys_tmp1675 = 32'sh00003366;
	assign w_sys_tmp1680 = (w_sys_tmp1681 + r_run_k_17);
	assign w_sys_tmp1681 = 32'sh000033e7;
	assign w_sys_tmp1686 = (w_sys_tmp1687 + r_run_k_17);
	assign w_sys_tmp1687 = 32'sh00003468;
	assign w_sys_tmp1692 = (w_sys_tmp1693 + r_run_k_17);
	assign w_sys_tmp1693 = 32'sh000034e9;
	assign w_sys_tmp1698 = (w_sys_tmp1699 + r_run_k_17);
	assign w_sys_tmp1699 = 32'sh0000356a;
	assign w_sys_tmp1704 = (w_sys_tmp1705 + r_run_k_17);
	assign w_sys_tmp1705 = 32'sh000035eb;
	assign w_sys_tmp1710 = (w_sys_tmp1711 + r_run_k_17);
	assign w_sys_tmp1711 = 32'sh0000366c;
	assign w_sys_tmp1716 = (w_sys_tmp1717 + r_run_k_17);
	assign w_sys_tmp1717 = 32'sh000036ed;
	assign w_sys_tmp1722 = (w_sys_tmp1723 + r_run_k_17);
	assign w_sys_tmp1723 = 32'sh0000376e;
	assign w_sys_tmp1728 = (w_sys_tmp1729 + r_run_k_17);
	assign w_sys_tmp1729 = 32'sh000037ef;
	assign w_sys_tmp1734 = (w_sys_tmp1735 + r_run_k_17);
	assign w_sys_tmp1735 = 32'sh00003870;
	assign w_sys_tmp1740 = (w_sys_tmp1741 + r_run_k_17);
	assign w_sys_tmp1741 = 32'sh000038f1;
	assign w_sys_tmp1746 = (w_sys_tmp1747 + r_run_k_17);
	assign w_sys_tmp1747 = 32'sh00003972;
	assign w_sys_tmp1752 = (w_sys_tmp1753 + r_run_k_17);
	assign w_sys_tmp1753 = 32'sh000039f3;
	assign w_sys_tmp1758 = (w_sys_tmp1759 + r_run_k_17);
	assign w_sys_tmp1759 = 32'sh00003a74;
	assign w_sys_tmp1764 = (w_sys_tmp1765 + r_run_k_17);
	assign w_sys_tmp1765 = 32'sh00003af5;
	assign w_sys_tmp1770 = (w_sys_tmp1771 + r_run_k_17);
	assign w_sys_tmp1771 = 32'sh00003b76;
	assign w_sys_tmp1776 = (w_sys_tmp1777 + r_run_k_17);
	assign w_sys_tmp1777 = 32'sh00003bf7;
	assign w_sys_tmp1782 = (w_sys_tmp1783 + r_run_k_17);
	assign w_sys_tmp1783 = 32'sh00003c78;
	assign w_sys_tmp1788 = (w_sys_tmp1789 + r_run_k_17);
	assign w_sys_tmp1789 = 32'sh00003cf9;
	assign w_sys_tmp1794 = (w_sys_tmp1795 + r_run_k_17);
	assign w_sys_tmp1795 = 32'sh00003d7a;
	assign w_sys_tmp1800 = (w_sys_tmp1801 + r_run_k_17);
	assign w_sys_tmp1801 = 32'sh00003dfb;
	assign w_sys_tmp1806 = (w_sys_tmp1807 + r_run_k_17);
	assign w_sys_tmp1807 = 32'sh00003e7c;
	assign w_sys_tmp1812 = (w_sys_tmp1813 + r_run_k_17);
	assign w_sys_tmp1813 = 32'sh00003efd;
	assign w_sys_tmp1818 = (w_sys_tmp1819 + r_run_k_17);
	assign w_sys_tmp1819 = 32'sh00003f7e;
	assign w_sys_tmp1824 = (w_sys_tmp1825 + r_run_k_17);
	assign w_sys_tmp1825 = 32'sh00003fff;
	assign w_sys_tmp1830 = (w_sys_tmp1831 + r_run_k_17);
	assign w_sys_tmp1831 = 32'sh00004080;
	assign w_sys_tmp1836 = (w_sys_tmp1837 + r_run_k_17);
	assign w_sys_tmp1837 = 32'sh00004101;
	assign w_sys_tmp1842 = (w_sys_tmp1843 + r_run_k_17);
	assign w_sys_tmp1843 = 32'sh000000a1;
	assign w_sys_tmp1848 = (w_sys_tmp1849 + r_run_k_17);
	assign w_sys_tmp1849 = 32'sh00000122;
	assign w_sys_tmp1854 = (w_sys_tmp1855 + r_run_k_17);
	assign w_sys_tmp1855 = 32'sh000001a3;
	assign w_sys_tmp1860 = (w_sys_tmp1861 + r_run_k_17);
	assign w_sys_tmp1861 = 32'sh00000224;
	assign w_sys_tmp1866 = (w_sys_tmp1867 + r_run_k_17);
	assign w_sys_tmp1867 = 32'sh000002a5;
	assign w_sys_tmp1872 = (w_sys_tmp1873 + r_run_k_17);
	assign w_sys_tmp1873 = 32'sh00000326;
	assign w_sys_tmp1878 = (w_sys_tmp1879 + r_run_k_17);
	assign w_sys_tmp1879 = 32'sh000003a7;
	assign w_sys_tmp1884 = (w_sys_tmp1885 + r_run_k_17);
	assign w_sys_tmp1885 = 32'sh00000428;
	assign w_sys_tmp1890 = (w_sys_tmp1891 + r_run_k_17);
	assign w_sys_tmp1891 = 32'sh000004a9;
	assign w_sys_tmp1896 = (w_sys_tmp1897 + r_run_k_17);
	assign w_sys_tmp1897 = 32'sh0000052a;
	assign w_sys_tmp1902 = (w_sys_tmp1903 + r_run_k_17);
	assign w_sys_tmp1903 = 32'sh000005ab;
	assign w_sys_tmp1908 = (w_sys_tmp1909 + r_run_k_17);
	assign w_sys_tmp1909 = 32'sh0000062c;
	assign w_sys_tmp1914 = (w_sys_tmp1915 + r_run_k_17);
	assign w_sys_tmp1915 = 32'sh000006ad;
	assign w_sys_tmp1920 = (w_sys_tmp1921 + r_run_k_17);
	assign w_sys_tmp1921 = 32'sh0000072e;
	assign w_sys_tmp1926 = (w_sys_tmp1927 + r_run_k_17);
	assign w_sys_tmp1927 = 32'sh000007af;
	assign w_sys_tmp1932 = (w_sys_tmp1933 + r_run_k_17);
	assign w_sys_tmp1933 = 32'sh00000830;
	assign w_sys_tmp1938 = (w_sys_tmp1939 + r_run_k_17);
	assign w_sys_tmp1939 = 32'sh000008b1;
	assign w_sys_tmp1944 = (w_sys_tmp1945 + r_run_k_17);
	assign w_sys_tmp1945 = 32'sh00000932;
	assign w_sys_tmp1950 = (w_sys_tmp1951 + r_run_k_17);
	assign w_sys_tmp1951 = 32'sh000009b3;
	assign w_sys_tmp1956 = (w_sys_tmp1957 + r_run_k_17);
	assign w_sys_tmp1957 = 32'sh00000a34;
	assign w_sys_tmp1962 = (w_sys_tmp1963 + r_run_k_17);
	assign w_sys_tmp1963 = 32'sh00000ab5;
	assign w_sys_tmp1968 = (w_sys_tmp1969 + r_run_k_17);
	assign w_sys_tmp1969 = 32'sh00000b36;
	assign w_sys_tmp1974 = (w_sys_tmp1975 + r_run_k_17);
	assign w_sys_tmp1975 = 32'sh00000bb7;
	assign w_sys_tmp1980 = (w_sys_tmp1981 + r_run_k_17);
	assign w_sys_tmp1981 = 32'sh00000c38;
	assign w_sys_tmp1986 = (w_sys_tmp1987 + r_run_k_17);
	assign w_sys_tmp1987 = 32'sh00000cb9;
	assign w_sys_tmp1992 = (w_sys_tmp1993 + r_run_k_17);
	assign w_sys_tmp1993 = 32'sh00000d3a;
	assign w_sys_tmp1998 = (w_sys_tmp1999 + r_run_k_17);
	assign w_sys_tmp1999 = 32'sh00000dbb;
	assign w_sys_tmp2004 = (w_sys_tmp2005 + r_run_k_17);
	assign w_sys_tmp2005 = 32'sh00000e3c;
	assign w_sys_tmp2010 = (w_sys_tmp2011 + r_run_k_17);
	assign w_sys_tmp2011 = 32'sh00000ebd;
	assign w_sys_tmp2016 = (w_sys_tmp2017 + r_run_k_17);
	assign w_sys_tmp2017 = 32'sh00000f3e;
	assign w_sys_tmp2022 = (w_sys_tmp2023 + r_run_k_17);
	assign w_sys_tmp2023 = 32'sh00000fbf;
	assign w_sys_tmp2028 = (w_sys_tmp2029 + r_run_k_17);
	assign w_sys_tmp2029 = 32'sh00001040;
	assign w_sys_tmp2034 = (w_sys_tmp2035 + r_run_k_17);
	assign w_sys_tmp2035 = 32'sh000010c1;
	assign w_sys_tmp2052 = (w_sys_tmp2053 + r_run_k_17);
	assign w_sys_tmp2053 = 32'sh00001142;
	assign w_sys_tmp2058 = (w_sys_tmp2059 + r_run_k_17);
	assign w_sys_tmp2059 = 32'sh000011c3;
	assign w_sys_tmp2064 = (w_sys_tmp2065 + r_run_k_17);
	assign w_sys_tmp2065 = 32'sh00001244;
	assign w_sys_tmp2070 = (w_sys_tmp2071 + r_run_k_17);
	assign w_sys_tmp2071 = 32'sh000012c5;
	assign w_sys_tmp2076 = (w_sys_tmp2077 + r_run_k_17);
	assign w_sys_tmp2077 = 32'sh00001346;
	assign w_sys_tmp2082 = (w_sys_tmp2083 + r_run_k_17);
	assign w_sys_tmp2083 = 32'sh000013c7;
	assign w_sys_tmp2088 = (w_sys_tmp2089 + r_run_k_17);
	assign w_sys_tmp2089 = 32'sh00001448;
	assign w_sys_tmp2094 = (w_sys_tmp2095 + r_run_k_17);
	assign w_sys_tmp2095 = 32'sh000014c9;
	assign w_sys_tmp2100 = (w_sys_tmp2101 + r_run_k_17);
	assign w_sys_tmp2101 = 32'sh0000154a;
	assign w_sys_tmp2106 = (w_sys_tmp2107 + r_run_k_17);
	assign w_sys_tmp2107 = 32'sh000015cb;
	assign w_sys_tmp2112 = (w_sys_tmp2113 + r_run_k_17);
	assign w_sys_tmp2113 = 32'sh0000164c;
	assign w_sys_tmp2118 = (w_sys_tmp2119 + r_run_k_17);
	assign w_sys_tmp2119 = 32'sh000016cd;
	assign w_sys_tmp2124 = (w_sys_tmp2125 + r_run_k_17);
	assign w_sys_tmp2125 = 32'sh0000174e;
	assign w_sys_tmp2130 = (w_sys_tmp2131 + r_run_k_17);
	assign w_sys_tmp2131 = 32'sh000017cf;
	assign w_sys_tmp2136 = (w_sys_tmp2137 + r_run_k_17);
	assign w_sys_tmp2137 = 32'sh00001850;
	assign w_sys_tmp2142 = (w_sys_tmp2143 + r_run_k_17);
	assign w_sys_tmp2143 = 32'sh000018d1;
	assign w_sys_tmp2148 = (w_sys_tmp2149 + r_run_k_17);
	assign w_sys_tmp2149 = 32'sh00001952;
	assign w_sys_tmp2154 = (w_sys_tmp2155 + r_run_k_17);
	assign w_sys_tmp2155 = 32'sh000019d3;
	assign w_sys_tmp2160 = (w_sys_tmp2161 + r_run_k_17);
	assign w_sys_tmp2161 = 32'sh00001a54;
	assign w_sys_tmp2166 = (w_sys_tmp2167 + r_run_k_17);
	assign w_sys_tmp2167 = 32'sh00001ad5;
	assign w_sys_tmp2172 = (w_sys_tmp2173 + r_run_k_17);
	assign w_sys_tmp2173 = 32'sh00001b56;
	assign w_sys_tmp2178 = (w_sys_tmp2179 + r_run_k_17);
	assign w_sys_tmp2179 = 32'sh00001bd7;
	assign w_sys_tmp2184 = (w_sys_tmp2185 + r_run_k_17);
	assign w_sys_tmp2185 = 32'sh00001c58;
	assign w_sys_tmp2190 = (w_sys_tmp2191 + r_run_k_17);
	assign w_sys_tmp2191 = 32'sh00001cd9;
	assign w_sys_tmp2196 = (w_sys_tmp2197 + r_run_k_17);
	assign w_sys_tmp2197 = 32'sh00001d5a;
	assign w_sys_tmp2202 = (w_sys_tmp2203 + r_run_k_17);
	assign w_sys_tmp2203 = 32'sh00001ddb;
	assign w_sys_tmp2208 = (w_sys_tmp2209 + r_run_k_17);
	assign w_sys_tmp2209 = 32'sh00001e5c;
	assign w_sys_tmp2214 = (w_sys_tmp2215 + r_run_k_17);
	assign w_sys_tmp2215 = 32'sh00001edd;
	assign w_sys_tmp2220 = (w_sys_tmp2221 + r_run_k_17);
	assign w_sys_tmp2221 = 32'sh00001f5e;
	assign w_sys_tmp2226 = (w_sys_tmp2227 + r_run_k_17);
	assign w_sys_tmp2227 = 32'sh00001fdf;
	assign w_sys_tmp2232 = (w_sys_tmp2233 + r_run_k_17);
	assign w_sys_tmp2233 = 32'sh00002060;
	assign w_sys_tmp2238 = (w_sys_tmp2239 + r_run_k_17);
	assign w_sys_tmp2239 = 32'sh000020e1;
	assign w_sys_tmp2256 = (w_sys_tmp2257 + r_run_k_17);
	assign w_sys_tmp2257 = 32'sh00002162;
	assign w_sys_tmp2262 = (w_sys_tmp2263 + r_run_k_17);
	assign w_sys_tmp2263 = 32'sh000021e3;
	assign w_sys_tmp2268 = (w_sys_tmp2269 + r_run_k_17);
	assign w_sys_tmp2269 = 32'sh00002264;
	assign w_sys_tmp2274 = (w_sys_tmp2275 + r_run_k_17);
	assign w_sys_tmp2275 = 32'sh000022e5;
	assign w_sys_tmp2280 = (w_sys_tmp2281 + r_run_k_17);
	assign w_sys_tmp2281 = 32'sh00002366;
	assign w_sys_tmp2286 = (w_sys_tmp2287 + r_run_k_17);
	assign w_sys_tmp2287 = 32'sh000023e7;
	assign w_sys_tmp2292 = (w_sys_tmp2293 + r_run_k_17);
	assign w_sys_tmp2293 = 32'sh00002468;
	assign w_sys_tmp2298 = (w_sys_tmp2299 + r_run_k_17);
	assign w_sys_tmp2299 = 32'sh000024e9;
	assign w_sys_tmp2304 = (w_sys_tmp2305 + r_run_k_17);
	assign w_sys_tmp2305 = 32'sh0000256a;
	assign w_sys_tmp2310 = (w_sys_tmp2311 + r_run_k_17);
	assign w_sys_tmp2311 = 32'sh000025eb;
	assign w_sys_tmp2316 = (w_sys_tmp2317 + r_run_k_17);
	assign w_sys_tmp2317 = 32'sh0000266c;
	assign w_sys_tmp2322 = (w_sys_tmp2323 + r_run_k_17);
	assign w_sys_tmp2323 = 32'sh000026ed;
	assign w_sys_tmp2328 = (w_sys_tmp2329 + r_run_k_17);
	assign w_sys_tmp2329 = 32'sh0000276e;
	assign w_sys_tmp2334 = (w_sys_tmp2335 + r_run_k_17);
	assign w_sys_tmp2335 = 32'sh000027ef;
	assign w_sys_tmp2340 = (w_sys_tmp2341 + r_run_k_17);
	assign w_sys_tmp2341 = 32'sh00002870;
	assign w_sys_tmp2346 = (w_sys_tmp2347 + r_run_k_17);
	assign w_sys_tmp2347 = 32'sh000028f1;
	assign w_sys_tmp2352 = (w_sys_tmp2353 + r_run_k_17);
	assign w_sys_tmp2353 = 32'sh00002972;
	assign w_sys_tmp2358 = (w_sys_tmp2359 + r_run_k_17);
	assign w_sys_tmp2359 = 32'sh000029f3;
	assign w_sys_tmp2364 = (w_sys_tmp2365 + r_run_k_17);
	assign w_sys_tmp2365 = 32'sh00002a74;
	assign w_sys_tmp2370 = (w_sys_tmp2371 + r_run_k_17);
	assign w_sys_tmp2371 = 32'sh00002af5;
	assign w_sys_tmp2376 = (w_sys_tmp2377 + r_run_k_17);
	assign w_sys_tmp2377 = 32'sh00002b76;
	assign w_sys_tmp2382 = (w_sys_tmp2383 + r_run_k_17);
	assign w_sys_tmp2383 = 32'sh00002bf7;
	assign w_sys_tmp2388 = (w_sys_tmp2389 + r_run_k_17);
	assign w_sys_tmp2389 = 32'sh00002c78;
	assign w_sys_tmp2394 = (w_sys_tmp2395 + r_run_k_17);
	assign w_sys_tmp2395 = 32'sh00002cf9;
	assign w_sys_tmp2400 = (w_sys_tmp2401 + r_run_k_17);
	assign w_sys_tmp2401 = 32'sh00002d7a;
	assign w_sys_tmp2406 = (w_sys_tmp2407 + r_run_k_17);
	assign w_sys_tmp2407 = 32'sh00002dfb;
	assign w_sys_tmp2412 = (w_sys_tmp2413 + r_run_k_17);
	assign w_sys_tmp2413 = 32'sh00002e7c;
	assign w_sys_tmp2418 = (w_sys_tmp2419 + r_run_k_17);
	assign w_sys_tmp2419 = 32'sh00002efd;
	assign w_sys_tmp2424 = (w_sys_tmp2425 + r_run_k_17);
	assign w_sys_tmp2425 = 32'sh00002f7e;
	assign w_sys_tmp2430 = (w_sys_tmp2431 + r_run_k_17);
	assign w_sys_tmp2431 = 32'sh00002fff;
	assign w_sys_tmp2436 = (w_sys_tmp2437 + r_run_k_17);
	assign w_sys_tmp2437 = 32'sh00003080;
	assign w_sys_tmp2442 = (w_sys_tmp2443 + r_run_k_17);
	assign w_sys_tmp2443 = 32'sh00003101;
	assign w_sys_tmp2460 = (w_sys_tmp2461 + r_run_k_17);
	assign w_sys_tmp2461 = 32'sh00003182;
	assign w_sys_tmp2466 = (w_sys_tmp2467 + r_run_k_17);
	assign w_sys_tmp2467 = 32'sh00003203;
	assign w_sys_tmp2472 = (w_sys_tmp2473 + r_run_k_17);
	assign w_sys_tmp2473 = 32'sh00003284;
	assign w_sys_tmp2478 = (w_sys_tmp2479 + r_run_k_17);
	assign w_sys_tmp2479 = 32'sh00003305;
	assign w_sys_tmp2484 = (w_sys_tmp2485 + r_run_k_17);
	assign w_sys_tmp2485 = 32'sh00003386;
	assign w_sys_tmp2490 = (w_sys_tmp2491 + r_run_k_17);
	assign w_sys_tmp2491 = 32'sh00003407;
	assign w_sys_tmp2496 = (w_sys_tmp2497 + r_run_k_17);
	assign w_sys_tmp2497 = 32'sh00003488;
	assign w_sys_tmp2502 = (w_sys_tmp2503 + r_run_k_17);
	assign w_sys_tmp2503 = 32'sh00003509;
	assign w_sys_tmp2508 = (w_sys_tmp2509 + r_run_k_17);
	assign w_sys_tmp2509 = 32'sh0000358a;
	assign w_sys_tmp2514 = (w_sys_tmp2515 + r_run_k_17);
	assign w_sys_tmp2515 = 32'sh0000360b;
	assign w_sys_tmp2520 = (w_sys_tmp2521 + r_run_k_17);
	assign w_sys_tmp2521 = 32'sh0000368c;
	assign w_sys_tmp2526 = (w_sys_tmp2527 + r_run_k_17);
	assign w_sys_tmp2527 = 32'sh0000370d;
	assign w_sys_tmp2532 = (w_sys_tmp2533 + r_run_k_17);
	assign w_sys_tmp2533 = 32'sh0000378e;
	assign w_sys_tmp2538 = (w_sys_tmp2539 + r_run_k_17);
	assign w_sys_tmp2539 = 32'sh0000380f;
	assign w_sys_tmp2544 = (w_sys_tmp2545 + r_run_k_17);
	assign w_sys_tmp2545 = 32'sh00003890;
	assign w_sys_tmp2550 = (w_sys_tmp2551 + r_run_k_17);
	assign w_sys_tmp2551 = 32'sh00003911;
	assign w_sys_tmp2556 = (w_sys_tmp2557 + r_run_k_17);
	assign w_sys_tmp2557 = 32'sh00003992;
	assign w_sys_tmp2562 = (w_sys_tmp2563 + r_run_k_17);
	assign w_sys_tmp2563 = 32'sh00003a13;
	assign w_sys_tmp2568 = (w_sys_tmp2569 + r_run_k_17);
	assign w_sys_tmp2569 = 32'sh00003a94;
	assign w_sys_tmp2574 = (w_sys_tmp2575 + r_run_k_17);
	assign w_sys_tmp2575 = 32'sh00003b15;
	assign w_sys_tmp2580 = (w_sys_tmp2581 + r_run_k_17);
	assign w_sys_tmp2581 = 32'sh00003b96;
	assign w_sys_tmp2586 = (w_sys_tmp2587 + r_run_k_17);
	assign w_sys_tmp2587 = 32'sh00003c17;
	assign w_sys_tmp2592 = (w_sys_tmp2593 + r_run_k_17);
	assign w_sys_tmp2593 = 32'sh00003c98;
	assign w_sys_tmp2598 = (w_sys_tmp2599 + r_run_k_17);
	assign w_sys_tmp2599 = 32'sh00003d19;
	assign w_sys_tmp2604 = (w_sys_tmp2605 + r_run_k_17);
	assign w_sys_tmp2605 = 32'sh00003d9a;
	assign w_sys_tmp2610 = (w_sys_tmp2611 + r_run_k_17);
	assign w_sys_tmp2611 = 32'sh00003e1b;
	assign w_sys_tmp2616 = (w_sys_tmp2617 + r_run_k_17);
	assign w_sys_tmp2617 = 32'sh00003e9c;
	assign w_sys_tmp2622 = (w_sys_tmp2623 + r_run_k_17);
	assign w_sys_tmp2623 = 32'sh00003f1d;
	assign w_sys_tmp2628 = (w_sys_tmp2629 + r_run_k_17);
	assign w_sys_tmp2629 = 32'sh00003f9e;
	assign w_sys_tmp2634 = (w_sys_tmp2635 + r_run_k_17);
	assign w_sys_tmp2635 = 32'sh0000401f;
	assign w_sys_tmp2640 = (w_sys_tmp2641 + r_run_k_17);
	assign w_sys_tmp2641 = 32'sh000040a0;
	assign w_sys_tmp2646 = (w_sys_tmp2647 + r_run_k_17);
	assign w_sys_tmp2647 = 32'sh00004121;
	assign w_sys_tmp2652 = (w_sys_tmp2653 + r_run_k_17);
	assign w_sys_tmp2653 = 32'sh000000c1;
	assign w_sys_tmp2658 = (w_sys_tmp2659 + r_run_k_17);
	assign w_sys_tmp2659 = 32'sh00000142;
	assign w_sys_tmp2664 = (w_sys_tmp2665 + r_run_k_17);
	assign w_sys_tmp2665 = 32'sh000001c3;
	assign w_sys_tmp2670 = (w_sys_tmp2671 + r_run_k_17);
	assign w_sys_tmp2671 = 32'sh00000244;
	assign w_sys_tmp2676 = (w_sys_tmp2677 + r_run_k_17);
	assign w_sys_tmp2677 = 32'sh000002c5;
	assign w_sys_tmp2682 = (w_sys_tmp2683 + r_run_k_17);
	assign w_sys_tmp2683 = 32'sh00000346;
	assign w_sys_tmp2688 = (w_sys_tmp2689 + r_run_k_17);
	assign w_sys_tmp2689 = 32'sh000003c7;
	assign w_sys_tmp2694 = (w_sys_tmp2695 + r_run_k_17);
	assign w_sys_tmp2695 = 32'sh00000448;
	assign w_sys_tmp2700 = (w_sys_tmp2701 + r_run_k_17);
	assign w_sys_tmp2701 = 32'sh000004c9;
	assign w_sys_tmp2706 = (w_sys_tmp2707 + r_run_k_17);
	assign w_sys_tmp2707 = 32'sh0000054a;
	assign w_sys_tmp2712 = (w_sys_tmp2713 + r_run_k_17);
	assign w_sys_tmp2713 = 32'sh000005cb;
	assign w_sys_tmp2718 = (w_sys_tmp2719 + r_run_k_17);
	assign w_sys_tmp2719 = 32'sh0000064c;
	assign w_sys_tmp2724 = (w_sys_tmp2725 + r_run_k_17);
	assign w_sys_tmp2725 = 32'sh000006cd;
	assign w_sys_tmp2730 = (w_sys_tmp2731 + r_run_k_17);
	assign w_sys_tmp2731 = 32'sh0000074e;
	assign w_sys_tmp2736 = (w_sys_tmp2737 + r_run_k_17);
	assign w_sys_tmp2737 = 32'sh000007cf;
	assign w_sys_tmp2742 = (w_sys_tmp2743 + r_run_k_17);
	assign w_sys_tmp2743 = 32'sh00000850;
	assign w_sys_tmp2748 = (w_sys_tmp2749 + r_run_k_17);
	assign w_sys_tmp2749 = 32'sh000008d1;
	assign w_sys_tmp2754 = (w_sys_tmp2755 + r_run_k_17);
	assign w_sys_tmp2755 = 32'sh00000952;
	assign w_sys_tmp2760 = (w_sys_tmp2761 + r_run_k_17);
	assign w_sys_tmp2761 = 32'sh000009d3;
	assign w_sys_tmp2766 = (w_sys_tmp2767 + r_run_k_17);
	assign w_sys_tmp2767 = 32'sh00000a54;
	assign w_sys_tmp2772 = (w_sys_tmp2773 + r_run_k_17);
	assign w_sys_tmp2773 = 32'sh00000ad5;
	assign w_sys_tmp2778 = (w_sys_tmp2779 + r_run_k_17);
	assign w_sys_tmp2779 = 32'sh00000b56;
	assign w_sys_tmp2784 = (w_sys_tmp2785 + r_run_k_17);
	assign w_sys_tmp2785 = 32'sh00000bd7;
	assign w_sys_tmp2790 = (w_sys_tmp2791 + r_run_k_17);
	assign w_sys_tmp2791 = 32'sh00000c58;
	assign w_sys_tmp2796 = (w_sys_tmp2797 + r_run_k_17);
	assign w_sys_tmp2797 = 32'sh00000cd9;
	assign w_sys_tmp2802 = (w_sys_tmp2803 + r_run_k_17);
	assign w_sys_tmp2803 = 32'sh00000d5a;
	assign w_sys_tmp2808 = (w_sys_tmp2809 + r_run_k_17);
	assign w_sys_tmp2809 = 32'sh00000ddb;
	assign w_sys_tmp2814 = (w_sys_tmp2815 + r_run_k_17);
	assign w_sys_tmp2815 = 32'sh00000e5c;
	assign w_sys_tmp2820 = (w_sys_tmp2821 + r_run_k_17);
	assign w_sys_tmp2821 = 32'sh00000edd;
	assign w_sys_tmp2826 = (w_sys_tmp2827 + r_run_k_17);
	assign w_sys_tmp2827 = 32'sh00000f5e;
	assign w_sys_tmp2832 = (w_sys_tmp2833 + r_run_k_17);
	assign w_sys_tmp2833 = 32'sh00000fdf;
	assign w_sys_tmp2838 = (w_sys_tmp2839 + r_run_k_17);
	assign w_sys_tmp2839 = 32'sh00001060;
	assign w_sys_tmp2844 = (w_sys_tmp2845 + r_run_k_17);
	assign w_sys_tmp2845 = 32'sh000010e1;
	assign w_sys_tmp2862 = (w_sys_tmp2863 + r_run_k_17);
	assign w_sys_tmp2863 = 32'sh00001162;
	assign w_sys_tmp2868 = (w_sys_tmp2869 + r_run_k_17);
	assign w_sys_tmp2869 = 32'sh000011e3;
	assign w_sys_tmp2874 = (w_sys_tmp2875 + r_run_k_17);
	assign w_sys_tmp2875 = 32'sh00001264;
	assign w_sys_tmp2880 = (w_sys_tmp2881 + r_run_k_17);
	assign w_sys_tmp2881 = 32'sh000012e5;
	assign w_sys_tmp2886 = (w_sys_tmp2887 + r_run_k_17);
	assign w_sys_tmp2887 = 32'sh00001366;
	assign w_sys_tmp2892 = (w_sys_tmp2893 + r_run_k_17);
	assign w_sys_tmp2893 = 32'sh000013e7;
	assign w_sys_tmp2898 = (w_sys_tmp2899 + r_run_k_17);
	assign w_sys_tmp2899 = 32'sh00001468;
	assign w_sys_tmp2904 = (w_sys_tmp2905 + r_run_k_17);
	assign w_sys_tmp2905 = 32'sh000014e9;
	assign w_sys_tmp2910 = (w_sys_tmp2911 + r_run_k_17);
	assign w_sys_tmp2911 = 32'sh0000156a;
	assign w_sys_tmp2916 = (w_sys_tmp2917 + r_run_k_17);
	assign w_sys_tmp2917 = 32'sh000015eb;
	assign w_sys_tmp2922 = (w_sys_tmp2923 + r_run_k_17);
	assign w_sys_tmp2923 = 32'sh0000166c;
	assign w_sys_tmp2928 = (w_sys_tmp2929 + r_run_k_17);
	assign w_sys_tmp2929 = 32'sh000016ed;
	assign w_sys_tmp2934 = (w_sys_tmp2935 + r_run_k_17);
	assign w_sys_tmp2935 = 32'sh0000176e;
	assign w_sys_tmp2940 = (w_sys_tmp2941 + r_run_k_17);
	assign w_sys_tmp2941 = 32'sh000017ef;
	assign w_sys_tmp2946 = (w_sys_tmp2947 + r_run_k_17);
	assign w_sys_tmp2947 = 32'sh00001870;
	assign w_sys_tmp2952 = (w_sys_tmp2953 + r_run_k_17);
	assign w_sys_tmp2953 = 32'sh000018f1;
	assign w_sys_tmp2958 = (w_sys_tmp2959 + r_run_k_17);
	assign w_sys_tmp2959 = 32'sh00001972;
	assign w_sys_tmp2964 = (w_sys_tmp2965 + r_run_k_17);
	assign w_sys_tmp2965 = 32'sh000019f3;
	assign w_sys_tmp2970 = (w_sys_tmp2971 + r_run_k_17);
	assign w_sys_tmp2971 = 32'sh00001a74;
	assign w_sys_tmp2976 = (w_sys_tmp2977 + r_run_k_17);
	assign w_sys_tmp2977 = 32'sh00001af5;
	assign w_sys_tmp2982 = (w_sys_tmp2983 + r_run_k_17);
	assign w_sys_tmp2983 = 32'sh00001b76;
	assign w_sys_tmp2988 = (w_sys_tmp2989 + r_run_k_17);
	assign w_sys_tmp2989 = 32'sh00001bf7;
	assign w_sys_tmp2994 = (w_sys_tmp2995 + r_run_k_17);
	assign w_sys_tmp2995 = 32'sh00001c78;
	assign w_sys_tmp3000 = (w_sys_tmp3001 + r_run_k_17);
	assign w_sys_tmp3001 = 32'sh00001cf9;
	assign w_sys_tmp3006 = (w_sys_tmp3007 + r_run_k_17);
	assign w_sys_tmp3007 = 32'sh00001d7a;
	assign w_sys_tmp3012 = (w_sys_tmp3013 + r_run_k_17);
	assign w_sys_tmp3013 = 32'sh00001dfb;
	assign w_sys_tmp3018 = (w_sys_tmp3019 + r_run_k_17);
	assign w_sys_tmp3019 = 32'sh00001e7c;
	assign w_sys_tmp3024 = (w_sys_tmp3025 + r_run_k_17);
	assign w_sys_tmp3025 = 32'sh00001efd;
	assign w_sys_tmp3030 = (w_sys_tmp3031 + r_run_k_17);
	assign w_sys_tmp3031 = 32'sh00001f7e;
	assign w_sys_tmp3036 = (w_sys_tmp3037 + r_run_k_17);
	assign w_sys_tmp3037 = 32'sh00001fff;
	assign w_sys_tmp3042 = (w_sys_tmp3043 + r_run_k_17);
	assign w_sys_tmp3043 = 32'sh00002080;
	assign w_sys_tmp3048 = (w_sys_tmp3049 + r_run_k_17);
	assign w_sys_tmp3049 = 32'sh00002101;
	assign w_sys_tmp3066 = (w_sys_tmp3067 + r_run_k_17);
	assign w_sys_tmp3067 = 32'sh00002182;
	assign w_sys_tmp3072 = (w_sys_tmp3073 + r_run_k_17);
	assign w_sys_tmp3073 = 32'sh00002203;
	assign w_sys_tmp3078 = (w_sys_tmp3079 + r_run_k_17);
	assign w_sys_tmp3079 = 32'sh00002284;
	assign w_sys_tmp3084 = (w_sys_tmp3085 + r_run_k_17);
	assign w_sys_tmp3085 = 32'sh00002305;
	assign w_sys_tmp3090 = (w_sys_tmp3091 + r_run_k_17);
	assign w_sys_tmp3091 = 32'sh00002386;
	assign w_sys_tmp3096 = (w_sys_tmp3097 + r_run_k_17);
	assign w_sys_tmp3097 = 32'sh00002407;
	assign w_sys_tmp3102 = (w_sys_tmp3103 + r_run_k_17);
	assign w_sys_tmp3103 = 32'sh00002488;
	assign w_sys_tmp3108 = (w_sys_tmp3109 + r_run_k_17);
	assign w_sys_tmp3109 = 32'sh00002509;
	assign w_sys_tmp3114 = (w_sys_tmp3115 + r_run_k_17);
	assign w_sys_tmp3115 = 32'sh0000258a;
	assign w_sys_tmp3120 = (w_sys_tmp3121 + r_run_k_17);
	assign w_sys_tmp3121 = 32'sh0000260b;
	assign w_sys_tmp3126 = (w_sys_tmp3127 + r_run_k_17);
	assign w_sys_tmp3127 = 32'sh0000268c;
	assign w_sys_tmp3132 = (w_sys_tmp3133 + r_run_k_17);
	assign w_sys_tmp3133 = 32'sh0000270d;
	assign w_sys_tmp3138 = (w_sys_tmp3139 + r_run_k_17);
	assign w_sys_tmp3139 = 32'sh0000278e;
	assign w_sys_tmp3144 = (w_sys_tmp3145 + r_run_k_17);
	assign w_sys_tmp3145 = 32'sh0000280f;
	assign w_sys_tmp3150 = (w_sys_tmp3151 + r_run_k_17);
	assign w_sys_tmp3151 = 32'sh00002890;
	assign w_sys_tmp3156 = (w_sys_tmp3157 + r_run_k_17);
	assign w_sys_tmp3157 = 32'sh00002911;
	assign w_sys_tmp3162 = (w_sys_tmp3163 + r_run_k_17);
	assign w_sys_tmp3163 = 32'sh00002992;
	assign w_sys_tmp3168 = (w_sys_tmp3169 + r_run_k_17);
	assign w_sys_tmp3169 = 32'sh00002a13;
	assign w_sys_tmp3174 = (w_sys_tmp3175 + r_run_k_17);
	assign w_sys_tmp3175 = 32'sh00002a94;
	assign w_sys_tmp3180 = (w_sys_tmp3181 + r_run_k_17);
	assign w_sys_tmp3181 = 32'sh00002b15;
	assign w_sys_tmp3186 = (w_sys_tmp3187 + r_run_k_17);
	assign w_sys_tmp3187 = 32'sh00002b96;
	assign w_sys_tmp3192 = (w_sys_tmp3193 + r_run_k_17);
	assign w_sys_tmp3193 = 32'sh00002c17;
	assign w_sys_tmp3198 = (w_sys_tmp3199 + r_run_k_17);
	assign w_sys_tmp3199 = 32'sh00002c98;
	assign w_sys_tmp3204 = (w_sys_tmp3205 + r_run_k_17);
	assign w_sys_tmp3205 = 32'sh00002d19;
	assign w_sys_tmp3210 = (w_sys_tmp3211 + r_run_k_17);
	assign w_sys_tmp3211 = 32'sh00002d9a;
	assign w_sys_tmp3216 = (w_sys_tmp3217 + r_run_k_17);
	assign w_sys_tmp3217 = 32'sh00002e1b;
	assign w_sys_tmp3222 = (w_sys_tmp3223 + r_run_k_17);
	assign w_sys_tmp3223 = 32'sh00002e9c;
	assign w_sys_tmp3228 = (w_sys_tmp3229 + r_run_k_17);
	assign w_sys_tmp3229 = 32'sh00002f1d;
	assign w_sys_tmp3234 = (w_sys_tmp3235 + r_run_k_17);
	assign w_sys_tmp3235 = 32'sh00002f9e;
	assign w_sys_tmp3240 = (w_sys_tmp3241 + r_run_k_17);
	assign w_sys_tmp3241 = 32'sh0000301f;
	assign w_sys_tmp3246 = (w_sys_tmp3247 + r_run_k_17);
	assign w_sys_tmp3247 = 32'sh000030a0;
	assign w_sys_tmp3252 = (w_sys_tmp3253 + r_run_k_17);
	assign w_sys_tmp3253 = 32'sh00003121;
	assign w_sys_tmp3270 = (w_sys_tmp3271 + r_run_k_17);
	assign w_sys_tmp3271 = 32'sh000031a2;
	assign w_sys_tmp3276 = (w_sys_tmp3277 + r_run_k_17);
	assign w_sys_tmp3277 = 32'sh00003223;
	assign w_sys_tmp3282 = (w_sys_tmp3283 + r_run_k_17);
	assign w_sys_tmp3283 = 32'sh000032a4;
	assign w_sys_tmp3288 = (w_sys_tmp3289 + r_run_k_17);
	assign w_sys_tmp3289 = 32'sh00003325;
	assign w_sys_tmp3294 = (w_sys_tmp3295 + r_run_k_17);
	assign w_sys_tmp3295 = 32'sh000033a6;
	assign w_sys_tmp3300 = (w_sys_tmp3301 + r_run_k_17);
	assign w_sys_tmp3301 = 32'sh00003427;
	assign w_sys_tmp3306 = (w_sys_tmp3307 + r_run_k_17);
	assign w_sys_tmp3307 = 32'sh000034a8;
	assign w_sys_tmp3312 = (w_sys_tmp3313 + r_run_k_17);
	assign w_sys_tmp3313 = 32'sh00003529;
	assign w_sys_tmp3318 = (w_sys_tmp3319 + r_run_k_17);
	assign w_sys_tmp3319 = 32'sh000035aa;
	assign w_sys_tmp3324 = (w_sys_tmp3325 + r_run_k_17);
	assign w_sys_tmp3325 = 32'sh0000362b;
	assign w_sys_tmp3330 = (w_sys_tmp3331 + r_run_k_17);
	assign w_sys_tmp3331 = 32'sh000036ac;
	assign w_sys_tmp3336 = (w_sys_tmp3337 + r_run_k_17);
	assign w_sys_tmp3337 = 32'sh0000372d;
	assign w_sys_tmp3342 = (w_sys_tmp3343 + r_run_k_17);
	assign w_sys_tmp3343 = 32'sh000037ae;
	assign w_sys_tmp3348 = (w_sys_tmp3349 + r_run_k_17);
	assign w_sys_tmp3349 = 32'sh0000382f;
	assign w_sys_tmp3354 = (w_sys_tmp3355 + r_run_k_17);
	assign w_sys_tmp3355 = 32'sh000038b0;
	assign w_sys_tmp3360 = (w_sys_tmp3361 + r_run_k_17);
	assign w_sys_tmp3361 = 32'sh00003931;
	assign w_sys_tmp3366 = (w_sys_tmp3367 + r_run_k_17);
	assign w_sys_tmp3367 = 32'sh000039b2;
	assign w_sys_tmp3372 = (w_sys_tmp3373 + r_run_k_17);
	assign w_sys_tmp3373 = 32'sh00003a33;
	assign w_sys_tmp3378 = (w_sys_tmp3379 + r_run_k_17);
	assign w_sys_tmp3379 = 32'sh00003ab4;
	assign w_sys_tmp3384 = (w_sys_tmp3385 + r_run_k_17);
	assign w_sys_tmp3385 = 32'sh00003b35;
	assign w_sys_tmp3390 = (w_sys_tmp3391 + r_run_k_17);
	assign w_sys_tmp3391 = 32'sh00003bb6;
	assign w_sys_tmp3396 = (w_sys_tmp3397 + r_run_k_17);
	assign w_sys_tmp3397 = 32'sh00003c37;
	assign w_sys_tmp3402 = (w_sys_tmp3403 + r_run_k_17);
	assign w_sys_tmp3403 = 32'sh00003cb8;
	assign w_sys_tmp3408 = (w_sys_tmp3409 + r_run_k_17);
	assign w_sys_tmp3409 = 32'sh00003d39;
	assign w_sys_tmp3414 = (w_sys_tmp3415 + r_run_k_17);
	assign w_sys_tmp3415 = 32'sh00003dba;
	assign w_sys_tmp3420 = (w_sys_tmp3421 + r_run_k_17);
	assign w_sys_tmp3421 = 32'sh00003e3b;
	assign w_sys_tmp3426 = (w_sys_tmp3427 + r_run_k_17);
	assign w_sys_tmp3427 = 32'sh00003ebc;
	assign w_sys_tmp3432 = (w_sys_tmp3433 + r_run_k_17);
	assign w_sys_tmp3433 = 32'sh00003f3d;
	assign w_sys_tmp3438 = (w_sys_tmp3439 + r_run_k_17);
	assign w_sys_tmp3439 = 32'sh00003fbe;
	assign w_sys_tmp3444 = (w_sys_tmp3445 + r_run_k_17);
	assign w_sys_tmp3445 = 32'sh0000403f;
	assign w_sys_tmp3450 = (w_sys_tmp3451 + r_run_k_17);
	assign w_sys_tmp3451 = 32'sh000040c0;
	assign w_sys_tmp3456 = (w_sys_tmp3457 + r_run_k_17);
	assign w_sys_tmp3457 = 32'sh00004141;
	assign w_sys_tmp3461 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp3462 = 32'sh00000002;
	assign w_sys_tmp3463 = ( !w_sys_tmp3464 );
	assign w_sys_tmp3464 = (w_sys_tmp3465 < r_run_k_17);
	assign w_sys_tmp3465 = 32'sh00000020;
	assign w_sys_tmp3468 = (w_sys_tmp3469 + r_run_k_17);
	assign w_sys_tmp3469 = 32'sh00000102;
	assign w_sys_tmp3470 = w_sub00_result_dataout;
	assign w_sys_tmp3474 = (w_sys_tmp3475 + r_run_k_17);
	assign w_sys_tmp3475 = 32'sh00000183;
	assign w_sys_tmp3480 = (w_sys_tmp3481 + r_run_k_17);
	assign w_sys_tmp3481 = 32'sh00000204;
	assign w_sys_tmp3486 = (w_sys_tmp3487 + r_run_k_17);
	assign w_sys_tmp3487 = 32'sh00000285;
	assign w_sys_tmp3492 = (w_sys_tmp3493 + r_run_k_17);
	assign w_sys_tmp3493 = 32'sh00000306;
	assign w_sys_tmp3498 = (w_sys_tmp3499 + r_run_k_17);
	assign w_sys_tmp3499 = 32'sh00000387;
	assign w_sys_tmp3504 = (w_sys_tmp3505 + r_run_k_17);
	assign w_sys_tmp3505 = 32'sh00000408;
	assign w_sys_tmp3510 = (w_sys_tmp3511 + r_run_k_17);
	assign w_sys_tmp3511 = 32'sh00000489;
	assign w_sys_tmp3516 = (w_sys_tmp3517 + r_run_k_17);
	assign w_sys_tmp3517 = 32'sh0000050a;
	assign w_sys_tmp3522 = (w_sys_tmp3523 + r_run_k_17);
	assign w_sys_tmp3523 = 32'sh0000058b;
	assign w_sys_tmp3528 = (w_sys_tmp3529 + r_run_k_17);
	assign w_sys_tmp3529 = 32'sh0000060c;
	assign w_sys_tmp3534 = (w_sys_tmp3535 + r_run_k_17);
	assign w_sys_tmp3535 = 32'sh0000068d;
	assign w_sys_tmp3540 = (w_sys_tmp3541 + r_run_k_17);
	assign w_sys_tmp3541 = 32'sh0000070e;
	assign w_sys_tmp3546 = (w_sys_tmp3547 + r_run_k_17);
	assign w_sys_tmp3547 = 32'sh0000078f;
	assign w_sys_tmp3552 = (w_sys_tmp3553 + r_run_k_17);
	assign w_sys_tmp3553 = 32'sh00000810;
	assign w_sys_tmp3558 = (w_sys_tmp3559 + r_run_k_17);
	assign w_sys_tmp3559 = 32'sh00000891;
	assign w_sys_tmp3564 = (w_sys_tmp3565 + r_run_k_17);
	assign w_sys_tmp3565 = 32'sh00000912;
	assign w_sys_tmp3570 = (w_sys_tmp3571 + r_run_k_17);
	assign w_sys_tmp3571 = 32'sh00000993;
	assign w_sys_tmp3576 = (w_sys_tmp3577 + r_run_k_17);
	assign w_sys_tmp3577 = 32'sh00000a14;
	assign w_sys_tmp3582 = (w_sys_tmp3583 + r_run_k_17);
	assign w_sys_tmp3583 = 32'sh00000a95;
	assign w_sys_tmp3588 = (w_sys_tmp3589 + r_run_k_17);
	assign w_sys_tmp3589 = 32'sh00000b16;
	assign w_sys_tmp3594 = (w_sys_tmp3595 + r_run_k_17);
	assign w_sys_tmp3595 = 32'sh00000b97;
	assign w_sys_tmp3600 = (w_sys_tmp3601 + r_run_k_17);
	assign w_sys_tmp3601 = 32'sh00000c18;
	assign w_sys_tmp3606 = (w_sys_tmp3607 + r_run_k_17);
	assign w_sys_tmp3607 = 32'sh00000c99;
	assign w_sys_tmp3612 = (w_sys_tmp3613 + r_run_k_17);
	assign w_sys_tmp3613 = 32'sh00000d1a;
	assign w_sys_tmp3618 = (w_sys_tmp3619 + r_run_k_17);
	assign w_sys_tmp3619 = 32'sh00000d9b;
	assign w_sys_tmp3624 = (w_sys_tmp3625 + r_run_k_17);
	assign w_sys_tmp3625 = 32'sh00000e1c;
	assign w_sys_tmp3630 = (w_sys_tmp3631 + r_run_k_17);
	assign w_sys_tmp3631 = 32'sh00000e9d;
	assign w_sys_tmp3636 = (w_sys_tmp3637 + r_run_k_17);
	assign w_sys_tmp3637 = 32'sh00000f1e;
	assign w_sys_tmp3642 = (w_sys_tmp3643 + r_run_k_17);
	assign w_sys_tmp3643 = 32'sh00000f9f;
	assign w_sys_tmp3648 = (w_sys_tmp3649 + r_run_k_17);
	assign w_sys_tmp3649 = 32'sh00001020;
	assign w_sys_tmp3654 = (w_sys_tmp3655 + r_run_k_17);
	assign w_sys_tmp3655 = 32'sh000010a1;
	assign w_sys_tmp3659 = (w_sys_tmp3660 + r_run_k_17);
	assign w_sys_tmp3660 = 32'sh00001122;
	assign w_sys_tmp3664 = (w_sys_tmp3665 + r_run_k_17);
	assign w_sys_tmp3665 = 32'sh000011a3;
	assign w_sys_tmp3669 = (w_sys_tmp3670 + r_run_k_17);
	assign w_sys_tmp3670 = 32'sh00001224;
	assign w_sys_tmp3674 = (w_sys_tmp3675 + r_run_k_17);
	assign w_sys_tmp3675 = 32'sh000012a5;
	assign w_sys_tmp3679 = (w_sys_tmp3680 + r_run_k_17);
	assign w_sys_tmp3680 = 32'sh00001326;
	assign w_sys_tmp3684 = (w_sys_tmp3685 + r_run_k_17);
	assign w_sys_tmp3685 = 32'sh000013a7;
	assign w_sys_tmp3689 = (w_sys_tmp3690 + r_run_k_17);
	assign w_sys_tmp3690 = 32'sh00001428;
	assign w_sys_tmp3694 = (w_sys_tmp3695 + r_run_k_17);
	assign w_sys_tmp3695 = 32'sh000014a9;
	assign w_sys_tmp3699 = (w_sys_tmp3700 + r_run_k_17);
	assign w_sys_tmp3700 = 32'sh0000152a;
	assign w_sys_tmp3704 = (w_sys_tmp3705 + r_run_k_17);
	assign w_sys_tmp3705 = 32'sh000015ab;
	assign w_sys_tmp3709 = (w_sys_tmp3710 + r_run_k_17);
	assign w_sys_tmp3710 = 32'sh0000162c;
	assign w_sys_tmp3714 = (w_sys_tmp3715 + r_run_k_17);
	assign w_sys_tmp3715 = 32'sh000016ad;
	assign w_sys_tmp3719 = (w_sys_tmp3720 + r_run_k_17);
	assign w_sys_tmp3720 = 32'sh0000172e;
	assign w_sys_tmp3724 = (w_sys_tmp3725 + r_run_k_17);
	assign w_sys_tmp3725 = 32'sh000017af;
	assign w_sys_tmp3729 = (w_sys_tmp3730 + r_run_k_17);
	assign w_sys_tmp3730 = 32'sh00001830;
	assign w_sys_tmp3734 = (w_sys_tmp3735 + r_run_k_17);
	assign w_sys_tmp3735 = 32'sh000018b1;
	assign w_sys_tmp3739 = (w_sys_tmp3740 + r_run_k_17);
	assign w_sys_tmp3740 = 32'sh00001932;
	assign w_sys_tmp3744 = (w_sys_tmp3745 + r_run_k_17);
	assign w_sys_tmp3745 = 32'sh000019b3;
	assign w_sys_tmp3749 = (w_sys_tmp3750 + r_run_k_17);
	assign w_sys_tmp3750 = 32'sh00001a34;
	assign w_sys_tmp3754 = (w_sys_tmp3755 + r_run_k_17);
	assign w_sys_tmp3755 = 32'sh00001ab5;
	assign w_sys_tmp3759 = (w_sys_tmp3760 + r_run_k_17);
	assign w_sys_tmp3760 = 32'sh00001b36;
	assign w_sys_tmp3764 = (w_sys_tmp3765 + r_run_k_17);
	assign w_sys_tmp3765 = 32'sh00001bb7;
	assign w_sys_tmp3769 = (w_sys_tmp3770 + r_run_k_17);
	assign w_sys_tmp3770 = 32'sh00001c38;
	assign w_sys_tmp3774 = (w_sys_tmp3775 + r_run_k_17);
	assign w_sys_tmp3775 = 32'sh00001cb9;
	assign w_sys_tmp3779 = (w_sys_tmp3780 + r_run_k_17);
	assign w_sys_tmp3780 = 32'sh00001d3a;
	assign w_sys_tmp3784 = (w_sys_tmp3785 + r_run_k_17);
	assign w_sys_tmp3785 = 32'sh00001dbb;
	assign w_sys_tmp3789 = (w_sys_tmp3790 + r_run_k_17);
	assign w_sys_tmp3790 = 32'sh00001e3c;
	assign w_sys_tmp3794 = (w_sys_tmp3795 + r_run_k_17);
	assign w_sys_tmp3795 = 32'sh00001ebd;
	assign w_sys_tmp3799 = (w_sys_tmp3800 + r_run_k_17);
	assign w_sys_tmp3800 = 32'sh00001f3e;
	assign w_sys_tmp3804 = (w_sys_tmp3805 + r_run_k_17);
	assign w_sys_tmp3805 = 32'sh00001fbf;
	assign w_sys_tmp3809 = (w_sys_tmp3810 + r_run_k_17);
	assign w_sys_tmp3810 = 32'sh00002040;
	assign w_sys_tmp3814 = (w_sys_tmp3815 + r_run_k_17);
	assign w_sys_tmp3815 = 32'sh000020c1;
	assign w_sys_tmp3819 = (w_sys_tmp3820 + r_run_k_17);
	assign w_sys_tmp3820 = 32'sh00002142;
	assign w_sys_tmp3824 = (w_sys_tmp3825 + r_run_k_17);
	assign w_sys_tmp3825 = 32'sh000021c3;
	assign w_sys_tmp3829 = (w_sys_tmp3830 + r_run_k_17);
	assign w_sys_tmp3830 = 32'sh00002244;
	assign w_sys_tmp3834 = (w_sys_tmp3835 + r_run_k_17);
	assign w_sys_tmp3835 = 32'sh000022c5;
	assign w_sys_tmp3839 = (w_sys_tmp3840 + r_run_k_17);
	assign w_sys_tmp3840 = 32'sh00002346;
	assign w_sys_tmp3844 = (w_sys_tmp3845 + r_run_k_17);
	assign w_sys_tmp3845 = 32'sh000023c7;
	assign w_sys_tmp3849 = (w_sys_tmp3850 + r_run_k_17);
	assign w_sys_tmp3850 = 32'sh00002448;
	assign w_sys_tmp3854 = (w_sys_tmp3855 + r_run_k_17);
	assign w_sys_tmp3855 = 32'sh000024c9;
	assign w_sys_tmp3859 = (w_sys_tmp3860 + r_run_k_17);
	assign w_sys_tmp3860 = 32'sh0000254a;
	assign w_sys_tmp3864 = (w_sys_tmp3865 + r_run_k_17);
	assign w_sys_tmp3865 = 32'sh000025cb;
	assign w_sys_tmp3869 = (w_sys_tmp3870 + r_run_k_17);
	assign w_sys_tmp3870 = 32'sh0000264c;
	assign w_sys_tmp3874 = (w_sys_tmp3875 + r_run_k_17);
	assign w_sys_tmp3875 = 32'sh000026cd;
	assign w_sys_tmp3879 = (w_sys_tmp3880 + r_run_k_17);
	assign w_sys_tmp3880 = 32'sh0000274e;
	assign w_sys_tmp3884 = (w_sys_tmp3885 + r_run_k_17);
	assign w_sys_tmp3885 = 32'sh000027cf;
	assign w_sys_tmp3889 = (w_sys_tmp3890 + r_run_k_17);
	assign w_sys_tmp3890 = 32'sh00002850;
	assign w_sys_tmp3894 = (w_sys_tmp3895 + r_run_k_17);
	assign w_sys_tmp3895 = 32'sh000028d1;
	assign w_sys_tmp3899 = (w_sys_tmp3900 + r_run_k_17);
	assign w_sys_tmp3900 = 32'sh00002952;
	assign w_sys_tmp3904 = (w_sys_tmp3905 + r_run_k_17);
	assign w_sys_tmp3905 = 32'sh000029d3;
	assign w_sys_tmp3909 = (w_sys_tmp3910 + r_run_k_17);
	assign w_sys_tmp3910 = 32'sh00002a54;
	assign w_sys_tmp3914 = (w_sys_tmp3915 + r_run_k_17);
	assign w_sys_tmp3915 = 32'sh00002ad5;
	assign w_sys_tmp3919 = (w_sys_tmp3920 + r_run_k_17);
	assign w_sys_tmp3920 = 32'sh00002b56;
	assign w_sys_tmp3924 = (w_sys_tmp3925 + r_run_k_17);
	assign w_sys_tmp3925 = 32'sh00002bd7;
	assign w_sys_tmp3929 = (w_sys_tmp3930 + r_run_k_17);
	assign w_sys_tmp3930 = 32'sh00002c58;
	assign w_sys_tmp3934 = (w_sys_tmp3935 + r_run_k_17);
	assign w_sys_tmp3935 = 32'sh00002cd9;
	assign w_sys_tmp3939 = (w_sys_tmp3940 + r_run_k_17);
	assign w_sys_tmp3940 = 32'sh00002d5a;
	assign w_sys_tmp3944 = (w_sys_tmp3945 + r_run_k_17);
	assign w_sys_tmp3945 = 32'sh00002ddb;
	assign w_sys_tmp3949 = (w_sys_tmp3950 + r_run_k_17);
	assign w_sys_tmp3950 = 32'sh00002e5c;
	assign w_sys_tmp3954 = (w_sys_tmp3955 + r_run_k_17);
	assign w_sys_tmp3955 = 32'sh00002edd;
	assign w_sys_tmp3959 = (w_sys_tmp3960 + r_run_k_17);
	assign w_sys_tmp3960 = 32'sh00002f5e;
	assign w_sys_tmp3964 = (w_sys_tmp3965 + r_run_k_17);
	assign w_sys_tmp3965 = 32'sh00002fdf;
	assign w_sys_tmp3969 = (w_sys_tmp3970 + r_run_k_17);
	assign w_sys_tmp3970 = 32'sh00003060;
	assign w_sys_tmp3974 = (w_sys_tmp3975 + r_run_k_17);
	assign w_sys_tmp3975 = 32'sh000030e1;
	assign w_sys_tmp3979 = (w_sys_tmp3980 + r_run_k_17);
	assign w_sys_tmp3980 = 32'sh00003162;
	assign w_sys_tmp3984 = (w_sys_tmp3985 + r_run_k_17);
	assign w_sys_tmp3985 = 32'sh000031e3;
	assign w_sys_tmp3989 = (w_sys_tmp3990 + r_run_k_17);
	assign w_sys_tmp3990 = 32'sh00003264;
	assign w_sys_tmp3994 = (w_sys_tmp3995 + r_run_k_17);
	assign w_sys_tmp3995 = 32'sh000032e5;
	assign w_sys_tmp3999 = (w_sys_tmp4000 + r_run_k_17);
	assign w_sys_tmp4000 = 32'sh00003366;
	assign w_sys_tmp4004 = (w_sys_tmp4005 + r_run_k_17);
	assign w_sys_tmp4005 = 32'sh000033e7;
	assign w_sys_tmp4009 = (w_sys_tmp4010 + r_run_k_17);
	assign w_sys_tmp4010 = 32'sh00003468;
	assign w_sys_tmp4014 = (w_sys_tmp4015 + r_run_k_17);
	assign w_sys_tmp4015 = 32'sh000034e9;
	assign w_sys_tmp4019 = (w_sys_tmp4020 + r_run_k_17);
	assign w_sys_tmp4020 = 32'sh0000356a;
	assign w_sys_tmp4024 = (w_sys_tmp4025 + r_run_k_17);
	assign w_sys_tmp4025 = 32'sh000035eb;
	assign w_sys_tmp4029 = (w_sys_tmp4030 + r_run_k_17);
	assign w_sys_tmp4030 = 32'sh0000366c;
	assign w_sys_tmp4034 = (w_sys_tmp4035 + r_run_k_17);
	assign w_sys_tmp4035 = 32'sh000036ed;
	assign w_sys_tmp4039 = (w_sys_tmp4040 + r_run_k_17);
	assign w_sys_tmp4040 = 32'sh0000376e;
	assign w_sys_tmp4044 = (w_sys_tmp4045 + r_run_k_17);
	assign w_sys_tmp4045 = 32'sh000037ef;
	assign w_sys_tmp4049 = (w_sys_tmp4050 + r_run_k_17);
	assign w_sys_tmp4050 = 32'sh00003870;
	assign w_sys_tmp4054 = (w_sys_tmp4055 + r_run_k_17);
	assign w_sys_tmp4055 = 32'sh000038f1;
	assign w_sys_tmp4059 = (w_sys_tmp4060 + r_run_k_17);
	assign w_sys_tmp4060 = 32'sh00003972;
	assign w_sys_tmp4064 = (w_sys_tmp4065 + r_run_k_17);
	assign w_sys_tmp4065 = 32'sh000039f3;
	assign w_sys_tmp4069 = (w_sys_tmp4070 + r_run_k_17);
	assign w_sys_tmp4070 = 32'sh00003a74;
	assign w_sys_tmp4074 = (w_sys_tmp4075 + r_run_k_17);
	assign w_sys_tmp4075 = 32'sh00003af5;
	assign w_sys_tmp4079 = (w_sys_tmp4080 + r_run_k_17);
	assign w_sys_tmp4080 = 32'sh00003b76;
	assign w_sys_tmp4084 = (w_sys_tmp4085 + r_run_k_17);
	assign w_sys_tmp4085 = 32'sh00003bf7;
	assign w_sys_tmp4089 = (w_sys_tmp4090 + r_run_k_17);
	assign w_sys_tmp4090 = 32'sh00003c78;
	assign w_sys_tmp4094 = (w_sys_tmp4095 + r_run_k_17);
	assign w_sys_tmp4095 = 32'sh00003cf9;
	assign w_sys_tmp4099 = (w_sys_tmp4100 + r_run_k_17);
	assign w_sys_tmp4100 = 32'sh00003d7a;
	assign w_sys_tmp4104 = (w_sys_tmp4105 + r_run_k_17);
	assign w_sys_tmp4105 = 32'sh00003dfb;
	assign w_sys_tmp4109 = (w_sys_tmp4110 + r_run_k_17);
	assign w_sys_tmp4110 = 32'sh00003e7c;
	assign w_sys_tmp4114 = (w_sys_tmp4115 + r_run_k_17);
	assign w_sys_tmp4115 = 32'sh00003efd;
	assign w_sys_tmp4119 = (w_sys_tmp4120 + r_run_k_17);
	assign w_sys_tmp4120 = 32'sh00003f7e;
	assign w_sys_tmp4124 = (w_sys_tmp4125 + r_run_k_17);
	assign w_sys_tmp4125 = 32'sh00003fff;
	assign w_sys_tmp4129 = (w_sys_tmp4130 + r_run_k_17);
	assign w_sys_tmp4130 = 32'sh00004080;
	assign w_sys_tmp4133 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp4134 = 32'sh00000006;
	assign w_sys_tmp4135 = ( !w_sys_tmp4136 );
	assign w_sys_tmp4136 = (w_sys_tmp4137 < r_run_k_17);
	assign w_sys_tmp4137 = 32'sh00000040;
	assign w_sys_tmp4140 = (w_sys_tmp4141 + r_run_k_17);
	assign w_sys_tmp4141 = 32'sh00000102;
	assign w_sys_tmp4142 = w_sub04_result_dataout;
	assign w_sys_tmp4146 = (w_sys_tmp4147 + r_run_k_17);
	assign w_sys_tmp4147 = 32'sh00000183;
	assign w_sys_tmp4152 = (w_sys_tmp4153 + r_run_k_17);
	assign w_sys_tmp4153 = 32'sh00000204;
	assign w_sys_tmp4158 = (w_sys_tmp4159 + r_run_k_17);
	assign w_sys_tmp4159 = 32'sh00000285;
	assign w_sys_tmp4164 = (w_sys_tmp4165 + r_run_k_17);
	assign w_sys_tmp4165 = 32'sh00000306;
	assign w_sys_tmp4170 = (w_sys_tmp4171 + r_run_k_17);
	assign w_sys_tmp4171 = 32'sh00000387;
	assign w_sys_tmp4176 = (w_sys_tmp4177 + r_run_k_17);
	assign w_sys_tmp4177 = 32'sh00000408;
	assign w_sys_tmp4182 = (w_sys_tmp4183 + r_run_k_17);
	assign w_sys_tmp4183 = 32'sh00000489;
	assign w_sys_tmp4188 = (w_sys_tmp4189 + r_run_k_17);
	assign w_sys_tmp4189 = 32'sh0000050a;
	assign w_sys_tmp4194 = (w_sys_tmp4195 + r_run_k_17);
	assign w_sys_tmp4195 = 32'sh0000058b;
	assign w_sys_tmp4200 = (w_sys_tmp4201 + r_run_k_17);
	assign w_sys_tmp4201 = 32'sh0000060c;
	assign w_sys_tmp4206 = (w_sys_tmp4207 + r_run_k_17);
	assign w_sys_tmp4207 = 32'sh0000068d;
	assign w_sys_tmp4212 = (w_sys_tmp4213 + r_run_k_17);
	assign w_sys_tmp4213 = 32'sh0000070e;
	assign w_sys_tmp4218 = (w_sys_tmp4219 + r_run_k_17);
	assign w_sys_tmp4219 = 32'sh0000078f;
	assign w_sys_tmp4224 = (w_sys_tmp4225 + r_run_k_17);
	assign w_sys_tmp4225 = 32'sh00000810;
	assign w_sys_tmp4230 = (w_sys_tmp4231 + r_run_k_17);
	assign w_sys_tmp4231 = 32'sh00000891;
	assign w_sys_tmp4236 = (w_sys_tmp4237 + r_run_k_17);
	assign w_sys_tmp4237 = 32'sh00000912;
	assign w_sys_tmp4242 = (w_sys_tmp4243 + r_run_k_17);
	assign w_sys_tmp4243 = 32'sh00000993;
	assign w_sys_tmp4248 = (w_sys_tmp4249 + r_run_k_17);
	assign w_sys_tmp4249 = 32'sh00000a14;
	assign w_sys_tmp4254 = (w_sys_tmp4255 + r_run_k_17);
	assign w_sys_tmp4255 = 32'sh00000a95;
	assign w_sys_tmp4260 = (w_sys_tmp4261 + r_run_k_17);
	assign w_sys_tmp4261 = 32'sh00000b16;
	assign w_sys_tmp4266 = (w_sys_tmp4267 + r_run_k_17);
	assign w_sys_tmp4267 = 32'sh00000b97;
	assign w_sys_tmp4272 = (w_sys_tmp4273 + r_run_k_17);
	assign w_sys_tmp4273 = 32'sh00000c18;
	assign w_sys_tmp4278 = (w_sys_tmp4279 + r_run_k_17);
	assign w_sys_tmp4279 = 32'sh00000c99;
	assign w_sys_tmp4284 = (w_sys_tmp4285 + r_run_k_17);
	assign w_sys_tmp4285 = 32'sh00000d1a;
	assign w_sys_tmp4290 = (w_sys_tmp4291 + r_run_k_17);
	assign w_sys_tmp4291 = 32'sh00000d9b;
	assign w_sys_tmp4296 = (w_sys_tmp4297 + r_run_k_17);
	assign w_sys_tmp4297 = 32'sh00000e1c;
	assign w_sys_tmp4302 = (w_sys_tmp4303 + r_run_k_17);
	assign w_sys_tmp4303 = 32'sh00000e9d;
	assign w_sys_tmp4308 = (w_sys_tmp4309 + r_run_k_17);
	assign w_sys_tmp4309 = 32'sh00000f1e;
	assign w_sys_tmp4314 = (w_sys_tmp4315 + r_run_k_17);
	assign w_sys_tmp4315 = 32'sh00000f9f;
	assign w_sys_tmp4320 = (w_sys_tmp4321 + r_run_k_17);
	assign w_sys_tmp4321 = 32'sh00001020;
	assign w_sys_tmp4326 = (w_sys_tmp4327 + r_run_k_17);
	assign w_sys_tmp4327 = 32'sh000010a1;
	assign w_sys_tmp4331 = (w_sys_tmp4332 + r_run_k_17);
	assign w_sys_tmp4332 = 32'sh00001122;
	assign w_sys_tmp4336 = (w_sys_tmp4337 + r_run_k_17);
	assign w_sys_tmp4337 = 32'sh000011a3;
	assign w_sys_tmp4341 = (w_sys_tmp4342 + r_run_k_17);
	assign w_sys_tmp4342 = 32'sh00001224;
	assign w_sys_tmp4346 = (w_sys_tmp4347 + r_run_k_17);
	assign w_sys_tmp4347 = 32'sh000012a5;
	assign w_sys_tmp4351 = (w_sys_tmp4352 + r_run_k_17);
	assign w_sys_tmp4352 = 32'sh00001326;
	assign w_sys_tmp4356 = (w_sys_tmp4357 + r_run_k_17);
	assign w_sys_tmp4357 = 32'sh000013a7;
	assign w_sys_tmp4361 = (w_sys_tmp4362 + r_run_k_17);
	assign w_sys_tmp4362 = 32'sh00001428;
	assign w_sys_tmp4366 = (w_sys_tmp4367 + r_run_k_17);
	assign w_sys_tmp4367 = 32'sh000014a9;
	assign w_sys_tmp4371 = (w_sys_tmp4372 + r_run_k_17);
	assign w_sys_tmp4372 = 32'sh0000152a;
	assign w_sys_tmp4376 = (w_sys_tmp4377 + r_run_k_17);
	assign w_sys_tmp4377 = 32'sh000015ab;
	assign w_sys_tmp4381 = (w_sys_tmp4382 + r_run_k_17);
	assign w_sys_tmp4382 = 32'sh0000162c;
	assign w_sys_tmp4386 = (w_sys_tmp4387 + r_run_k_17);
	assign w_sys_tmp4387 = 32'sh000016ad;
	assign w_sys_tmp4391 = (w_sys_tmp4392 + r_run_k_17);
	assign w_sys_tmp4392 = 32'sh0000172e;
	assign w_sys_tmp4396 = (w_sys_tmp4397 + r_run_k_17);
	assign w_sys_tmp4397 = 32'sh000017af;
	assign w_sys_tmp4401 = (w_sys_tmp4402 + r_run_k_17);
	assign w_sys_tmp4402 = 32'sh00001830;
	assign w_sys_tmp4406 = (w_sys_tmp4407 + r_run_k_17);
	assign w_sys_tmp4407 = 32'sh000018b1;
	assign w_sys_tmp4411 = (w_sys_tmp4412 + r_run_k_17);
	assign w_sys_tmp4412 = 32'sh00001932;
	assign w_sys_tmp4416 = (w_sys_tmp4417 + r_run_k_17);
	assign w_sys_tmp4417 = 32'sh000019b3;
	assign w_sys_tmp4421 = (w_sys_tmp4422 + r_run_k_17);
	assign w_sys_tmp4422 = 32'sh00001a34;
	assign w_sys_tmp4426 = (w_sys_tmp4427 + r_run_k_17);
	assign w_sys_tmp4427 = 32'sh00001ab5;
	assign w_sys_tmp4431 = (w_sys_tmp4432 + r_run_k_17);
	assign w_sys_tmp4432 = 32'sh00001b36;
	assign w_sys_tmp4436 = (w_sys_tmp4437 + r_run_k_17);
	assign w_sys_tmp4437 = 32'sh00001bb7;
	assign w_sys_tmp4441 = (w_sys_tmp4442 + r_run_k_17);
	assign w_sys_tmp4442 = 32'sh00001c38;
	assign w_sys_tmp4446 = (w_sys_tmp4447 + r_run_k_17);
	assign w_sys_tmp4447 = 32'sh00001cb9;
	assign w_sys_tmp4451 = (w_sys_tmp4452 + r_run_k_17);
	assign w_sys_tmp4452 = 32'sh00001d3a;
	assign w_sys_tmp4456 = (w_sys_tmp4457 + r_run_k_17);
	assign w_sys_tmp4457 = 32'sh00001dbb;
	assign w_sys_tmp4461 = (w_sys_tmp4462 + r_run_k_17);
	assign w_sys_tmp4462 = 32'sh00001e3c;
	assign w_sys_tmp4466 = (w_sys_tmp4467 + r_run_k_17);
	assign w_sys_tmp4467 = 32'sh00001ebd;
	assign w_sys_tmp4471 = (w_sys_tmp4472 + r_run_k_17);
	assign w_sys_tmp4472 = 32'sh00001f3e;
	assign w_sys_tmp4476 = (w_sys_tmp4477 + r_run_k_17);
	assign w_sys_tmp4477 = 32'sh00001fbf;
	assign w_sys_tmp4481 = (w_sys_tmp4482 + r_run_k_17);
	assign w_sys_tmp4482 = 32'sh00002040;
	assign w_sys_tmp4486 = (w_sys_tmp4487 + r_run_k_17);
	assign w_sys_tmp4487 = 32'sh000020c1;
	assign w_sys_tmp4491 = (w_sys_tmp4492 + r_run_k_17);
	assign w_sys_tmp4492 = 32'sh00002142;
	assign w_sys_tmp4496 = (w_sys_tmp4497 + r_run_k_17);
	assign w_sys_tmp4497 = 32'sh000021c3;
	assign w_sys_tmp4501 = (w_sys_tmp4502 + r_run_k_17);
	assign w_sys_tmp4502 = 32'sh00002244;
	assign w_sys_tmp4506 = (w_sys_tmp4507 + r_run_k_17);
	assign w_sys_tmp4507 = 32'sh000022c5;
	assign w_sys_tmp4511 = (w_sys_tmp4512 + r_run_k_17);
	assign w_sys_tmp4512 = 32'sh00002346;
	assign w_sys_tmp4516 = (w_sys_tmp4517 + r_run_k_17);
	assign w_sys_tmp4517 = 32'sh000023c7;
	assign w_sys_tmp4521 = (w_sys_tmp4522 + r_run_k_17);
	assign w_sys_tmp4522 = 32'sh00002448;
	assign w_sys_tmp4526 = (w_sys_tmp4527 + r_run_k_17);
	assign w_sys_tmp4527 = 32'sh000024c9;
	assign w_sys_tmp4531 = (w_sys_tmp4532 + r_run_k_17);
	assign w_sys_tmp4532 = 32'sh0000254a;
	assign w_sys_tmp4536 = (w_sys_tmp4537 + r_run_k_17);
	assign w_sys_tmp4537 = 32'sh000025cb;
	assign w_sys_tmp4541 = (w_sys_tmp4542 + r_run_k_17);
	assign w_sys_tmp4542 = 32'sh0000264c;
	assign w_sys_tmp4546 = (w_sys_tmp4547 + r_run_k_17);
	assign w_sys_tmp4547 = 32'sh000026cd;
	assign w_sys_tmp4551 = (w_sys_tmp4552 + r_run_k_17);
	assign w_sys_tmp4552 = 32'sh0000274e;
	assign w_sys_tmp4556 = (w_sys_tmp4557 + r_run_k_17);
	assign w_sys_tmp4557 = 32'sh000027cf;
	assign w_sys_tmp4561 = (w_sys_tmp4562 + r_run_k_17);
	assign w_sys_tmp4562 = 32'sh00002850;
	assign w_sys_tmp4566 = (w_sys_tmp4567 + r_run_k_17);
	assign w_sys_tmp4567 = 32'sh000028d1;
	assign w_sys_tmp4571 = (w_sys_tmp4572 + r_run_k_17);
	assign w_sys_tmp4572 = 32'sh00002952;
	assign w_sys_tmp4576 = (w_sys_tmp4577 + r_run_k_17);
	assign w_sys_tmp4577 = 32'sh000029d3;
	assign w_sys_tmp4581 = (w_sys_tmp4582 + r_run_k_17);
	assign w_sys_tmp4582 = 32'sh00002a54;
	assign w_sys_tmp4586 = (w_sys_tmp4587 + r_run_k_17);
	assign w_sys_tmp4587 = 32'sh00002ad5;
	assign w_sys_tmp4591 = (w_sys_tmp4592 + r_run_k_17);
	assign w_sys_tmp4592 = 32'sh00002b56;
	assign w_sys_tmp4596 = (w_sys_tmp4597 + r_run_k_17);
	assign w_sys_tmp4597 = 32'sh00002bd7;
	assign w_sys_tmp4601 = (w_sys_tmp4602 + r_run_k_17);
	assign w_sys_tmp4602 = 32'sh00002c58;
	assign w_sys_tmp4606 = (w_sys_tmp4607 + r_run_k_17);
	assign w_sys_tmp4607 = 32'sh00002cd9;
	assign w_sys_tmp4611 = (w_sys_tmp4612 + r_run_k_17);
	assign w_sys_tmp4612 = 32'sh00002d5a;
	assign w_sys_tmp4616 = (w_sys_tmp4617 + r_run_k_17);
	assign w_sys_tmp4617 = 32'sh00002ddb;
	assign w_sys_tmp4621 = (w_sys_tmp4622 + r_run_k_17);
	assign w_sys_tmp4622 = 32'sh00002e5c;
	assign w_sys_tmp4626 = (w_sys_tmp4627 + r_run_k_17);
	assign w_sys_tmp4627 = 32'sh00002edd;
	assign w_sys_tmp4631 = (w_sys_tmp4632 + r_run_k_17);
	assign w_sys_tmp4632 = 32'sh00002f5e;
	assign w_sys_tmp4636 = (w_sys_tmp4637 + r_run_k_17);
	assign w_sys_tmp4637 = 32'sh00002fdf;
	assign w_sys_tmp4641 = (w_sys_tmp4642 + r_run_k_17);
	assign w_sys_tmp4642 = 32'sh00003060;
	assign w_sys_tmp4646 = (w_sys_tmp4647 + r_run_k_17);
	assign w_sys_tmp4647 = 32'sh000030e1;
	assign w_sys_tmp4651 = (w_sys_tmp4652 + r_run_k_17);
	assign w_sys_tmp4652 = 32'sh00003162;
	assign w_sys_tmp4656 = (w_sys_tmp4657 + r_run_k_17);
	assign w_sys_tmp4657 = 32'sh000031e3;
	assign w_sys_tmp4661 = (w_sys_tmp4662 + r_run_k_17);
	assign w_sys_tmp4662 = 32'sh00003264;
	assign w_sys_tmp4666 = (w_sys_tmp4667 + r_run_k_17);
	assign w_sys_tmp4667 = 32'sh000032e5;
	assign w_sys_tmp4671 = (w_sys_tmp4672 + r_run_k_17);
	assign w_sys_tmp4672 = 32'sh00003366;
	assign w_sys_tmp4676 = (w_sys_tmp4677 + r_run_k_17);
	assign w_sys_tmp4677 = 32'sh000033e7;
	assign w_sys_tmp4681 = (w_sys_tmp4682 + r_run_k_17);
	assign w_sys_tmp4682 = 32'sh00003468;
	assign w_sys_tmp4686 = (w_sys_tmp4687 + r_run_k_17);
	assign w_sys_tmp4687 = 32'sh000034e9;
	assign w_sys_tmp4691 = (w_sys_tmp4692 + r_run_k_17);
	assign w_sys_tmp4692 = 32'sh0000356a;
	assign w_sys_tmp4696 = (w_sys_tmp4697 + r_run_k_17);
	assign w_sys_tmp4697 = 32'sh000035eb;
	assign w_sys_tmp4701 = (w_sys_tmp4702 + r_run_k_17);
	assign w_sys_tmp4702 = 32'sh0000366c;
	assign w_sys_tmp4706 = (w_sys_tmp4707 + r_run_k_17);
	assign w_sys_tmp4707 = 32'sh000036ed;
	assign w_sys_tmp4711 = (w_sys_tmp4712 + r_run_k_17);
	assign w_sys_tmp4712 = 32'sh0000376e;
	assign w_sys_tmp4716 = (w_sys_tmp4717 + r_run_k_17);
	assign w_sys_tmp4717 = 32'sh000037ef;
	assign w_sys_tmp4721 = (w_sys_tmp4722 + r_run_k_17);
	assign w_sys_tmp4722 = 32'sh00003870;
	assign w_sys_tmp4726 = (w_sys_tmp4727 + r_run_k_17);
	assign w_sys_tmp4727 = 32'sh000038f1;
	assign w_sys_tmp4731 = (w_sys_tmp4732 + r_run_k_17);
	assign w_sys_tmp4732 = 32'sh00003972;
	assign w_sys_tmp4736 = (w_sys_tmp4737 + r_run_k_17);
	assign w_sys_tmp4737 = 32'sh000039f3;
	assign w_sys_tmp4741 = (w_sys_tmp4742 + r_run_k_17);
	assign w_sys_tmp4742 = 32'sh00003a74;
	assign w_sys_tmp4746 = (w_sys_tmp4747 + r_run_k_17);
	assign w_sys_tmp4747 = 32'sh00003af5;
	assign w_sys_tmp4751 = (w_sys_tmp4752 + r_run_k_17);
	assign w_sys_tmp4752 = 32'sh00003b76;
	assign w_sys_tmp4756 = (w_sys_tmp4757 + r_run_k_17);
	assign w_sys_tmp4757 = 32'sh00003bf7;
	assign w_sys_tmp4761 = (w_sys_tmp4762 + r_run_k_17);
	assign w_sys_tmp4762 = 32'sh00003c78;
	assign w_sys_tmp4766 = (w_sys_tmp4767 + r_run_k_17);
	assign w_sys_tmp4767 = 32'sh00003cf9;
	assign w_sys_tmp4771 = (w_sys_tmp4772 + r_run_k_17);
	assign w_sys_tmp4772 = 32'sh00003d7a;
	assign w_sys_tmp4776 = (w_sys_tmp4777 + r_run_k_17);
	assign w_sys_tmp4777 = 32'sh00003dfb;
	assign w_sys_tmp4781 = (w_sys_tmp4782 + r_run_k_17);
	assign w_sys_tmp4782 = 32'sh00003e7c;
	assign w_sys_tmp4786 = (w_sys_tmp4787 + r_run_k_17);
	assign w_sys_tmp4787 = 32'sh00003efd;
	assign w_sys_tmp4791 = (w_sys_tmp4792 + r_run_k_17);
	assign w_sys_tmp4792 = 32'sh00003f7e;
	assign w_sys_tmp4796 = (w_sys_tmp4797 + r_run_k_17);
	assign w_sys_tmp4797 = 32'sh00003fff;
	assign w_sys_tmp4801 = (w_sys_tmp4802 + r_run_k_17);
	assign w_sys_tmp4802 = 32'sh00004080;
	assign w_sys_tmp4806 = (w_sys_tmp4807 + r_run_k_17);
	assign w_sys_tmp4807 = 32'sh00000122;
	assign w_sys_tmp4811 = (w_sys_tmp4812 + r_run_k_17);
	assign w_sys_tmp4812 = 32'sh000001a3;
	assign w_sys_tmp4816 = (w_sys_tmp4817 + r_run_k_17);
	assign w_sys_tmp4817 = 32'sh00000224;
	assign w_sys_tmp4821 = (w_sys_tmp4822 + r_run_k_17);
	assign w_sys_tmp4822 = 32'sh000002a5;
	assign w_sys_tmp4826 = (w_sys_tmp4827 + r_run_k_17);
	assign w_sys_tmp4827 = 32'sh00000326;
	assign w_sys_tmp4831 = (w_sys_tmp4832 + r_run_k_17);
	assign w_sys_tmp4832 = 32'sh000003a7;
	assign w_sys_tmp4836 = (w_sys_tmp4837 + r_run_k_17);
	assign w_sys_tmp4837 = 32'sh00000428;
	assign w_sys_tmp4841 = (w_sys_tmp4842 + r_run_k_17);
	assign w_sys_tmp4842 = 32'sh000004a9;
	assign w_sys_tmp4846 = (w_sys_tmp4847 + r_run_k_17);
	assign w_sys_tmp4847 = 32'sh0000052a;
	assign w_sys_tmp4851 = (w_sys_tmp4852 + r_run_k_17);
	assign w_sys_tmp4852 = 32'sh000005ab;
	assign w_sys_tmp4856 = (w_sys_tmp4857 + r_run_k_17);
	assign w_sys_tmp4857 = 32'sh0000062c;
	assign w_sys_tmp4861 = (w_sys_tmp4862 + r_run_k_17);
	assign w_sys_tmp4862 = 32'sh000006ad;
	assign w_sys_tmp4866 = (w_sys_tmp4867 + r_run_k_17);
	assign w_sys_tmp4867 = 32'sh0000072e;
	assign w_sys_tmp4871 = (w_sys_tmp4872 + r_run_k_17);
	assign w_sys_tmp4872 = 32'sh000007af;
	assign w_sys_tmp4876 = (w_sys_tmp4877 + r_run_k_17);
	assign w_sys_tmp4877 = 32'sh00000830;
	assign w_sys_tmp4881 = (w_sys_tmp4882 + r_run_k_17);
	assign w_sys_tmp4882 = 32'sh000008b1;
	assign w_sys_tmp4886 = (w_sys_tmp4887 + r_run_k_17);
	assign w_sys_tmp4887 = 32'sh00000932;
	assign w_sys_tmp4891 = (w_sys_tmp4892 + r_run_k_17);
	assign w_sys_tmp4892 = 32'sh000009b3;
	assign w_sys_tmp4896 = (w_sys_tmp4897 + r_run_k_17);
	assign w_sys_tmp4897 = 32'sh00000a34;
	assign w_sys_tmp4901 = (w_sys_tmp4902 + r_run_k_17);
	assign w_sys_tmp4902 = 32'sh00000ab5;
	assign w_sys_tmp4906 = (w_sys_tmp4907 + r_run_k_17);
	assign w_sys_tmp4907 = 32'sh00000b36;
	assign w_sys_tmp4911 = (w_sys_tmp4912 + r_run_k_17);
	assign w_sys_tmp4912 = 32'sh00000bb7;
	assign w_sys_tmp4916 = (w_sys_tmp4917 + r_run_k_17);
	assign w_sys_tmp4917 = 32'sh00000c38;
	assign w_sys_tmp4921 = (w_sys_tmp4922 + r_run_k_17);
	assign w_sys_tmp4922 = 32'sh00000cb9;
	assign w_sys_tmp4926 = (w_sys_tmp4927 + r_run_k_17);
	assign w_sys_tmp4927 = 32'sh00000d3a;
	assign w_sys_tmp4931 = (w_sys_tmp4932 + r_run_k_17);
	assign w_sys_tmp4932 = 32'sh00000dbb;
	assign w_sys_tmp4936 = (w_sys_tmp4937 + r_run_k_17);
	assign w_sys_tmp4937 = 32'sh00000e3c;
	assign w_sys_tmp4941 = (w_sys_tmp4942 + r_run_k_17);
	assign w_sys_tmp4942 = 32'sh00000ebd;
	assign w_sys_tmp4946 = (w_sys_tmp4947 + r_run_k_17);
	assign w_sys_tmp4947 = 32'sh00000f3e;
	assign w_sys_tmp4951 = (w_sys_tmp4952 + r_run_k_17);
	assign w_sys_tmp4952 = 32'sh00000fbf;
	assign w_sys_tmp4956 = (w_sys_tmp4957 + r_run_k_17);
	assign w_sys_tmp4957 = 32'sh00001040;
	assign w_sys_tmp4961 = (w_sys_tmp4962 + r_run_k_17);
	assign w_sys_tmp4962 = 32'sh000010c1;
	assign w_sys_tmp4966 = (w_sys_tmp4967 + r_run_k_17);
	assign w_sys_tmp4967 = 32'sh00001142;
	assign w_sys_tmp4971 = (w_sys_tmp4972 + r_run_k_17);
	assign w_sys_tmp4972 = 32'sh000011c3;
	assign w_sys_tmp4976 = (w_sys_tmp4977 + r_run_k_17);
	assign w_sys_tmp4977 = 32'sh00001244;
	assign w_sys_tmp4981 = (w_sys_tmp4982 + r_run_k_17);
	assign w_sys_tmp4982 = 32'sh000012c5;
	assign w_sys_tmp4986 = (w_sys_tmp4987 + r_run_k_17);
	assign w_sys_tmp4987 = 32'sh00001346;
	assign w_sys_tmp4991 = (w_sys_tmp4992 + r_run_k_17);
	assign w_sys_tmp4992 = 32'sh000013c7;
	assign w_sys_tmp4996 = (w_sys_tmp4997 + r_run_k_17);
	assign w_sys_tmp4997 = 32'sh00001448;
	assign w_sys_tmp5001 = (w_sys_tmp5002 + r_run_k_17);
	assign w_sys_tmp5002 = 32'sh000014c9;
	assign w_sys_tmp5006 = (w_sys_tmp5007 + r_run_k_17);
	assign w_sys_tmp5007 = 32'sh0000154a;
	assign w_sys_tmp5011 = (w_sys_tmp5012 + r_run_k_17);
	assign w_sys_tmp5012 = 32'sh000015cb;
	assign w_sys_tmp5016 = (w_sys_tmp5017 + r_run_k_17);
	assign w_sys_tmp5017 = 32'sh0000164c;
	assign w_sys_tmp5021 = (w_sys_tmp5022 + r_run_k_17);
	assign w_sys_tmp5022 = 32'sh000016cd;
	assign w_sys_tmp5026 = (w_sys_tmp5027 + r_run_k_17);
	assign w_sys_tmp5027 = 32'sh0000174e;
	assign w_sys_tmp5031 = (w_sys_tmp5032 + r_run_k_17);
	assign w_sys_tmp5032 = 32'sh000017cf;
	assign w_sys_tmp5036 = (w_sys_tmp5037 + r_run_k_17);
	assign w_sys_tmp5037 = 32'sh00001850;
	assign w_sys_tmp5041 = (w_sys_tmp5042 + r_run_k_17);
	assign w_sys_tmp5042 = 32'sh000018d1;
	assign w_sys_tmp5046 = (w_sys_tmp5047 + r_run_k_17);
	assign w_sys_tmp5047 = 32'sh00001952;
	assign w_sys_tmp5051 = (w_sys_tmp5052 + r_run_k_17);
	assign w_sys_tmp5052 = 32'sh000019d3;
	assign w_sys_tmp5056 = (w_sys_tmp5057 + r_run_k_17);
	assign w_sys_tmp5057 = 32'sh00001a54;
	assign w_sys_tmp5061 = (w_sys_tmp5062 + r_run_k_17);
	assign w_sys_tmp5062 = 32'sh00001ad5;
	assign w_sys_tmp5066 = (w_sys_tmp5067 + r_run_k_17);
	assign w_sys_tmp5067 = 32'sh00001b56;
	assign w_sys_tmp5071 = (w_sys_tmp5072 + r_run_k_17);
	assign w_sys_tmp5072 = 32'sh00001bd7;
	assign w_sys_tmp5076 = (w_sys_tmp5077 + r_run_k_17);
	assign w_sys_tmp5077 = 32'sh00001c58;
	assign w_sys_tmp5081 = (w_sys_tmp5082 + r_run_k_17);
	assign w_sys_tmp5082 = 32'sh00001cd9;
	assign w_sys_tmp5086 = (w_sys_tmp5087 + r_run_k_17);
	assign w_sys_tmp5087 = 32'sh00001d5a;
	assign w_sys_tmp5091 = (w_sys_tmp5092 + r_run_k_17);
	assign w_sys_tmp5092 = 32'sh00001ddb;
	assign w_sys_tmp5096 = (w_sys_tmp5097 + r_run_k_17);
	assign w_sys_tmp5097 = 32'sh00001e5c;
	assign w_sys_tmp5101 = (w_sys_tmp5102 + r_run_k_17);
	assign w_sys_tmp5102 = 32'sh00001edd;
	assign w_sys_tmp5106 = (w_sys_tmp5107 + r_run_k_17);
	assign w_sys_tmp5107 = 32'sh00001f5e;
	assign w_sys_tmp5111 = (w_sys_tmp5112 + r_run_k_17);
	assign w_sys_tmp5112 = 32'sh00001fdf;
	assign w_sys_tmp5116 = (w_sys_tmp5117 + r_run_k_17);
	assign w_sys_tmp5117 = 32'sh00002060;
	assign w_sys_tmp5121 = (w_sys_tmp5122 + r_run_k_17);
	assign w_sys_tmp5122 = 32'sh000020e1;
	assign w_sys_tmp5126 = (w_sys_tmp5127 + r_run_k_17);
	assign w_sys_tmp5127 = 32'sh00002162;
	assign w_sys_tmp5131 = (w_sys_tmp5132 + r_run_k_17);
	assign w_sys_tmp5132 = 32'sh000021e3;
	assign w_sys_tmp5136 = (w_sys_tmp5137 + r_run_k_17);
	assign w_sys_tmp5137 = 32'sh00002264;
	assign w_sys_tmp5141 = (w_sys_tmp5142 + r_run_k_17);
	assign w_sys_tmp5142 = 32'sh000022e5;
	assign w_sys_tmp5146 = (w_sys_tmp5147 + r_run_k_17);
	assign w_sys_tmp5147 = 32'sh00002366;
	assign w_sys_tmp5151 = (w_sys_tmp5152 + r_run_k_17);
	assign w_sys_tmp5152 = 32'sh000023e7;
	assign w_sys_tmp5156 = (w_sys_tmp5157 + r_run_k_17);
	assign w_sys_tmp5157 = 32'sh00002468;
	assign w_sys_tmp5161 = (w_sys_tmp5162 + r_run_k_17);
	assign w_sys_tmp5162 = 32'sh000024e9;
	assign w_sys_tmp5166 = (w_sys_tmp5167 + r_run_k_17);
	assign w_sys_tmp5167 = 32'sh0000256a;
	assign w_sys_tmp5171 = (w_sys_tmp5172 + r_run_k_17);
	assign w_sys_tmp5172 = 32'sh000025eb;
	assign w_sys_tmp5176 = (w_sys_tmp5177 + r_run_k_17);
	assign w_sys_tmp5177 = 32'sh0000266c;
	assign w_sys_tmp5181 = (w_sys_tmp5182 + r_run_k_17);
	assign w_sys_tmp5182 = 32'sh000026ed;
	assign w_sys_tmp5186 = (w_sys_tmp5187 + r_run_k_17);
	assign w_sys_tmp5187 = 32'sh0000276e;
	assign w_sys_tmp5191 = (w_sys_tmp5192 + r_run_k_17);
	assign w_sys_tmp5192 = 32'sh000027ef;
	assign w_sys_tmp5196 = (w_sys_tmp5197 + r_run_k_17);
	assign w_sys_tmp5197 = 32'sh00002870;
	assign w_sys_tmp5201 = (w_sys_tmp5202 + r_run_k_17);
	assign w_sys_tmp5202 = 32'sh000028f1;
	assign w_sys_tmp5206 = (w_sys_tmp5207 + r_run_k_17);
	assign w_sys_tmp5207 = 32'sh00002972;
	assign w_sys_tmp5211 = (w_sys_tmp5212 + r_run_k_17);
	assign w_sys_tmp5212 = 32'sh000029f3;
	assign w_sys_tmp5216 = (w_sys_tmp5217 + r_run_k_17);
	assign w_sys_tmp5217 = 32'sh00002a74;
	assign w_sys_tmp5221 = (w_sys_tmp5222 + r_run_k_17);
	assign w_sys_tmp5222 = 32'sh00002af5;
	assign w_sys_tmp5226 = (w_sys_tmp5227 + r_run_k_17);
	assign w_sys_tmp5227 = 32'sh00002b76;
	assign w_sys_tmp5231 = (w_sys_tmp5232 + r_run_k_17);
	assign w_sys_tmp5232 = 32'sh00002bf7;
	assign w_sys_tmp5236 = (w_sys_tmp5237 + r_run_k_17);
	assign w_sys_tmp5237 = 32'sh00002c78;
	assign w_sys_tmp5241 = (w_sys_tmp5242 + r_run_k_17);
	assign w_sys_tmp5242 = 32'sh00002cf9;
	assign w_sys_tmp5246 = (w_sys_tmp5247 + r_run_k_17);
	assign w_sys_tmp5247 = 32'sh00002d7a;
	assign w_sys_tmp5251 = (w_sys_tmp5252 + r_run_k_17);
	assign w_sys_tmp5252 = 32'sh00002dfb;
	assign w_sys_tmp5256 = (w_sys_tmp5257 + r_run_k_17);
	assign w_sys_tmp5257 = 32'sh00002e7c;
	assign w_sys_tmp5261 = (w_sys_tmp5262 + r_run_k_17);
	assign w_sys_tmp5262 = 32'sh00002efd;
	assign w_sys_tmp5266 = (w_sys_tmp5267 + r_run_k_17);
	assign w_sys_tmp5267 = 32'sh00002f7e;
	assign w_sys_tmp5271 = (w_sys_tmp5272 + r_run_k_17);
	assign w_sys_tmp5272 = 32'sh00002fff;
	assign w_sys_tmp5276 = (w_sys_tmp5277 + r_run_k_17);
	assign w_sys_tmp5277 = 32'sh00003080;
	assign w_sys_tmp5281 = (w_sys_tmp5282 + r_run_k_17);
	assign w_sys_tmp5282 = 32'sh00003101;
	assign w_sys_tmp5286 = (w_sys_tmp5287 + r_run_k_17);
	assign w_sys_tmp5287 = 32'sh00003182;
	assign w_sys_tmp5291 = (w_sys_tmp5292 + r_run_k_17);
	assign w_sys_tmp5292 = 32'sh00003203;
	assign w_sys_tmp5296 = (w_sys_tmp5297 + r_run_k_17);
	assign w_sys_tmp5297 = 32'sh00003284;
	assign w_sys_tmp5301 = (w_sys_tmp5302 + r_run_k_17);
	assign w_sys_tmp5302 = 32'sh00003305;
	assign w_sys_tmp5306 = (w_sys_tmp5307 + r_run_k_17);
	assign w_sys_tmp5307 = 32'sh00003386;
	assign w_sys_tmp5311 = (w_sys_tmp5312 + r_run_k_17);
	assign w_sys_tmp5312 = 32'sh00003407;
	assign w_sys_tmp5316 = (w_sys_tmp5317 + r_run_k_17);
	assign w_sys_tmp5317 = 32'sh00003488;
	assign w_sys_tmp5321 = (w_sys_tmp5322 + r_run_k_17);
	assign w_sys_tmp5322 = 32'sh00003509;
	assign w_sys_tmp5326 = (w_sys_tmp5327 + r_run_k_17);
	assign w_sys_tmp5327 = 32'sh0000358a;
	assign w_sys_tmp5331 = (w_sys_tmp5332 + r_run_k_17);
	assign w_sys_tmp5332 = 32'sh0000360b;
	assign w_sys_tmp5336 = (w_sys_tmp5337 + r_run_k_17);
	assign w_sys_tmp5337 = 32'sh0000368c;
	assign w_sys_tmp5341 = (w_sys_tmp5342 + r_run_k_17);
	assign w_sys_tmp5342 = 32'sh0000370d;
	assign w_sys_tmp5346 = (w_sys_tmp5347 + r_run_k_17);
	assign w_sys_tmp5347 = 32'sh0000378e;
	assign w_sys_tmp5351 = (w_sys_tmp5352 + r_run_k_17);
	assign w_sys_tmp5352 = 32'sh0000380f;
	assign w_sys_tmp5356 = (w_sys_tmp5357 + r_run_k_17);
	assign w_sys_tmp5357 = 32'sh00003890;
	assign w_sys_tmp5361 = (w_sys_tmp5362 + r_run_k_17);
	assign w_sys_tmp5362 = 32'sh00003911;
	assign w_sys_tmp5366 = (w_sys_tmp5367 + r_run_k_17);
	assign w_sys_tmp5367 = 32'sh00003992;
	assign w_sys_tmp5371 = (w_sys_tmp5372 + r_run_k_17);
	assign w_sys_tmp5372 = 32'sh00003a13;
	assign w_sys_tmp5376 = (w_sys_tmp5377 + r_run_k_17);
	assign w_sys_tmp5377 = 32'sh00003a94;
	assign w_sys_tmp5381 = (w_sys_tmp5382 + r_run_k_17);
	assign w_sys_tmp5382 = 32'sh00003b15;
	assign w_sys_tmp5386 = (w_sys_tmp5387 + r_run_k_17);
	assign w_sys_tmp5387 = 32'sh00003b96;
	assign w_sys_tmp5391 = (w_sys_tmp5392 + r_run_k_17);
	assign w_sys_tmp5392 = 32'sh00003c17;
	assign w_sys_tmp5396 = (w_sys_tmp5397 + r_run_k_17);
	assign w_sys_tmp5397 = 32'sh00003c98;
	assign w_sys_tmp5401 = (w_sys_tmp5402 + r_run_k_17);
	assign w_sys_tmp5402 = 32'sh00003d19;
	assign w_sys_tmp5406 = (w_sys_tmp5407 + r_run_k_17);
	assign w_sys_tmp5407 = 32'sh00003d9a;
	assign w_sys_tmp5411 = (w_sys_tmp5412 + r_run_k_17);
	assign w_sys_tmp5412 = 32'sh00003e1b;
	assign w_sys_tmp5416 = (w_sys_tmp5417 + r_run_k_17);
	assign w_sys_tmp5417 = 32'sh00003e9c;
	assign w_sys_tmp5421 = (w_sys_tmp5422 + r_run_k_17);
	assign w_sys_tmp5422 = 32'sh00003f1d;
	assign w_sys_tmp5426 = (w_sys_tmp5427 + r_run_k_17);
	assign w_sys_tmp5427 = 32'sh00003f9e;
	assign w_sys_tmp5431 = (w_sys_tmp5432 + r_run_k_17);
	assign w_sys_tmp5432 = 32'sh0000401f;
	assign w_sys_tmp5436 = (w_sys_tmp5437 + r_run_k_17);
	assign w_sys_tmp5437 = 32'sh000040a0;
	assign w_sys_tmp5441 = (w_sys_tmp5442 + r_run_k_17);
	assign w_sys_tmp5442 = 32'sh00000142;
	assign w_sys_tmp5446 = (w_sys_tmp5447 + r_run_k_17);
	assign w_sys_tmp5447 = 32'sh000001c3;
	assign w_sys_tmp5451 = (w_sys_tmp5452 + r_run_k_17);
	assign w_sys_tmp5452 = 32'sh00000244;
	assign w_sys_tmp5456 = (w_sys_tmp5457 + r_run_k_17);
	assign w_sys_tmp5457 = 32'sh000002c5;
	assign w_sys_tmp5461 = (w_sys_tmp5462 + r_run_k_17);
	assign w_sys_tmp5462 = 32'sh00000346;
	assign w_sys_tmp5466 = (w_sys_tmp5467 + r_run_k_17);
	assign w_sys_tmp5467 = 32'sh000003c7;
	assign w_sys_tmp5471 = (w_sys_tmp5472 + r_run_k_17);
	assign w_sys_tmp5472 = 32'sh00000448;
	assign w_sys_tmp5476 = (w_sys_tmp5477 + r_run_k_17);
	assign w_sys_tmp5477 = 32'sh000004c9;
	assign w_sys_tmp5481 = (w_sys_tmp5482 + r_run_k_17);
	assign w_sys_tmp5482 = 32'sh0000054a;
	assign w_sys_tmp5486 = (w_sys_tmp5487 + r_run_k_17);
	assign w_sys_tmp5487 = 32'sh000005cb;
	assign w_sys_tmp5491 = (w_sys_tmp5492 + r_run_k_17);
	assign w_sys_tmp5492 = 32'sh0000064c;
	assign w_sys_tmp5496 = (w_sys_tmp5497 + r_run_k_17);
	assign w_sys_tmp5497 = 32'sh000006cd;
	assign w_sys_tmp5501 = (w_sys_tmp5502 + r_run_k_17);
	assign w_sys_tmp5502 = 32'sh0000074e;
	assign w_sys_tmp5506 = (w_sys_tmp5507 + r_run_k_17);
	assign w_sys_tmp5507 = 32'sh000007cf;
	assign w_sys_tmp5511 = (w_sys_tmp5512 + r_run_k_17);
	assign w_sys_tmp5512 = 32'sh00000850;
	assign w_sys_tmp5516 = (w_sys_tmp5517 + r_run_k_17);
	assign w_sys_tmp5517 = 32'sh000008d1;
	assign w_sys_tmp5521 = (w_sys_tmp5522 + r_run_k_17);
	assign w_sys_tmp5522 = 32'sh00000952;
	assign w_sys_tmp5526 = (w_sys_tmp5527 + r_run_k_17);
	assign w_sys_tmp5527 = 32'sh000009d3;
	assign w_sys_tmp5531 = (w_sys_tmp5532 + r_run_k_17);
	assign w_sys_tmp5532 = 32'sh00000a54;
	assign w_sys_tmp5536 = (w_sys_tmp5537 + r_run_k_17);
	assign w_sys_tmp5537 = 32'sh00000ad5;
	assign w_sys_tmp5541 = (w_sys_tmp5542 + r_run_k_17);
	assign w_sys_tmp5542 = 32'sh00000b56;
	assign w_sys_tmp5546 = (w_sys_tmp5547 + r_run_k_17);
	assign w_sys_tmp5547 = 32'sh00000bd7;
	assign w_sys_tmp5551 = (w_sys_tmp5552 + r_run_k_17);
	assign w_sys_tmp5552 = 32'sh00000c58;
	assign w_sys_tmp5556 = (w_sys_tmp5557 + r_run_k_17);
	assign w_sys_tmp5557 = 32'sh00000cd9;
	assign w_sys_tmp5561 = (w_sys_tmp5562 + r_run_k_17);
	assign w_sys_tmp5562 = 32'sh00000d5a;
	assign w_sys_tmp5566 = (w_sys_tmp5567 + r_run_k_17);
	assign w_sys_tmp5567 = 32'sh00000ddb;
	assign w_sys_tmp5571 = (w_sys_tmp5572 + r_run_k_17);
	assign w_sys_tmp5572 = 32'sh00000e5c;
	assign w_sys_tmp5576 = (w_sys_tmp5577 + r_run_k_17);
	assign w_sys_tmp5577 = 32'sh00000edd;
	assign w_sys_tmp5581 = (w_sys_tmp5582 + r_run_k_17);
	assign w_sys_tmp5582 = 32'sh00000f5e;
	assign w_sys_tmp5586 = (w_sys_tmp5587 + r_run_k_17);
	assign w_sys_tmp5587 = 32'sh00000fdf;
	assign w_sys_tmp5591 = (w_sys_tmp5592 + r_run_k_17);
	assign w_sys_tmp5592 = 32'sh00001060;
	assign w_sys_tmp5596 = (w_sys_tmp5597 + r_run_k_17);
	assign w_sys_tmp5597 = 32'sh000010e1;
	assign w_sys_tmp5601 = (w_sys_tmp5602 + r_run_k_17);
	assign w_sys_tmp5602 = 32'sh00001162;
	assign w_sys_tmp5606 = (w_sys_tmp5607 + r_run_k_17);
	assign w_sys_tmp5607 = 32'sh000011e3;
	assign w_sys_tmp5611 = (w_sys_tmp5612 + r_run_k_17);
	assign w_sys_tmp5612 = 32'sh00001264;
	assign w_sys_tmp5616 = (w_sys_tmp5617 + r_run_k_17);
	assign w_sys_tmp5617 = 32'sh000012e5;
	assign w_sys_tmp5621 = (w_sys_tmp5622 + r_run_k_17);
	assign w_sys_tmp5622 = 32'sh00001366;
	assign w_sys_tmp5626 = (w_sys_tmp5627 + r_run_k_17);
	assign w_sys_tmp5627 = 32'sh000013e7;
	assign w_sys_tmp5631 = (w_sys_tmp5632 + r_run_k_17);
	assign w_sys_tmp5632 = 32'sh00001468;
	assign w_sys_tmp5636 = (w_sys_tmp5637 + r_run_k_17);
	assign w_sys_tmp5637 = 32'sh000014e9;
	assign w_sys_tmp5641 = (w_sys_tmp5642 + r_run_k_17);
	assign w_sys_tmp5642 = 32'sh0000156a;
	assign w_sys_tmp5646 = (w_sys_tmp5647 + r_run_k_17);
	assign w_sys_tmp5647 = 32'sh000015eb;
	assign w_sys_tmp5651 = (w_sys_tmp5652 + r_run_k_17);
	assign w_sys_tmp5652 = 32'sh0000166c;
	assign w_sys_tmp5656 = (w_sys_tmp5657 + r_run_k_17);
	assign w_sys_tmp5657 = 32'sh000016ed;
	assign w_sys_tmp5661 = (w_sys_tmp5662 + r_run_k_17);
	assign w_sys_tmp5662 = 32'sh0000176e;
	assign w_sys_tmp5666 = (w_sys_tmp5667 + r_run_k_17);
	assign w_sys_tmp5667 = 32'sh000017ef;
	assign w_sys_tmp5671 = (w_sys_tmp5672 + r_run_k_17);
	assign w_sys_tmp5672 = 32'sh00001870;
	assign w_sys_tmp5676 = (w_sys_tmp5677 + r_run_k_17);
	assign w_sys_tmp5677 = 32'sh000018f1;
	assign w_sys_tmp5681 = (w_sys_tmp5682 + r_run_k_17);
	assign w_sys_tmp5682 = 32'sh00001972;
	assign w_sys_tmp5686 = (w_sys_tmp5687 + r_run_k_17);
	assign w_sys_tmp5687 = 32'sh000019f3;
	assign w_sys_tmp5691 = (w_sys_tmp5692 + r_run_k_17);
	assign w_sys_tmp5692 = 32'sh00001a74;
	assign w_sys_tmp5696 = (w_sys_tmp5697 + r_run_k_17);
	assign w_sys_tmp5697 = 32'sh00001af5;
	assign w_sys_tmp5701 = (w_sys_tmp5702 + r_run_k_17);
	assign w_sys_tmp5702 = 32'sh00001b76;
	assign w_sys_tmp5706 = (w_sys_tmp5707 + r_run_k_17);
	assign w_sys_tmp5707 = 32'sh00001bf7;
	assign w_sys_tmp5711 = (w_sys_tmp5712 + r_run_k_17);
	assign w_sys_tmp5712 = 32'sh00001c78;
	assign w_sys_tmp5716 = (w_sys_tmp5717 + r_run_k_17);
	assign w_sys_tmp5717 = 32'sh00001cf9;
	assign w_sys_tmp5721 = (w_sys_tmp5722 + r_run_k_17);
	assign w_sys_tmp5722 = 32'sh00001d7a;
	assign w_sys_tmp5726 = (w_sys_tmp5727 + r_run_k_17);
	assign w_sys_tmp5727 = 32'sh00001dfb;
	assign w_sys_tmp5731 = (w_sys_tmp5732 + r_run_k_17);
	assign w_sys_tmp5732 = 32'sh00001e7c;
	assign w_sys_tmp5736 = (w_sys_tmp5737 + r_run_k_17);
	assign w_sys_tmp5737 = 32'sh00001efd;
	assign w_sys_tmp5741 = (w_sys_tmp5742 + r_run_k_17);
	assign w_sys_tmp5742 = 32'sh00001f7e;
	assign w_sys_tmp5746 = (w_sys_tmp5747 + r_run_k_17);
	assign w_sys_tmp5747 = 32'sh00001fff;
	assign w_sys_tmp5751 = (w_sys_tmp5752 + r_run_k_17);
	assign w_sys_tmp5752 = 32'sh00002080;
	assign w_sys_tmp5756 = (w_sys_tmp5757 + r_run_k_17);
	assign w_sys_tmp5757 = 32'sh00002101;
	assign w_sys_tmp5761 = (w_sys_tmp5762 + r_run_k_17);
	assign w_sys_tmp5762 = 32'sh00002182;
	assign w_sys_tmp5766 = (w_sys_tmp5767 + r_run_k_17);
	assign w_sys_tmp5767 = 32'sh00002203;
	assign w_sys_tmp5771 = (w_sys_tmp5772 + r_run_k_17);
	assign w_sys_tmp5772 = 32'sh00002284;
	assign w_sys_tmp5776 = (w_sys_tmp5777 + r_run_k_17);
	assign w_sys_tmp5777 = 32'sh00002305;
	assign w_sys_tmp5781 = (w_sys_tmp5782 + r_run_k_17);
	assign w_sys_tmp5782 = 32'sh00002386;
	assign w_sys_tmp5786 = (w_sys_tmp5787 + r_run_k_17);
	assign w_sys_tmp5787 = 32'sh00002407;
	assign w_sys_tmp5791 = (w_sys_tmp5792 + r_run_k_17);
	assign w_sys_tmp5792 = 32'sh00002488;
	assign w_sys_tmp5796 = (w_sys_tmp5797 + r_run_k_17);
	assign w_sys_tmp5797 = 32'sh00002509;
	assign w_sys_tmp5801 = (w_sys_tmp5802 + r_run_k_17);
	assign w_sys_tmp5802 = 32'sh0000258a;
	assign w_sys_tmp5806 = (w_sys_tmp5807 + r_run_k_17);
	assign w_sys_tmp5807 = 32'sh0000260b;
	assign w_sys_tmp5811 = (w_sys_tmp5812 + r_run_k_17);
	assign w_sys_tmp5812 = 32'sh0000268c;
	assign w_sys_tmp5816 = (w_sys_tmp5817 + r_run_k_17);
	assign w_sys_tmp5817 = 32'sh0000270d;
	assign w_sys_tmp5821 = (w_sys_tmp5822 + r_run_k_17);
	assign w_sys_tmp5822 = 32'sh0000278e;
	assign w_sys_tmp5826 = (w_sys_tmp5827 + r_run_k_17);
	assign w_sys_tmp5827 = 32'sh0000280f;
	assign w_sys_tmp5831 = (w_sys_tmp5832 + r_run_k_17);
	assign w_sys_tmp5832 = 32'sh00002890;
	assign w_sys_tmp5836 = (w_sys_tmp5837 + r_run_k_17);
	assign w_sys_tmp5837 = 32'sh00002911;
	assign w_sys_tmp5841 = (w_sys_tmp5842 + r_run_k_17);
	assign w_sys_tmp5842 = 32'sh00002992;
	assign w_sys_tmp5846 = (w_sys_tmp5847 + r_run_k_17);
	assign w_sys_tmp5847 = 32'sh00002a13;
	assign w_sys_tmp5851 = (w_sys_tmp5852 + r_run_k_17);
	assign w_sys_tmp5852 = 32'sh00002a94;
	assign w_sys_tmp5856 = (w_sys_tmp5857 + r_run_k_17);
	assign w_sys_tmp5857 = 32'sh00002b15;
	assign w_sys_tmp5861 = (w_sys_tmp5862 + r_run_k_17);
	assign w_sys_tmp5862 = 32'sh00002b96;
	assign w_sys_tmp5866 = (w_sys_tmp5867 + r_run_k_17);
	assign w_sys_tmp5867 = 32'sh00002c17;
	assign w_sys_tmp5871 = (w_sys_tmp5872 + r_run_k_17);
	assign w_sys_tmp5872 = 32'sh00002c98;
	assign w_sys_tmp5876 = (w_sys_tmp5877 + r_run_k_17);
	assign w_sys_tmp5877 = 32'sh00002d19;
	assign w_sys_tmp5881 = (w_sys_tmp5882 + r_run_k_17);
	assign w_sys_tmp5882 = 32'sh00002d9a;
	assign w_sys_tmp5886 = (w_sys_tmp5887 + r_run_k_17);
	assign w_sys_tmp5887 = 32'sh00002e1b;
	assign w_sys_tmp5891 = (w_sys_tmp5892 + r_run_k_17);
	assign w_sys_tmp5892 = 32'sh00002e9c;
	assign w_sys_tmp5896 = (w_sys_tmp5897 + r_run_k_17);
	assign w_sys_tmp5897 = 32'sh00002f1d;
	assign w_sys_tmp5901 = (w_sys_tmp5902 + r_run_k_17);
	assign w_sys_tmp5902 = 32'sh00002f9e;
	assign w_sys_tmp5906 = (w_sys_tmp5907 + r_run_k_17);
	assign w_sys_tmp5907 = 32'sh0000301f;
	assign w_sys_tmp5911 = (w_sys_tmp5912 + r_run_k_17);
	assign w_sys_tmp5912 = 32'sh000030a0;
	assign w_sys_tmp5916 = (w_sys_tmp5917 + r_run_k_17);
	assign w_sys_tmp5917 = 32'sh00003121;
	assign w_sys_tmp5921 = (w_sys_tmp5922 + r_run_k_17);
	assign w_sys_tmp5922 = 32'sh000031a2;
	assign w_sys_tmp5926 = (w_sys_tmp5927 + r_run_k_17);
	assign w_sys_tmp5927 = 32'sh00003223;
	assign w_sys_tmp5931 = (w_sys_tmp5932 + r_run_k_17);
	assign w_sys_tmp5932 = 32'sh000032a4;
	assign w_sys_tmp5936 = (w_sys_tmp5937 + r_run_k_17);
	assign w_sys_tmp5937 = 32'sh00003325;
	assign w_sys_tmp5941 = (w_sys_tmp5942 + r_run_k_17);
	assign w_sys_tmp5942 = 32'sh000033a6;
	assign w_sys_tmp5946 = (w_sys_tmp5947 + r_run_k_17);
	assign w_sys_tmp5947 = 32'sh00003427;
	assign w_sys_tmp5951 = (w_sys_tmp5952 + r_run_k_17);
	assign w_sys_tmp5952 = 32'sh000034a8;
	assign w_sys_tmp5956 = (w_sys_tmp5957 + r_run_k_17);
	assign w_sys_tmp5957 = 32'sh00003529;
	assign w_sys_tmp5961 = (w_sys_tmp5962 + r_run_k_17);
	assign w_sys_tmp5962 = 32'sh000035aa;
	assign w_sys_tmp5966 = (w_sys_tmp5967 + r_run_k_17);
	assign w_sys_tmp5967 = 32'sh0000362b;
	assign w_sys_tmp5971 = (w_sys_tmp5972 + r_run_k_17);
	assign w_sys_tmp5972 = 32'sh000036ac;
	assign w_sys_tmp5976 = (w_sys_tmp5977 + r_run_k_17);
	assign w_sys_tmp5977 = 32'sh0000372d;
	assign w_sys_tmp5981 = (w_sys_tmp5982 + r_run_k_17);
	assign w_sys_tmp5982 = 32'sh000037ae;
	assign w_sys_tmp5986 = (w_sys_tmp5987 + r_run_k_17);
	assign w_sys_tmp5987 = 32'sh0000382f;
	assign w_sys_tmp5991 = (w_sys_tmp5992 + r_run_k_17);
	assign w_sys_tmp5992 = 32'sh000038b0;
	assign w_sys_tmp5996 = (w_sys_tmp5997 + r_run_k_17);
	assign w_sys_tmp5997 = 32'sh00003931;
	assign w_sys_tmp6001 = (w_sys_tmp6002 + r_run_k_17);
	assign w_sys_tmp6002 = 32'sh000039b2;
	assign w_sys_tmp6006 = (w_sys_tmp6007 + r_run_k_17);
	assign w_sys_tmp6007 = 32'sh00003a33;
	assign w_sys_tmp6011 = (w_sys_tmp6012 + r_run_k_17);
	assign w_sys_tmp6012 = 32'sh00003ab4;
	assign w_sys_tmp6016 = (w_sys_tmp6017 + r_run_k_17);
	assign w_sys_tmp6017 = 32'sh00003b35;
	assign w_sys_tmp6021 = (w_sys_tmp6022 + r_run_k_17);
	assign w_sys_tmp6022 = 32'sh00003bb6;
	assign w_sys_tmp6026 = (w_sys_tmp6027 + r_run_k_17);
	assign w_sys_tmp6027 = 32'sh00003c37;
	assign w_sys_tmp6031 = (w_sys_tmp6032 + r_run_k_17);
	assign w_sys_tmp6032 = 32'sh00003cb8;
	assign w_sys_tmp6036 = (w_sys_tmp6037 + r_run_k_17);
	assign w_sys_tmp6037 = 32'sh00003d39;
	assign w_sys_tmp6041 = (w_sys_tmp6042 + r_run_k_17);
	assign w_sys_tmp6042 = 32'sh00003dba;
	assign w_sys_tmp6046 = (w_sys_tmp6047 + r_run_k_17);
	assign w_sys_tmp6047 = 32'sh00003e3b;
	assign w_sys_tmp6051 = (w_sys_tmp6052 + r_run_k_17);
	assign w_sys_tmp6052 = 32'sh00003ebc;
	assign w_sys_tmp6056 = (w_sys_tmp6057 + r_run_k_17);
	assign w_sys_tmp6057 = 32'sh00003f3d;
	assign w_sys_tmp6061 = (w_sys_tmp6062 + r_run_k_17);
	assign w_sys_tmp6062 = 32'sh00003fbe;
	assign w_sys_tmp6066 = (w_sys_tmp6067 + r_run_k_17);
	assign w_sys_tmp6067 = 32'sh0000403f;
	assign w_sys_tmp6071 = (w_sys_tmp6072 + r_run_k_17);
	assign w_sys_tmp6072 = 32'sh000040c0;
	assign w_sys_tmp6075 = (r_run_k_17 + w_sys_intOne);


	sub09
		sub09_inst(
			.i_fld_result_1_addr_0 (w_sub09_result_addr),
			.i_fld_result_1_datain_0 (w_sub09_result_datain),
			.o_fld_result_1_dataout_0 (w_sub09_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub09_result_r_w),
			.i_fld_u_0_addr_0 (w_sub09_u_addr),
			.i_fld_u_0_datain_0 (w_sub09_u_datain),
			.o_fld_u_0_dataout_0 (w_sub09_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub09_u_r_w),
			.o_run_busy (w_sub09_run_busy),
			.i_run_req (r_sub09_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub08
		sub08_inst(
			.i_fld_result_1_addr_0 (w_sub08_result_addr),
			.i_fld_result_1_datain_0 (w_sub08_result_datain),
			.o_fld_result_1_dataout_0 (w_sub08_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub08_result_r_w),
			.i_fld_u_0_addr_0 (w_sub08_u_addr),
			.i_fld_u_0_datain_0 (w_sub08_u_datain),
			.o_fld_u_0_dataout_0 (w_sub08_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub08_u_r_w),
			.o_run_busy (w_sub08_run_busy),
			.i_run_req (r_sub08_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub12
		sub12_inst(
			.i_fld_result_1_addr_0 (w_sub12_result_addr),
			.i_fld_result_1_datain_0 (w_sub12_result_datain),
			.o_fld_result_1_dataout_0 (w_sub12_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub12_result_r_w),
			.i_fld_u_0_addr_0 (w_sub12_u_addr),
			.i_fld_u_0_datain_0 (w_sub12_u_datain),
			.o_fld_u_0_dataout_0 (w_sub12_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub12_u_r_w),
			.o_run_busy (w_sub12_run_busy),
			.i_run_req (r_sub12_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub03
		sub03_inst(
			.i_fld_result_1_addr_0 (w_sub03_result_addr),
			.i_fld_result_1_datain_0 (w_sub03_result_datain),
			.o_fld_result_1_dataout_0 (w_sub03_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub03_result_r_w),
			.i_fld_u_0_addr_0 (w_sub03_u_addr),
			.i_fld_u_0_datain_0 (w_sub03_u_datain),
			.o_fld_u_0_dataout_0 (w_sub03_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub03_u_r_w),
			.o_run_busy (w_sub03_run_busy),
			.i_run_req (r_sub03_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub02
		sub02_inst(
			.i_fld_result_1_addr_0 (w_sub02_result_addr),
			.i_fld_result_1_datain_0 (w_sub02_result_datain),
			.o_fld_result_1_dataout_0 (w_sub02_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub02_result_r_w),
			.i_fld_u_0_addr_0 (w_sub02_u_addr),
			.i_fld_u_0_datain_0 (w_sub02_u_datain),
			.o_fld_u_0_dataout_0 (w_sub02_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub02_u_r_w),
			.o_run_busy (w_sub02_run_busy),
			.i_run_req (r_sub02_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub11
		sub11_inst(
			.i_fld_result_1_addr_0 (w_sub11_result_addr),
			.i_fld_result_1_datain_0 (w_sub11_result_datain),
			.o_fld_result_1_dataout_0 (w_sub11_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub11_result_r_w),
			.i_fld_u_0_addr_0 (w_sub11_u_addr),
			.i_fld_u_0_datain_0 (w_sub11_u_datain),
			.o_fld_u_0_dataout_0 (w_sub11_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub11_u_r_w),
			.o_run_busy (w_sub11_run_busy),
			.i_run_req (r_sub11_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub14
		sub14_inst(
			.i_fld_result_1_addr_0 (w_sub14_result_addr),
			.i_fld_result_1_datain_0 (w_sub14_result_datain),
			.o_fld_result_1_dataout_0 (w_sub14_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub14_result_r_w),
			.i_fld_u_0_addr_0 (w_sub14_u_addr),
			.i_fld_u_0_datain_0 (w_sub14_u_datain),
			.o_fld_u_0_dataout_0 (w_sub14_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub14_u_r_w),
			.o_run_busy (w_sub14_run_busy),
			.i_run_req (r_sub14_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub01
		sub01_inst(
			.i_fld_result_1_addr_0 (w_sub01_result_addr),
			.i_fld_result_1_datain_0 (w_sub01_result_datain),
			.o_fld_result_1_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub01_result_r_w),
			.i_fld_u_0_addr_0 (w_sub01_u_addr),
			.i_fld_u_0_datain_0 (w_sub01_u_datain),
			.o_fld_u_0_dataout_0 (w_sub01_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub01_u_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub13
		sub13_inst(
			.i_fld_result_1_addr_0 (w_sub13_result_addr),
			.i_fld_result_1_datain_0 (w_sub13_result_datain),
			.o_fld_result_1_dataout_0 (w_sub13_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub13_result_r_w),
			.i_fld_u_0_addr_0 (w_sub13_u_addr),
			.i_fld_u_0_datain_0 (w_sub13_u_datain),
			.o_fld_u_0_dataout_0 (w_sub13_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub13_u_r_w),
			.o_run_busy (w_sub13_run_busy),
			.i_run_req (r_sub13_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub00
		sub00_inst(
			.i_fld_result_1_addr_0 (w_sub00_result_addr),
			.i_fld_result_1_datain_0 (w_sub00_result_datain),
			.o_fld_result_1_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub00_result_r_w),
			.i_fld_u_0_addr_0 (w_sub00_u_addr),
			.i_fld_u_0_datain_0 (w_sub00_u_datain),
			.o_fld_u_0_dataout_0 (w_sub00_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub00_u_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub07
		sub07_inst(
			.i_fld_result_1_addr_0 (w_sub07_result_addr),
			.i_fld_result_1_datain_0 (w_sub07_result_datain),
			.o_fld_result_1_dataout_0 (w_sub07_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub07_result_r_w),
			.i_fld_u_0_addr_0 (w_sub07_u_addr),
			.i_fld_u_0_datain_0 (w_sub07_u_datain),
			.o_fld_u_0_dataout_0 (w_sub07_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub07_u_r_w),
			.o_run_busy (w_sub07_run_busy),
			.i_run_req (r_sub07_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub06
		sub06_inst(
			.i_fld_result_1_addr_0 (w_sub06_result_addr),
			.i_fld_result_1_datain_0 (w_sub06_result_datain),
			.o_fld_result_1_dataout_0 (w_sub06_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub06_result_r_w),
			.i_fld_u_0_addr_0 (w_sub06_u_addr),
			.i_fld_u_0_datain_0 (w_sub06_u_datain),
			.o_fld_u_0_dataout_0 (w_sub06_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub06_u_r_w),
			.o_run_busy (w_sub06_run_busy),
			.i_run_req (r_sub06_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub15
		sub15_inst(
			.i_fld_result_1_addr_0 (w_sub15_result_addr),
			.i_fld_result_1_datain_0 (w_sub15_result_datain),
			.o_fld_result_1_dataout_0 (w_sub15_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub15_result_r_w),
			.i_fld_u_0_addr_0 (w_sub15_u_addr),
			.i_fld_u_0_datain_0 (w_sub15_u_datain),
			.o_fld_u_0_dataout_0 (w_sub15_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub15_u_r_w),
			.o_run_busy (w_sub15_run_busy),
			.i_run_req (r_sub15_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub05
		sub05_inst(
			.i_fld_result_1_addr_0 (w_sub05_result_addr),
			.i_fld_result_1_datain_0 (w_sub05_result_datain),
			.o_fld_result_1_dataout_0 (w_sub05_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub05_result_r_w),
			.i_fld_u_0_addr_0 (w_sub05_u_addr),
			.i_fld_u_0_datain_0 (w_sub05_u_datain),
			.o_fld_u_0_dataout_0 (w_sub05_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub05_u_r_w),
			.o_run_busy (w_sub05_run_busy),
			.i_run_req (r_sub05_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub04
		sub04_inst(
			.i_fld_result_1_addr_0 (w_sub04_result_addr),
			.i_fld_result_1_datain_0 (w_sub04_result_datain),
			.o_fld_result_1_dataout_0 (w_sub04_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub04_result_r_w),
			.i_fld_u_0_addr_0 (w_sub04_u_addr),
			.i_fld_u_0_datain_0 (w_sub04_u_datain),
			.o_fld_u_0_dataout_0 (w_sub04_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub04_u_r_w),
			.o_run_busy (w_sub04_run_busy),
			.i_run_req (r_sub04_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub10
		sub10_inst(
			.i_fld_result_1_addr_0 (w_sub10_result_addr),
			.i_fld_result_1_datain_0 (w_sub10_result_datain),
			.o_fld_result_1_dataout_0 (w_sub10_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub10_result_r_w),
			.i_fld_u_0_addr_0 (w_sub10_u_addr),
			.i_fld_u_0_datain_0 (w_sub10_u_datain),
			.o_fld_u_0_dataout_0 (w_sub10_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub10_u_r_w),
			.o_run_busy (w_sub10_run_busy),
			.i_run_req (r_sub10_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_u_0(
			.clk (clock),
			.ce_0 (w_fld_u_0_ce_0),
			.addr_0 (w_fld_u_0_addr_0),
			.datain_0 (w_fld_u_0_datain_0),
			.dataout_0 (w_fld_u_0_dataout_0),
			.r_w_0 (w_fld_u_0_r_w_0),
			.ce_1 (w_fld_u_0_ce_1),
			.addr_1 (r_fld_u_0_addr_1),
			.datain_1 (r_fld_u_0_datain_1),
			.dataout_1 (w_fld_u_0_dataout_1),
			.r_w_1 (r_fld_u_0_r_w_1)
		);

	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h35: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 6'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_phase <= 6'h2;
						end

						6'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'h4;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3) ? 6'h9 : 6'hf);

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'ha;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6) ? 6'hd : 6'h6);

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_run_phase <= 6'ha;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'h10;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp51) ? 6'h14 : 6'h35);

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'h10;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'h15;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp54) ? 6'h18 : 6'h1a);

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sys_run_phase <= 6'h15;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'h1b;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp211) ? 6'h1e : 6'h20);

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h88)) begin
										r_sys_run_phase <= 6'h1b;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'h21;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1027) ? 6'h24 : 6'h25);

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h196)) begin
										r_sys_run_phase <= 6'h21;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h10: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_phase <= 6'h27;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_phase <= 6'h29;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'h2a;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3463) ? 6'h2d : 6'h2f);

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h80)) begin
										r_sys_run_phase <= 6'h2a;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 6'h30;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4135) ? 6'h33 : 6'h11);

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h17e)) begin
										r_sys_run_phase <= 6'h30;

									end
								end

							endcase
						end

						6'h35: begin
							r_sys_run_phase <= 6'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 5'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h88)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h196)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h80)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h17e)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 9'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h5)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1a)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h88)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h87)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h196)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h195)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub00_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub01_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub02_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub03_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub04_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub05_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub06_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub07_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub08_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub09_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub10_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub11_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub12_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub13_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub14_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub15_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h80)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h7f)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h17d)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==9'h17e)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						6'h35: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp10[14:0] );

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3) || (r_sys_run_step==9'h7) || (r_sys_run_step==9'hb) || (r_sys_run_step==9'hf) || (r_sys_run_step==9'h13) || (r_sys_run_step==9'h17) || (r_sys_run_step==9'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp71[14:0] );

									end
									else
									if((r_sys_run_step==9'h1) || (r_sys_run_step==9'h5) || (r_sys_run_step==9'h9) || (r_sys_run_step==9'hd) || (r_sys_run_step==9'h11) || (r_sys_run_step==9'h15) || (r_sys_run_step==9'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp62[14:0] );

									end
									else
									if((r_sys_run_step==9'h0) || (r_sys_run_step==9'h4) || (r_sys_run_step==9'h8) || (r_sys_run_step==9'hc) || (r_sys_run_step==9'h10) || (r_sys_run_step==9'h14) || (r_sys_run_step==9'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp58[14:0] );

									end
									else
									if((r_sys_run_step==9'h2) || (r_sys_run_step==9'h6) || (r_sys_run_step==9'ha) || (r_sys_run_step==9'he) || (r_sys_run_step==9'h12) || (r_sys_run_step==9'h16) || (r_sys_run_step==9'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp66[14:0] );

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp870[14:0] );

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp672[14:0] );

									end
									else
									if((r_sys_run_step==9'h7b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp954[14:0] );

									end
									else
									if((r_sys_run_step==9'h71)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp894[14:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp390[14:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp258[14:0] );

									end
									else
									if((r_sys_run_step==9'h2e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp492[14:0] );

									end
									else
									if((r_sys_run_step==9'h6a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp852[14:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp294[14:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp306[14:0] );

									end
									else
									if((r_sys_run_step==9'h3e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp588[14:0] );

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp708[14:0] );

									end
									else
									if((r_sys_run_step==9'h6f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp882[14:0] );

									end
									else
									if((r_sys_run_step==9'h6e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp876[14:0] );

									end
									else
									if((r_sys_run_step==9'h2d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp486[14:0] );

									end
									else
									if((r_sys_run_step==9'h68)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp840[14:0] );

									end
									else
									if((r_sys_run_step==9'h42) || (r_sys_run_step==9'h44)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp612[14:0] );

									end
									else
									if((r_sys_run_step==9'h62)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp804[14:0] );

									end
									else
									if((r_sys_run_step==9'h28)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp456[14:0] );

									end
									else
									if((r_sys_run_step==9'h5c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp768[14:0] );

									end
									else
									if((r_sys_run_step==9'h81)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp990[14:0] );

									end
									else
									if((r_sys_run_step==9'h3a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp564[14:0] );

									end
									else
									if((r_sys_run_step==9'h76)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp924[14:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp354[14:0] );

									end
									else
									if((r_sys_run_step==9'h41) || (r_sys_run_step==9'h43)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp606[14:0] );

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp642[14:0] );

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp684[14:0] );

									end
									else
									if((r_sys_run_step==9'h50)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp696[14:0] );

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp498[14:0] );

									end
									else
									if((r_sys_run_step==9'h30)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp504[14:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp366[14:0] );

									end
									else
									if((r_sys_run_step==9'h33)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp522[14:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp252[14:0] );

									end
									else
									if((r_sys_run_step==9'h40)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp600[14:0] );

									end
									else
									if((r_sys_run_step==9'h63) || (r_sys_run_step==9'h65)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp810[14:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp216[14:0] );

									end
									else
									if((r_sys_run_step==9'h80)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp984[14:0] );

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp432[14:0] );

									end
									else
									if((r_sys_run_step==9'h79)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp942[14:0] );

									end
									else
									if((r_sys_run_step==9'h84)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1008[14:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp372[14:0] );

									end
									else
									if((r_sys_run_step==9'h31)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp510[14:0] );

									end
									else
									if((r_sys_run_step==9'h67)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp834[14:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp330[14:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp282[14:0] );

									end
									else
									if((r_sys_run_step==9'h85)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1014[14:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp384[14:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp336[14:0] );

									end
									else
									if((r_sys_run_step==9'h35)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp534[14:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp318[14:0] );

									end
									else
									if((r_sys_run_step==9'h77)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp930[14:0] );

									end
									else
									if((r_sys_run_step==9'h32)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp516[14:0] );

									end
									else
									if((r_sys_run_step==9'h5f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp786[14:0] );

									end
									else
									if((r_sys_run_step==9'h7c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp960[14:0] );

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp666[14:0] );

									end
									else
									if((r_sys_run_step==9'h6b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp858[14:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp300[14:0] );

									end
									else
									if((r_sys_run_step==9'h2c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp480[14:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp240[14:0] );

									end
									else
									if((r_sys_run_step==9'h29)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp462[14:0] );

									end
									else
									if((r_sys_run_step==9'h5e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp780[14:0] );

									end
									else
									if((r_sys_run_step==9'h56)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp732[14:0] );

									end
									else
									if((r_sys_run_step==9'h45)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp630[14:0] );

									end
									else
									if((r_sys_run_step==9'h5b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp762[14:0] );

									end
									else
									if((r_sys_run_step==9'h36)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp540[14:0] );

									end
									else
									if((r_sys_run_step==9'h4a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp660[14:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp270[14:0] );

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp558[14:0] );

									end
									else
									if((r_sys_run_step==9'h2a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp468[14:0] );

									end
									else
									if((r_sys_run_step==9'h61)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp798[14:0] );

									end
									else
									if((r_sys_run_step==9'h58)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp744[14:0] );

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp582[14:0] );

									end
									else
									if((r_sys_run_step==9'h59)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp750[14:0] );

									end
									else
									if((r_sys_run_step==9'h27)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp450[14:0] );

									end
									else
									if((r_sys_run_step==9'h7e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp972[14:0] );

									end
									else
									if((r_sys_run_step==9'h46)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp636[14:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp264[14:0] );

									end
									else
									if((r_sys_run_step==9'h5a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp756[14:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp228[14:0] );

									end
									else
									if((r_sys_run_step==9'h57)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp738[14:0] );

									end
									else
									if((r_sys_run_step==9'h49)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp654[14:0] );

									end
									else
									if((r_sys_run_step==9'h60)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp792[14:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp378[14:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp312[14:0] );

									end
									else
									if((r_sys_run_step==9'h53)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp714[14:0] );

									end
									else
									if((r_sys_run_step==9'h48)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp648[14:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp276[14:0] );

									end
									else
									if((r_sys_run_step==9'h51)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp702[14:0] );

									end
									else
									if((r_sys_run_step==9'h75)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp918[14:0] );

									end
									else
									if((r_sys_run_step==9'h83)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1002[14:0] );

									end
									else
									if((r_sys_run_step==9'h38)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp552[14:0] );

									end
									else
									if((r_sys_run_step==9'h7f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp978[14:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp396[14:0] );

									end
									else
									if((r_sys_run_step==9'h74)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp912[14:0] );

									end
									else
									if((r_sys_run_step==9'h4f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp690[14:0] );

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp576[14:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp222[14:0] );

									end
									else
									if((r_sys_run_step==9'h72)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp900[14:0] );

									end
									else
									if((r_sys_run_step==9'h64) || (r_sys_run_step==9'h66)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp816[14:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp234[14:0] );

									end
									else
									if((r_sys_run_step==9'h82)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp996[14:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp324[14:0] );

									end
									else
									if((r_sys_run_step==9'h26)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp444[14:0] );

									end
									else
									if((r_sys_run_step==9'h37)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp546[14:0] );

									end
									else
									if((r_sys_run_step==9'h34)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp528[14:0] );

									end
									else
									if((r_sys_run_step==9'h4d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp678[14:0] );

									end
									else
									if((r_sys_run_step==9'h6c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp864[14:0] );

									end
									else
									if((r_sys_run_step==9'h70)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp888[14:0] );

									end
									else
									if((r_sys_run_step==9'h1f) || (r_sys_run_step==9'h21)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp402[14:0] );

									end
									else
									if((r_sys_run_step==9'h5d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp774[14:0] );

									end
									else
									if((r_sys_run_step==9'h23)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp426[14:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp360[14:0] );

									end
									else
									if((r_sys_run_step==9'h73)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp906[14:0] );

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp570[14:0] );

									end
									else
									if((r_sys_run_step==9'h78)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp936[14:0] );

									end
									else
									if((r_sys_run_step==9'h55)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp726[14:0] );

									end
									else
									if((r_sys_run_step==9'h86)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1020[14:0] );

									end
									else
									if((r_sys_run_step==9'h69)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp846[14:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp348[14:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp246[14:0] );

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp720[14:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp342[14:0] );

									end
									else
									if((r_sys_run_step==9'h20) || (r_sys_run_step==9'h22)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp408[14:0] );

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp438[14:0] );

									end
									else
									if((r_sys_run_step==9'h7d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp966[14:0] );

									end
									else
									if((r_sys_run_step==9'h2b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp474[14:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp288[14:0] );

									end
									else
									if((r_sys_run_step==9'h7a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp948[14:0] );

									end
									else
									if((r_sys_run_step==9'h3f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp594[14:0] );

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h28)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1272[14:0] );

									end
									else
									if((r_sys_run_step==9'h26)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1260[14:0] );

									end
									else
									if((r_sys_run_step==9'hfe)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2556[14:0] );

									end
									else
									if((r_sys_run_step==9'h87)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1842[14:0] );

									end
									else
									if((r_sys_run_step==9'h2d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1302[14:0] );

									end
									else
									if((r_sys_run_step==9'h94)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1920[14:0] );

									end
									else
									if((r_sys_run_step==9'he2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2388[14:0] );

									end
									else
									if((r_sys_run_step==9'h12e) || (r_sys_run_step==9'h130)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2844[14:0] );

									end
									else
									if((r_sys_run_step==9'h33)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1338[14:0] );

									end
									else
									if((r_sys_run_step==9'h16d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3222[14:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1110[14:0] );

									end
									else
									if((r_sys_run_step==9'h16e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3228[14:0] );

									end
									else
									if((r_sys_run_step==9'he9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2430[14:0] );

									end
									else
									if((r_sys_run_step==9'h101)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2574[14:0] );

									end
									else
									if((r_sys_run_step==9'h14e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3036[14:0] );

									end
									else
									if((r_sys_run_step==9'hc7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2226[14:0] );

									end
									else
									if((r_sys_run_step==9'h84)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1824[14:0] );

									end
									else
									if((r_sys_run_step==9'h11f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2754[14:0] );

									end
									else
									if((r_sys_run_step==9'h180)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3336[14:0] );

									end
									else
									if((r_sys_run_step==9'h134)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2880[14:0] );

									end
									else
									if((r_sys_run_step==9'h15f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3138[14:0] );

									end
									else
									if((r_sys_run_step==9'h112)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2676[14:0] );

									end
									else
									if((r_sys_run_step==9'h164)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3168[14:0] );

									end
									else
									if((r_sys_run_step==9'h7f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1794[14:0] );

									end
									else
									if((r_sys_run_step==9'h40)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1416[14:0] );

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1374[14:0] );

									end
									else
									if((r_sys_run_step==9'hd4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2304[14:0] );

									end
									else
									if((r_sys_run_step==9'hcc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2256[14:0] );

									end
									else
									if((r_sys_run_step==9'h167)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3186[14:0] );

									end
									else
									if((r_sys_run_step==9'h132)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2868[14:0] );

									end
									else
									if((r_sys_run_step==9'h12c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2832[14:0] );

									end
									else
									if((r_sys_run_step==9'hd1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2286[14:0] );

									end
									else
									if((r_sys_run_step==9'h16a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3204[14:0] );

									end
									else
									if((r_sys_run_step==9'h178)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3288[14:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1098[14:0] );

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1500[14:0] );

									end
									else
									if((r_sys_run_step==9'h8d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1878[14:0] );

									end
									else
									if((r_sys_run_step==9'h179)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3294[14:0] );

									end
									else
									if((r_sys_run_step==9'hd2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2292[14:0] );

									end
									else
									if((r_sys_run_step==9'h171) || (r_sys_run_step==9'h173)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3246[14:0] );

									end
									else
									if((r_sys_run_step==9'h103)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2586[14:0] );

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1398[14:0] );

									end
									else
									if((r_sys_run_step==9'h36)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1356[14:0] );

									end
									else
									if((r_sys_run_step==9'h18f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3426[14:0] );

									end
									else
									if((r_sys_run_step==9'h72)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1716[14:0] );

									end
									else
									if((r_sys_run_step==9'h73)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1722[14:0] );

									end
									else
									if((r_sys_run_step==9'h6d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1686[14:0] );

									end
									else
									if((r_sys_run_step==9'h13e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2940[14:0] );

									end
									else
									if((r_sys_run_step==9'h5f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1602[14:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1050[14:0] );

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1536[14:0] );

									end
									else
									if((r_sys_run_step==9'h23)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1242[14:0] );

									end
									else
									if((r_sys_run_step==9'he6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2412[14:0] );

									end
									else
									if((r_sys_run_step==9'h131)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2862[14:0] );

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1524[14:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1128[14:0] );

									end
									else
									if((r_sys_run_step==9'he7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2418[14:0] );

									end
									else
									if((r_sys_run_step==9'h9a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1956[14:0] );

									end
									else
									if((r_sys_run_step==9'h18b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3402[14:0] );

									end
									else
									if((r_sys_run_step==9'h4f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1506[14:0] );

									end
									else
									if((r_sys_run_step==9'hc9) || (r_sys_run_step==9'hcb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2238[14:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1134[14:0] );

									end
									else
									if((r_sys_run_step==9'h11e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2748[14:0] );

									end
									else
									if((r_sys_run_step==9'h60)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1608[14:0] );

									end
									else
									if((r_sys_run_step==9'h69)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1662[14:0] );

									end
									else
									if((r_sys_run_step==9'he8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2424[14:0] );

									end
									else
									if((r_sys_run_step==9'hbc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2160[14:0] );

									end
									else
									if((r_sys_run_step==9'ha5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2022[14:0] );

									end
									else
									if((r_sys_run_step==9'h7e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1788[14:0] );

									end
									else
									if((r_sys_run_step==9'hbd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2166[14:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1176[14:0] );

									end
									else
									if((r_sys_run_step==9'h183)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3354[14:0] );

									end
									else
									if((r_sys_run_step==9'ha6) || (r_sys_run_step==9'ha8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2028[14:0] );

									end
									else
									if((r_sys_run_step==9'h5b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1578[14:0] );

									end
									else
									if((r_sys_run_step==9'hd5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2310[14:0] );

									end
									else
									if((r_sys_run_step==9'h17c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3312[14:0] );

									end
									else
									if((r_sys_run_step==9'hff)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2562[14:0] );

									end
									else
									if((r_sys_run_step==9'h5e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1596[14:0] );

									end
									else
									if((r_sys_run_step==9'h139)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2910[14:0] );

									end
									else
									if((r_sys_run_step==9'hfc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2544[14:0] );

									end
									else
									if((r_sys_run_step==9'hbb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2154[14:0] );

									end
									else
									if((r_sys_run_step==9'h5c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1584[14:0] );

									end
									else
									if((r_sys_run_step==9'h186)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3372[14:0] );

									end
									else
									if((r_sys_run_step==9'h172) || (r_sys_run_step==9'h174)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3252[14:0] );

									end
									else
									if((r_sys_run_step==9'h71)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1710[14:0] );

									end
									else
									if((r_sys_run_step==9'hf1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2478[14:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1170[14:0] );

									end
									else
									if((r_sys_run_step==9'hc3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2202[14:0] );

									end
									else
									if((r_sys_run_step==9'h10f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2658[14:0] );

									end
									else
									if((r_sys_run_step==9'h7c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1776[14:0] );

									end
									else
									if((r_sys_run_step==9'h92)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1908[14:0] );

									end
									else
									if((r_sys_run_step==9'h177)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3282[14:0] );

									end
									else
									if((r_sys_run_step==9'h106)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2604[14:0] );

									end
									else
									if((r_sys_run_step==9'hb4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2112[14:0] );

									end
									else
									if((r_sys_run_step==9'h125)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2790[14:0] );

									end
									else
									if((r_sys_run_step==9'h32)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1332[14:0] );

									end
									else
									if((r_sys_run_step==9'h93)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1914[14:0] );

									end
									else
									if((r_sys_run_step==9'h111)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2670[14:0] );

									end
									else
									if((r_sys_run_step==9'h121)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2766[14:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1062[14:0] );

									end
									else
									if((r_sys_run_step==9'h16c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3216[14:0] );

									end
									else
									if((r_sys_run_step==9'h108)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2616[14:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1074[14:0] );

									end
									else
									if((r_sys_run_step==9'hc1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2190[14:0] );

									end
									else
									if((r_sys_run_step==9'h82)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1812[14:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1188[14:0] );

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1254[14:0] );

									end
									else
									if((r_sys_run_step==9'h75)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1734[14:0] );

									end
									else
									if((r_sys_run_step==9'h9d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1974[14:0] );

									end
									else
									if((r_sys_run_step==9'h163)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3162[14:0] );

									end
									else
									if((r_sys_run_step==9'h10a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2628[14:0] );

									end
									else
									if((r_sys_run_step==9'h70)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1704[14:0] );

									end
									else
									if((r_sys_run_step==9'hdc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2352[14:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1158[14:0] );

									end
									else
									if((r_sys_run_step==9'h137)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2898[14:0] );

									end
									else
									if((r_sys_run_step==9'h42) || (r_sys_run_step==9'h44)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1428[14:0] );

									end
									else
									if((r_sys_run_step==9'h34)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1344[14:0] );

									end
									else
									if((r_sys_run_step==9'hbe)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2172[14:0] );

									end
									else
									if((r_sys_run_step==9'h185)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3366[14:0] );

									end
									else
									if((r_sys_run_step==9'h181)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3342[14:0] );

									end
									else
									if((r_sys_run_step==9'hf6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2508[14:0] );

									end
									else
									if((r_sys_run_step==9'h140)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2952[14:0] );

									end
									else
									if((r_sys_run_step==9'h17b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3306[14:0] );

									end
									else
									if((r_sys_run_step==9'h17d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3318[14:0] );

									end
									else
									if((r_sys_run_step==9'hf7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2514[14:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1200[14:0] );

									end
									else
									if((r_sys_run_step==9'hab)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2058[14:0] );

									end
									else
									if((r_sys_run_step==9'h17e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3324[14:0] );

									end
									else
									if((r_sys_run_step==9'h41) || (r_sys_run_step==9'h43)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1422[14:0] );

									end
									else
									if((r_sys_run_step==9'h11c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2736[14:0] );

									end
									else
									if((r_sys_run_step==9'h11b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2730[14:0] );

									end
									else
									if((r_sys_run_step==9'h187)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3378[14:0] );

									end
									else
									if((r_sys_run_step==9'h15d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3126[14:0] );

									end
									else
									if((r_sys_run_step==9'h148)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3000[14:0] );

									end
									else
									if((r_sys_run_step==9'h4d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1494[14:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1182[14:0] );

									end
									else
									if((r_sys_run_step==9'h119)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2718[14:0] );

									end
									else
									if((r_sys_run_step==9'he5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2406[14:0] );

									end
									else
									if((r_sys_run_step==9'h49)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1470[14:0] );

									end
									else
									if((r_sys_run_step==9'h17a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3300[14:0] );

									end
									else
									if((r_sys_run_step==9'h168)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3192[14:0] );

									end
									else
									if((r_sys_run_step==9'h123)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2778[14:0] );

									end
									else
									if((r_sys_run_step==9'h128)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2808[14:0] );

									end
									else
									if((r_sys_run_step==9'h20) || (r_sys_run_step==9'h22)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1224[14:0] );

									end
									else
									if((r_sys_run_step==9'hd3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2298[14:0] );

									end
									else
									if((r_sys_run_step==9'h86)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1836[14:0] );

									end
									else
									if((r_sys_run_step==9'hef)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2466[14:0] );

									end
									else
									if((r_sys_run_step==9'hce)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2268[14:0] );

									end
									else
									if((r_sys_run_step==9'h192)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3444[14:0] );

									end
									else
									if((r_sys_run_step==9'ha3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2010[14:0] );

									end
									else
									if((r_sys_run_step==9'h2b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1290[14:0] );

									end
									else
									if((r_sys_run_step==9'h96)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1932[14:0] );

									end
									else
									if((r_sys_run_step==9'h18c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3408[14:0] );

									end
									else
									if((r_sys_run_step==9'h6e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1692[14:0] );

									end
									else
									if((r_sys_run_step==9'h77)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1746[14:0] );

									end
									else
									if((r_sys_run_step==9'ha4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2016[14:0] );

									end
									else
									if((r_sys_run_step==9'h10d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2646[14:0] );

									end
									else
									if((r_sys_run_step==9'hdd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2358[14:0] );

									end
									else
									if((r_sys_run_step==9'hd0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2280[14:0] );

									end
									else
									if((r_sys_run_step==9'h188)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3384[14:0] );

									end
									else
									if((r_sys_run_step==9'hf9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2526[14:0] );

									end
									else
									if((r_sys_run_step==9'h13f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2946[14:0] );

									end
									else
									if((r_sys_run_step==9'hb0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2088[14:0] );

									end
									else
									if((r_sys_run_step==9'h170)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3240[14:0] );

									end
									else
									if((r_sys_run_step==9'hc0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2184[14:0] );

									end
									else
									if((r_sys_run_step==9'h45)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1446[14:0] );

									end
									else
									if((r_sys_run_step==9'hf0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2472[14:0] );

									end
									else
									if((r_sys_run_step==9'h3a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1380[14:0] );

									end
									else
									if((r_sys_run_step==9'hfb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2538[14:0] );

									end
									else
									if((r_sys_run_step==9'hfa)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2532[14:0] );

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1482[14:0] );

									end
									else
									if((r_sys_run_step==9'h6c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1680[14:0] );

									end
									else
									if((r_sys_run_step==9'h144)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2976[14:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1080[14:0] );

									end
									else
									if((r_sys_run_step==9'h95)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1926[14:0] );

									end
									else
									if((r_sys_run_step==9'hf8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2520[14:0] );

									end
									else
									if((r_sys_run_step==9'h18e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3420[14:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1146[14:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1056[14:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1116[14:0] );

									end
									else
									if((r_sys_run_step==9'h50)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1512[14:0] );

									end
									else
									if((r_sys_run_step==9'h138)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2904[14:0] );

									end
									else
									if((r_sys_run_step==9'h102)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2580[14:0] );

									end
									else
									if((r_sys_run_step==9'h14a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3012[14:0] );

									end
									else
									if((r_sys_run_step==9'h2c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1296[14:0] );

									end
									else
									if((r_sys_run_step==9'h16f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3234[14:0] );

									end
									else
									if((r_sys_run_step==9'h38)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1368[14:0] );

									end
									else
									if((r_sys_run_step==9'h27)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1266[14:0] );

									end
									else
									if((r_sys_run_step==9'h2a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1284[14:0] );

									end
									else
									if((r_sys_run_step==9'h136)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2892[14:0] );

									end
									else
									if((r_sys_run_step==9'h81)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1806[14:0] );

									end
									else
									if((r_sys_run_step==9'had)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2070[14:0] );

									end
									else
									if((r_sys_run_step==9'h13d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2934[14:0] );

									end
									else
									if((r_sys_run_step==9'h8b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1866[14:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1164[14:0] );

									end
									else
									if((r_sys_run_step==9'h191)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3438[14:0] );

									end
									else
									if((r_sys_run_step==9'hf4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2496[14:0] );

									end
									else
									if((r_sys_run_step==9'h147)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2994[14:0] );

									end
									else
									if((r_sys_run_step==9'h133)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2874[14:0] );

									end
									else
									if((r_sys_run_step==9'h56)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1548[14:0] );

									end
									else
									if((r_sys_run_step==9'h53)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1530[14:0] );

									end
									else
									if((r_sys_run_step==9'hb3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2106[14:0] );

									end
									else
									if((r_sys_run_step==9'h13a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2916[14:0] );

									end
									else
									if((r_sys_run_step==9'h15a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3108[14:0] );

									end
									else
									if((r_sys_run_step==9'h29)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1278[14:0] );

									end
									else
									if((r_sys_run_step==9'h78)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1752[14:0] );

									end
									else
									if((r_sys_run_step==9'h175)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3270[14:0] );

									end
									else
									if((r_sys_run_step==9'ha7) || (r_sys_run_step==9'ha9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2034[14:0] );

									end
									else
									if((r_sys_run_step==9'h114)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2688[14:0] );

									end
									else
									if((r_sys_run_step==9'hc4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2208[14:0] );

									end
									else
									if((r_sys_run_step==9'h88)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1848[14:0] );

									end
									else
									if((r_sys_run_step==9'h165)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3174[14:0] );

									end
									else
									if((r_sys_run_step==9'hee)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2460[14:0] );

									end
									else
									if((r_sys_run_step==9'h7d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1782[14:0] );

									end
									else
									if((r_sys_run_step==9'hc5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2214[14:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1104[14:0] );

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1314[14:0] );

									end
									else
									if((r_sys_run_step==9'h129)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2814[14:0] );

									end
									else
									if((r_sys_run_step==9'h8c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1872[14:0] );

									end
									else
									if((r_sys_run_step==9'h5d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1590[14:0] );

									end
									else
									if((r_sys_run_step==9'h51)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1518[14:0] );

									end
									else
									if((r_sys_run_step==9'h12a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2820[14:0] );

									end
									else
									if((r_sys_run_step==9'h142)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2964[14:0] );

									end
									else
									if((r_sys_run_step==9'h14b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3018[14:0] );

									end
									else
									if((r_sys_run_step==9'h91)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1902[14:0] );

									end
									else
									if((r_sys_run_step==9'h158)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3096[14:0] );

									end
									else
									if((r_sys_run_step==9'h11a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2724[14:0] );

									end
									else
									if((r_sys_run_step==9'h48)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1464[14:0] );

									end
									else
									if((r_sys_run_step==9'hac)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2064[14:0] );

									end
									else
									if((r_sys_run_step==9'he0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2376[14:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1122[14:0] );

									end
									else
									if((r_sys_run_step==9'h90)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1896[14:0] );

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1488[14:0] );

									end
									else
									if((r_sys_run_step==9'h149)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3006[14:0] );

									end
									else
									if((r_sys_run_step==9'hb9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2142[14:0] );

									end
									else
									if((r_sys_run_step==9'h162)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3156[14:0] );

									end
									else
									if((r_sys_run_step==9'h57)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1554[14:0] );

									end
									else
									if((r_sys_run_step==9'h105)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2598[14:0] );

									end
									else
									if((r_sys_run_step==9'hc8) || (r_sys_run_step==9'hca)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2232[14:0] );

									end
									else
									if((r_sys_run_step==9'h67)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1650[14:0] );

									end
									else
									if((r_sys_run_step==9'h74)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1728[14:0] );

									end
									else
									if((r_sys_run_step==9'h143)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2970[14:0] );

									end
									else
									if((r_sys_run_step==9'hf5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2502[14:0] );

									end
									else
									if((r_sys_run_step==9'hdf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2370[14:0] );

									end
									else
									if((r_sys_run_step==9'hf2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2484[14:0] );

									end
									else
									if((r_sys_run_step==9'h46)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1452[14:0] );

									end
									else
									if((r_sys_run_step==9'h98)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1944[14:0] );

									end
									else
									if((r_sys_run_step==9'h14f) || (r_sys_run_step==9'h151)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3042[14:0] );

									end
									else
									if((r_sys_run_step==9'hdb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2346[14:0] );

									end
									else
									if((r_sys_run_step==9'h80)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1800[14:0] );

									end
									else
									if((r_sys_run_step==9'h146)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2988[14:0] );

									end
									else
									if((r_sys_run_step==9'heb) || (r_sys_run_step==9'hed)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2442[14:0] );

									end
									else
									if((r_sys_run_step==9'h15c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3120[14:0] );

									end
									else
									if((r_sys_run_step==9'h13b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2922[14:0] );

									end
									else
									if((r_sys_run_step==9'h76)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1740[14:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1068[14:0] );

									end
									else
									if((r_sys_run_step==9'hbf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2178[14:0] );

									end
									else
									if((r_sys_run_step==9'h12b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2826[14:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1206[14:0] );

									end
									else
									if((r_sys_run_step==9'hcd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2262[14:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1140[14:0] );

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1386[14:0] );

									end
									else
									if((r_sys_run_step==9'hd6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2316[14:0] );

									end
									else
									if((r_sys_run_step==9'h99)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1950[14:0] );

									end
									else
									if((r_sys_run_step==9'h62)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1620[14:0] );

									end
									else
									if((r_sys_run_step==9'hb5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2118[14:0] );

									end
									else
									if((r_sys_run_step==9'h189)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3390[14:0] );

									end
									else
									if((r_sys_run_step==9'h117)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2706[14:0] );

									end
									else
									if((r_sys_run_step==9'h10c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2640[14:0] );

									end
									else
									if((r_sys_run_step==9'h109)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2622[14:0] );

									end
									else
									if((r_sys_run_step==9'hd7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2322[14:0] );

									end
									else
									if((r_sys_run_step==9'h55)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1542[14:0] );

									end
									else
									if((r_sys_run_step==9'h9e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1980[14:0] );

									end
									else
									if((r_sys_run_step==9'he3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2394[14:0] );

									end
									else
									if((r_sys_run_step==9'h37)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1362[14:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1212[14:0] );

									end
									else
									if((r_sys_run_step==9'h18d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3414[14:0] );

									end
									else
									if((r_sys_run_step==9'he4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2400[14:0] );

									end
									else
									if((r_sys_run_step==9'h6a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1668[14:0] );

									end
									else
									if((r_sys_run_step==9'h2e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1308[14:0] );

									end
									else
									if((r_sys_run_step==9'h194)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3456[14:0] );

									end
									else
									if((r_sys_run_step==9'h3f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1410[14:0] );

									end
									else
									if((r_sys_run_step==9'hae)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2076[14:0] );

									end
									else
									if((r_sys_run_step==9'h68)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1656[14:0] );

									end
									else
									if((r_sys_run_step==9'h3e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1404[14:0] );

									end
									else
									if((r_sys_run_step==9'h113)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2682[14:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1044[14:0] );

									end
									else
									if((r_sys_run_step==9'h14d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3030[14:0] );

									end
									else
									if((r_sys_run_step==9'h18a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3396[14:0] );

									end
									else
									if((r_sys_run_step==9'h169)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3198[14:0] );

									end
									else
									if((r_sys_run_step==9'h120)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2760[14:0] );

									end
									else
									if((r_sys_run_step==9'h14c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3024[14:0] );

									end
									else
									if((r_sys_run_step==9'h126)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2796[14:0] );

									end
									else
									if((r_sys_run_step==9'h9c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1968[14:0] );

									end
									else
									if((r_sys_run_step==9'haf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2082[14:0] );

									end
									else
									if((r_sys_run_step==9'h59)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1566[14:0] );

									end
									else
									if((r_sys_run_step==9'h154)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3072[14:0] );

									end
									else
									if((r_sys_run_step==9'h110)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2664[14:0] );

									end
									else
									if((r_sys_run_step==9'h190)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3432[14:0] );

									end
									else
									if((r_sys_run_step==9'h6f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1698[14:0] );

									end
									else
									if((r_sys_run_step==9'h79)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1758[14:0] );

									end
									else
									if((r_sys_run_step==9'h15b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3114[14:0] );

									end
									else
									if((r_sys_run_step==9'h145)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2982[14:0] );

									end
									else
									if((r_sys_run_step==9'h124)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2784[14:0] );

									end
									else
									if((r_sys_run_step==9'h11d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2742[14:0] );

									end
									else
									if((r_sys_run_step==9'h100)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2568[14:0] );

									end
									else
									if((r_sys_run_step==9'ha0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1992[14:0] );

									end
									else
									if((r_sys_run_step==9'hc6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2220[14:0] );

									end
									else
									if((r_sys_run_step==9'h107)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2610[14:0] );

									end
									else
									if((r_sys_run_step==9'hb7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2130[14:0] );

									end
									else
									if((r_sys_run_step==9'h15e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3132[14:0] );

									end
									else
									if((r_sys_run_step==9'h155)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3078[14:0] );

									end
									else
									if((r_sys_run_step==9'hde)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2364[14:0] );

									end
									else
									if((r_sys_run_step==9'h31)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1326[14:0] );

									end
									else
									if((r_sys_run_step==9'h8f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1890[14:0] );

									end
									else
									if((r_sys_run_step==9'h122)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2772[14:0] );

									end
									else
									if((r_sys_run_step==9'h10e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2652[14:0] );

									end
									else
									if((r_sys_run_step==9'h16b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3210[14:0] );

									end
									else
									if((r_sys_run_step==9'hcf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2274[14:0] );

									end
									else
									if((r_sys_run_step==9'ha1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1998[14:0] );

									end
									else
									if((r_sys_run_step==9'h156)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3084[14:0] );

									end
									else
									if((r_sys_run_step==9'h85)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1830[14:0] );

									end
									else
									if((r_sys_run_step==9'hea) || (r_sys_run_step==9'hec)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2436[14:0] );

									end
									else
									if((r_sys_run_step==9'hb6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2124[14:0] );

									end
									else
									if((r_sys_run_step==9'h176)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3276[14:0] );

									end
									else
									if((r_sys_run_step==9'h160)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3144[14:0] );

									end
									else
									if((r_sys_run_step==9'h17f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3330[14:0] );

									end
									else
									if((r_sys_run_step==9'h116)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2700[14:0] );

									end
									else
									if((r_sys_run_step==9'h141)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2958[14:0] );

									end
									else
									if((r_sys_run_step==9'h4a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1476[14:0] );

									end
									else
									if((r_sys_run_step==9'h182)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3348[14:0] );

									end
									else
									if((r_sys_run_step==9'h13c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2928[14:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1194[14:0] );

									end
									else
									if((r_sys_run_step==9'h135)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2886[14:0] );

									end
									else
									if((r_sys_run_step==9'h12d) || (r_sys_run_step==9'h12f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2838[14:0] );

									end
									else
									if((r_sys_run_step==9'h115)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2694[14:0] );

									end
									else
									if((r_sys_run_step==9'h10b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2634[14:0] );

									end
									else
									if((r_sys_run_step==9'he1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2382[14:0] );

									end
									else
									if((r_sys_run_step==9'h8e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1884[14:0] );

									end
									else
									if((r_sys_run_step==9'h118)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2712[14:0] );

									end
									else
									if((r_sys_run_step==9'hfd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2550[14:0] );

									end
									else
									if((r_sys_run_step==9'h35)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1350[14:0] );

									end
									else
									if((r_sys_run_step==9'h6b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1674[14:0] );

									end
									else
									if((r_sys_run_step==9'h9f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1986[14:0] );

									end
									else
									if((r_sys_run_step==9'h153)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3066[14:0] );

									end
									else
									if((r_sys_run_step==9'h150) || (r_sys_run_step==9'h152)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3048[14:0] );

									end
									else
									if((r_sys_run_step==9'h159)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3102[14:0] );

									end
									else
									if((r_sys_run_step==9'hc2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2196[14:0] );

									end
									else
									if((r_sys_run_step==9'h63) || (r_sys_run_step==9'h65)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1626[14:0] );

									end
									else
									if((r_sys_run_step==9'h30)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1320[14:0] );

									end
									else
									if((r_sys_run_step==9'h157)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3090[14:0] );

									end
									else
									if((r_sys_run_step==9'h97)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1938[14:0] );

									end
									else
									if((r_sys_run_step==9'h64) || (r_sys_run_step==9'h66)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1632[14:0] );

									end
									else
									if((r_sys_run_step==9'h184)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3360[14:0] );

									end
									else
									if((r_sys_run_step==9'hb8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2136[14:0] );

									end
									else
									if((r_sys_run_step==9'hd8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2328[14:0] );

									end
									else
									if((r_sys_run_step==9'h7a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1764[14:0] );

									end
									else
									if((r_sys_run_step==9'h61)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1614[14:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1032[14:0] );

									end
									else
									if((r_sys_run_step==9'hd9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2334[14:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1038[14:0] );

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1392[14:0] );

									end
									else
									if((r_sys_run_step==9'h161)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3150[14:0] );

									end
									else
									if((r_sys_run_step==9'hda)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2340[14:0] );

									end
									else
									if((r_sys_run_step==9'h8a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1860[14:0] );

									end
									else
									if((r_sys_run_step==9'h104)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2592[14:0] );

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1248[14:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1086[14:0] );

									end
									else
									if((r_sys_run_step==9'hf3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2490[14:0] );

									end
									else
									if((r_sys_run_step==9'h9b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1962[14:0] );

									end
									else
									if((r_sys_run_step==9'haa)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2052[14:0] );

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1458[14:0] );

									end
									else
									if((r_sys_run_step==9'h1f) || (r_sys_run_step==9'h21)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1218[14:0] );

									end
									else
									if((r_sys_run_step==9'h83)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1818[14:0] );

									end
									else
									if((r_sys_run_step==9'h193)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3450[14:0] );

									end
									else
									if((r_sys_run_step==9'hba)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2148[14:0] );

									end
									else
									if((r_sys_run_step==9'ha2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2004[14:0] );

									end
									else
									if((r_sys_run_step==9'h127)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2802[14:0] );

									end
									else
									if((r_sys_run_step==9'h5a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1572[14:0] );

									end
									else
									if((r_sys_run_step==9'h7b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1770[14:0] );

									end
									else
									if((r_sys_run_step==9'hb2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2100[14:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1092[14:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1152[14:0] );

									end
									else
									if((r_sys_run_step==9'h89)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1854[14:0] );

									end
									else
									if((r_sys_run_step==9'h166)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3180[14:0] );

									end
									else
									if((r_sys_run_step==9'h58)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1560[14:0] );

									end
									else
									if((r_sys_run_step==9'hb1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2094[14:0] );

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h69)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4014[14:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3510[14:0] );

									end
									else
									if((r_sys_run_step==9'h7f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4124[14:0] );

									end
									else
									if((r_sys_run_step==9'h23)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3664[14:0] );

									end
									else
									if((r_sys_run_step==9'h61)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3974[14:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3558[14:0] );

									end
									else
									if((r_sys_run_step==9'h4d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3874[14:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3504[14:0] );

									end
									else
									if((r_sys_run_step==9'h6f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4044[14:0] );

									end
									else
									if((r_sys_run_step==9'h22)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3659[14:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3576[14:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3516[14:0] );

									end
									else
									if((r_sys_run_step==9'h6a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4019[14:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3630[14:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3642[14:0] );

									end
									else
									if((r_sys_run_step==9'h73)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4064[14:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3546[14:0] );

									end
									else
									if((r_sys_run_step==9'h64)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3989[14:0] );

									end
									else
									if((r_sys_run_step==9'h79)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4094[14:0] );

									end
									else
									if((r_sys_run_step==9'h20)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3648[14:0] );

									end
									else
									if((r_sys_run_step==9'h40)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3809[14:0] );

									end
									else
									if((r_sys_run_step==9'h42)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3819[14:0] );

									end
									else
									if((r_sys_run_step==9'h5a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3939[14:0] );

									end
									else
									if((r_sys_run_step==9'h27)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3684[14:0] );

									end
									else
									if((r_sys_run_step==9'h58)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3929[14:0] );

									end
									else
									if((r_sys_run_step==9'h35)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3754[14:0] );

									end
									else
									if((r_sys_run_step==9'h7a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4099[14:0] );

									end
									else
									if((r_sys_run_step==9'h6b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4024[14:0] );

									end
									else
									if((r_sys_run_step==9'h59)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3934[14:0] );

									end
									else
									if((r_sys_run_step==9'h77)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4084[14:0] );

									end
									else
									if((r_sys_run_step==9'h7e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4119[14:0] );

									end
									else
									if((r_sys_run_step==9'h3f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3804[14:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3618[14:0] );

									end
									else
									if((r_sys_run_step==9'h75)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4074[14:0] );

									end
									else
									if((r_sys_run_step==9'h78)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4089[14:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3528[14:0] );

									end
									else
									if((r_sys_run_step==9'h7d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4114[14:0] );

									end
									else
									if((r_sys_run_step==9'h71)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4054[14:0] );

									end
									else
									if((r_sys_run_step==9'h2a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3699[14:0] );

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3784[14:0] );

									end
									else
									if((r_sys_run_step==9'h51)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3894[14:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3492[14:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3600[14:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3588[14:0] );

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3864[14:0] );

									end
									else
									if((r_sys_run_step==9'h60)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3969[14:0] );

									end
									else
									if((r_sys_run_step==9'h32)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3739[14:0] );

									end
									else
									if((r_sys_run_step==9'h41)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3814[14:0] );

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3674[14:0] );

									end
									else
									if((r_sys_run_step==9'h21)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3654[14:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3486[14:0] );

									end
									else
									if((r_sys_run_step==9'h48)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3849[14:0] );

									end
									else
									if((r_sys_run_step==9'h68)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4009[14:0] );

									end
									else
									if((r_sys_run_step==9'h7b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4104[14:0] );

									end
									else
									if((r_sys_run_step==9'h33)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3744[14:0] );

									end
									else
									if((r_sys_run_step==9'h43)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3824[14:0] );

									end
									else
									if((r_sys_run_step==9'h56)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3919[14:0] );

									end
									else
									if((r_sys_run_step==9'h5d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3954[14:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3540[14:0] );

									end
									else
									if((r_sys_run_step==9'h50)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3889[14:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3468[14:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3594[14:0] );

									end
									else
									if((r_sys_run_step==9'h6e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4039[14:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3612[14:0] );

									end
									else
									if((r_sys_run_step==9'h65)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3994[14:0] );

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3844[14:0] );

									end
									else
									if((r_sys_run_step==9'h63)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3984[14:0] );

									end
									else
									if((r_sys_run_step==9'h57)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3924[14:0] );

									end
									else
									if((r_sys_run_step==9'h45)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3834[14:0] );

									end
									else
									if((r_sys_run_step==9'h2b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3704[14:0] );

									end
									else
									if((r_sys_run_step==9'h31)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3734[14:0] );

									end
									else
									if((r_sys_run_step==9'h34)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3749[14:0] );

									end
									else
									if((r_sys_run_step==9'h49)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3854[14:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3534[14:0] );

									end
									else
									if((r_sys_run_step==9'h5e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3959[14:0] );

									end
									else
									if((r_sys_run_step==9'h7c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4109[14:0] );

									end
									else
									if((r_sys_run_step==9'h5f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3964[14:0] );

									end
									else
									if((r_sys_run_step==9'h4a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3859[14:0] );

									end
									else
									if((r_sys_run_step==9'h2e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3719[14:0] );

									end
									else
									if((r_sys_run_step==9'h2c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3709[14:0] );

									end
									else
									if((r_sys_run_step==9'h66)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3999[14:0] );

									end
									else
									if((r_sys_run_step==9'h30)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3729[14:0] );

									end
									else
									if((r_sys_run_step==9'h36)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3759[14:0] );

									end
									else
									if((r_sys_run_step==9'h76)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4079[14:0] );

									end
									else
									if((r_sys_run_step==9'h6d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4034[14:0] );

									end
									else
									if((r_sys_run_step==9'h6c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4029[14:0] );

									end
									else
									if((r_sys_run_step==9'h53)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3904[14:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3564[14:0] );

									end
									else
									if((r_sys_run_step==9'h37)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3764[14:0] );

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3899[14:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3582[14:0] );

									end
									else
									if((r_sys_run_step==9'h29)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3694[14:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3552[14:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3480[14:0] );

									end
									else
									if((r_sys_run_step==9'h72)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4059[14:0] );

									end
									else
									if((r_sys_run_step==9'h67)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4004[14:0] );

									end
									else
									if((r_sys_run_step==9'h62)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3979[14:0] );

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3669[14:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3498[14:0] );

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3794[14:0] );

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3909[14:0] );

									end
									else
									if((r_sys_run_step==9'h3e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3799[14:0] );

									end
									else
									if((r_sys_run_step==9'h5b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3944[14:0] );

									end
									else
									if((r_sys_run_step==9'h28)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3689[14:0] );

									end
									else
									if((r_sys_run_step==9'h55)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3914[14:0] );

									end
									else
									if((r_sys_run_step==9'h2d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3714[14:0] );

									end
									else
									if((r_sys_run_step==9'h46)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3839[14:0] );

									end
									else
									if((r_sys_run_step==9'h5c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3949[14:0] );

									end
									else
									if((r_sys_run_step==9'h44)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3829[14:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3636[14:0] );

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3869[14:0] );

									end
									else
									if((r_sys_run_step==9'h26)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3679[14:0] );

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3789[14:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3474[14:0] );

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3879[14:0] );

									end
									else
									if((r_sys_run_step==9'h38)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3769[14:0] );

									end
									else
									if((r_sys_run_step==9'h3a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3779[14:0] );

									end
									else
									if((r_sys_run_step==9'h4f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3884[14:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3570[14:0] );

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3774[14:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3624[14:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3606[14:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3522[14:0] );

									end
									else
									if((r_sys_run_step==9'h80)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4129[14:0] );

									end
									else
									if((r_sys_run_step==9'h70)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4049[14:0] );

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3724[14:0] );

									end
									else
									if((r_sys_run_step==9'h74)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4069[14:0] );

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h65)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4666[14:0] );

									end
									else
									if((r_sys_run_step==9'h9f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4956[14:0] );

									end
									else
									if((r_sys_run_step==9'h8d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4866[14:0] );

									end
									else
									if((r_sys_run_step==9'h97)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4916[14:0] );

									end
									else
									if((r_sys_run_step==9'hde)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5271[14:0] );

									end
									else
									if((r_sys_run_step==9'hdb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5256[14:0] );

									end
									else
									if((r_sys_run_step==9'h42)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4491[14:0] );

									end
									else
									if((r_sys_run_step==9'h149)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5806[14:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4254[14:0] );

									end
									else
									if((r_sys_run_step==9'h5e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4631[14:0] );

									end
									else
									if((r_sys_run_step==9'h8f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4876[14:0] );

									end
									else
									if((r_sys_run_step==9'h11c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5581[14:0] );

									end
									else
									if((r_sys_run_step==9'h107)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5476[14:0] );

									end
									else
									if((r_sys_run_step==9'h8e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4871[14:0] );

									end
									else
									if((r_sys_run_step==9'hcc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5181[14:0] );

									end
									else
									if((r_sys_run_step==9'h62)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4651[14:0] );

									end
									else
									if((r_sys_run_step==9'h6e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4711[14:0] );

									end
									else
									if((r_sys_run_step==9'h6a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4691[14:0] );

									end
									else
									if((r_sys_run_step==9'h59)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4606[14:0] );

									end
									else
									if((r_sys_run_step==9'h17d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp6066[14:0] );

									end
									else
									if((r_sys_run_step==9'h13c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5741[14:0] );

									end
									else
									if((r_sys_run_step==9'hbd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5106[14:0] );

									end
									else
									if((r_sys_run_step==9'h167)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5956[14:0] );

									end
									else
									if((r_sys_run_step==9'hf1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5366[14:0] );

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4581[14:0] );

									end
									else
									if((r_sys_run_step==9'h5c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4621[14:0] );

									end
									else
									if((r_sys_run_step==9'h105)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5466[14:0] );

									end
									else
									if((r_sys_run_step==9'h4f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4556[14:0] );

									end
									else
									if((r_sys_run_step==9'h14f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5836[14:0] );

									end
									else
									if((r_sys_run_step==9'h92)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4891[14:0] );

									end
									else
									if((r_sys_run_step==9'h9b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4936[14:0] );

									end
									else
									if((r_sys_run_step==9'h71)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4726[14:0] );

									end
									else
									if((r_sys_run_step==9'hf4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5381[14:0] );

									end
									else
									if((r_sys_run_step==9'h46)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4511[14:0] );

									end
									else
									if((r_sys_run_step==9'hd9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5246[14:0] );

									end
									else
									if((r_sys_run_step==9'h9a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4931[14:0] );

									end
									else
									if((r_sys_run_step==9'h11e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5591[14:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4170[14:0] );

									end
									else
									if((r_sys_run_step==9'h127)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5636[14:0] );

									end
									else
									if((r_sys_run_step==9'hfb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5416[14:0] );

									end
									else
									if((r_sys_run_step==9'h63)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4656[14:0] );

									end
									else
									if((r_sys_run_step==9'h10c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5501[14:0] );

									end
									else
									if((r_sys_run_step==9'h12f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5676[14:0] );

									end
									else
									if((r_sys_run_step==9'he1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5286[14:0] );

									end
									else
									if((r_sys_run_step==9'hb1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5046[14:0] );

									end
									else
									if((r_sys_run_step==9'h5d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4626[14:0] );

									end
									else
									if((r_sys_run_step==9'h51)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4566[14:0] );

									end
									else
									if((r_sys_run_step==9'ha7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4996[14:0] );

									end
									else
									if((r_sys_run_step==9'h170)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp6001[14:0] );

									end
									else
									if((r_sys_run_step==9'ha6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4991[14:0] );

									end
									else
									if((r_sys_run_step==9'h169)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5966[14:0] );

									end
									else
									if((r_sys_run_step==9'h12b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5656[14:0] );

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4551[14:0] );

									end
									else
									if((r_sys_run_step==9'h53)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4576[14:0] );

									end
									else
									if((r_sys_run_step==9'he0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5281[14:0] );

									end
									else
									if((r_sys_run_step==9'h82)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4811[14:0] );

									end
									else
									if((r_sys_run_step==9'h112)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5531[14:0] );

									end
									else
									if((r_sys_run_step==9'h2d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4386[14:0] );

									end
									else
									if((r_sys_run_step==9'h94)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4901[14:0] );

									end
									else
									if((r_sys_run_step==9'hab)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5016[14:0] );

									end
									else
									if((r_sys_run_step==9'hce)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5191[14:0] );

									end
									else
									if((r_sys_run_step==9'h61)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4646[14:0] );

									end
									else
									if((r_sys_run_step==9'h99)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4926[14:0] );

									end
									else
									if((r_sys_run_step==9'h103)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5456[14:0] );

									end
									else
									if((r_sys_run_step==9'h2e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4391[14:0] );

									end
									else
									if((r_sys_run_step==9'he3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5296[14:0] );

									end
									else
									if((r_sys_run_step==9'h9c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4941[14:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4248[14:0] );

									end
									else
									if((r_sys_run_step==9'h171)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp6006[14:0] );

									end
									else
									if((r_sys_run_step==9'h120)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5601[14:0] );

									end
									else
									if((r_sys_run_step==9'hd5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5226[14:0] );

									end
									else
									if((r_sys_run_step==9'h60)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4641[14:0] );

									end
									else
									if((r_sys_run_step==9'h115)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5546[14:0] );

									end
									else
									if((r_sys_run_step==9'hae)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5031[14:0] );

									end
									else
									if((r_sys_run_step==9'h7f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4796[14:0] );

									end
									else
									if((r_sys_run_step==9'h126)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5631[14:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4242[14:0] );

									end
									else
									if((r_sys_run_step==9'h132)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5691[14:0] );

									end
									else
									if((r_sys_run_step==9'h55)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4586[14:0] );

									end
									else
									if((r_sys_run_step==9'h32)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4411[14:0] );

									end
									else
									if((r_sys_run_step==9'hd4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5221[14:0] );

									end
									else
									if((r_sys_run_step==9'h40)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4481[14:0] );

									end
									else
									if((r_sys_run_step==9'h83)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4816[14:0] );

									end
									else
									if((r_sys_run_step==9'h37)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4436[14:0] );

									end
									else
									if((r_sys_run_step==9'h86)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4831[14:0] );

									end
									else
									if((r_sys_run_step==9'ha2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4971[14:0] );

									end
									else
									if((r_sys_run_step==9'h8b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4856[14:0] );

									end
									else
									if((r_sys_run_step==9'h98)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4921[14:0] );

									end
									else
									if((r_sys_run_step==9'h176)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp6031[14:0] );

									end
									else
									if((r_sys_run_step==9'h108)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5481[14:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4200[14:0] );

									end
									else
									if((r_sys_run_step==9'hfa)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5411[14:0] );

									end
									else
									if((r_sys_run_step==9'h106)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5471[14:0] );

									end
									else
									if((r_sys_run_step==9'h122)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5611[14:0] );

									end
									else
									if((r_sys_run_step==9'hc7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5156[14:0] );

									end
									else
									if((r_sys_run_step==9'h15a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5891[14:0] );

									end
									else
									if((r_sys_run_step==9'h100)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5441[14:0] );

									end
									else
									if((r_sys_run_step==9'had)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5026[14:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4236[14:0] );

									end
									else
									if((r_sys_run_step==9'h23)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4336[14:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4314[14:0] );

									end
									else
									if((r_sys_run_step==9'hcf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5196[14:0] );

									end
									else
									if((r_sys_run_step==9'hb5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5066[14:0] );

									end
									else
									if((r_sys_run_step==9'hb8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5081[14:0] );

									end
									else
									if((r_sys_run_step==9'h17b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp6056[14:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4230[14:0] );

									end
									else
									if((r_sys_run_step==9'h77)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4756[14:0] );

									end
									else
									if((r_sys_run_step==9'h80)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4801[14:0] );

									end
									else
									if((r_sys_run_step==9'h155)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5866[14:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4224[14:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4290[14:0] );

									end
									else
									if((r_sys_run_step==9'h15d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5906[14:0] );

									end
									else
									if((r_sys_run_step==9'h4d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4546[14:0] );

									end
									else
									if((r_sys_run_step==9'h150)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5841[14:0] );

									end
									else
									if((r_sys_run_step==9'h20)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4320[14:0] );

									end
									else
									if((r_sys_run_step==9'h123)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5616[14:0] );

									end
									else
									if((r_sys_run_step==9'h2c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4381[14:0] );

									end
									else
									if((r_sys_run_step==9'h96)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4911[14:0] );

									end
									else
									if((r_sys_run_step==9'heb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5336[14:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4146[14:0] );

									end
									else
									if((r_sys_run_step==9'h35)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4426[14:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4176[14:0] );

									end
									else
									if((r_sys_run_step==9'h156)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5871[14:0] );

									end
									else
									if((r_sys_run_step==9'h102)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5451[14:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4272[14:0] );

									end
									else
									if((r_sys_run_step==9'ha1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4966[14:0] );

									end
									else
									if((r_sys_run_step==9'hb6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5071[14:0] );

									end
									else
									if((r_sys_run_step==9'hcb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5176[14:0] );

									end
									else
									if((r_sys_run_step==9'h30)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4401[14:0] );

									end
									else
									if((r_sys_run_step==9'h34)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4421[14:0] );

									end
									else
									if((r_sys_run_step==9'h27)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4356[14:0] );

									end
									else
									if((r_sys_run_step==9'h10f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5516[14:0] );

									end
									else
									if((r_sys_run_step==9'h6c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4701[14:0] );

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4461[14:0] );

									end
									else
									if((r_sys_run_step==9'h133)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5696[14:0] );

									end
									else
									if((r_sys_run_step==9'h131)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5686[14:0] );

									end
									else
									if((r_sys_run_step==9'h163)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5936[14:0] );

									end
									else
									if((r_sys_run_step==9'h14a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5811[14:0] );

									end
									else
									if((r_sys_run_step==9'h12e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5671[14:0] );

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4516[14:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4194[14:0] );

									end
									else
									if((r_sys_run_step==9'h9e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4951[14:0] );

									end
									else
									if((r_sys_run_step==9'h101)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5446[14:0] );

									end
									else
									if((r_sys_run_step==9'hc9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5166[14:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4284[14:0] );

									end
									else
									if((r_sys_run_step==9'hb2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5051[14:0] );

									end
									else
									if((r_sys_run_step==9'h43)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4496[14:0] );

									end
									else
									if((r_sys_run_step==9'h74)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4741[14:0] );

									end
									else
									if((r_sys_run_step==9'hb3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5056[14:0] );

									end
									else
									if((r_sys_run_step==9'h67)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4676[14:0] );

									end
									else
									if((r_sys_run_step==9'h5f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4636[14:0] );

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4466[14:0] );

									end
									else
									if((r_sys_run_step==9'h178)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp6041[14:0] );

									end
									else
									if((r_sys_run_step==9'hc3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5136[14:0] );

									end
									else
									if((r_sys_run_step==9'h143)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5776[14:0] );

									end
									else
									if((r_sys_run_step==9'h79)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4766[14:0] );

									end
									else
									if((r_sys_run_step==9'h118)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5561[14:0] );

									end
									else
									if((r_sys_run_step==9'h3f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4476[14:0] );

									end
									else
									if((r_sys_run_step==9'h84)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4821[14:0] );

									end
									else
									if((r_sys_run_step==9'hac)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5021[14:0] );

									end
									else
									if((r_sys_run_step==9'hf8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5401[14:0] );

									end
									else
									if((r_sys_run_step==9'hd1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5206[14:0] );

									end
									else
									if((r_sys_run_step==9'h10d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5506[14:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4260[14:0] );

									end
									else
									if((r_sys_run_step==9'h8c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4861[14:0] );

									end
									else
									if((r_sys_run_step==9'hff)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5436[14:0] );

									end
									else
									if((r_sys_run_step==9'h179)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp6046[14:0] );

									end
									else
									if((r_sys_run_step==9'h113)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5536[14:0] );

									end
									else
									if((r_sys_run_step==9'h10b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5496[14:0] );

									end
									else
									if((r_sys_run_step==9'h6b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4696[14:0] );

									end
									else
									if((r_sys_run_step==9'hcd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5186[14:0] );

									end
									else
									if((r_sys_run_step==9'h17e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp6071[14:0] );

									end
									else
									if((r_sys_run_step==9'h158)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5881[14:0] );

									end
									else
									if((r_sys_run_step==9'h16b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5976[14:0] );

									end
									else
									if((r_sys_run_step==9'hc6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5151[14:0] );

									end
									else
									if((r_sys_run_step==9'h11a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5571[14:0] );

									end
									else
									if((r_sys_run_step==9'h164)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5941[14:0] );

									end
									else
									if((r_sys_run_step==9'h142)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5771[14:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4182[14:0] );

									end
									else
									if((r_sys_run_step==9'h12c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5661[14:0] );

									end
									else
									if((r_sys_run_step==9'hfd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5426[14:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4212[14:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4188[14:0] );

									end
									else
									if((r_sys_run_step==9'hb4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5061[14:0] );

									end
									else
									if((r_sys_run_step==9'h148)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5801[14:0] );

									end
									else
									if((r_sys_run_step==9'h13e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5751[14:0] );

									end
									else
									if((r_sys_run_step==9'h130)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5681[14:0] );

									end
									else
									if((r_sys_run_step==9'hf3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5376[14:0] );

									end
									else
									if((r_sys_run_step==9'h144)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5781[14:0] );

									end
									else
									if((r_sys_run_step==9'ha9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5006[14:0] );

									end
									else
									if((r_sys_run_step==9'h128)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5641[14:0] );

									end
									else
									if((r_sys_run_step==9'h16c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5981[14:0] );

									end
									else
									if((r_sys_run_step==9'h75)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4746[14:0] );

									end
									else
									if((r_sys_run_step==9'h7c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4781[14:0] );

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4446[14:0] );

									end
									else
									if((r_sys_run_step==9'ha4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4981[14:0] );

									end
									else
									if((r_sys_run_step==9'h26)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4351[14:0] );

									end
									else
									if((r_sys_run_step==9'hc1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5126[14:0] );

									end
									else
									if((r_sys_run_step==9'h85)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4826[14:0] );

									end
									else
									if((r_sys_run_step==9'h16a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5971[14:0] );

									end
									else
									if((r_sys_run_step==9'hca)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5171[14:0] );

									end
									else
									if((r_sys_run_step==9'h49)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4526[14:0] );

									end
									else
									if((r_sys_run_step==9'h45)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4506[14:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4308[14:0] );

									end
									else
									if((r_sys_run_step==9'he9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5326[14:0] );

									end
									else
									if((r_sys_run_step==9'h78)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4761[14:0] );

									end
									else
									if((r_sys_run_step==9'h12a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5651[14:0] );

									end
									else
									if((r_sys_run_step==9'hef)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5356[14:0] );

									end
									else
									if((r_sys_run_step==9'h29)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4366[14:0] );

									end
									else
									if((r_sys_run_step==9'h13d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5746[14:0] );

									end
									else
									if((r_sys_run_step==9'h145)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5786[14:0] );

									end
									else
									if((r_sys_run_step==9'hfc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5421[14:0] );

									end
									else
									if((r_sys_run_step==9'h172)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp6011[14:0] );

									end
									else
									if((r_sys_run_step==9'hd2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5211[14:0] );

									end
									else
									if((r_sys_run_step==9'h7a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4771[14:0] );

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4396[14:0] );

									end
									else
									if((r_sys_run_step==9'h157)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5876[14:0] );

									end
									else
									if((r_sys_run_step==9'ha5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4986[14:0] );

									end
									else
									if((r_sys_run_step==9'h16d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5986[14:0] );

									end
									else
									if((r_sys_run_step==9'h66)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4671[14:0] );

									end
									else
									if((r_sys_run_step==9'hb7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5076[14:0] );

									end
									else
									if((r_sys_run_step==9'he5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5306[14:0] );

									end
									else
									if((r_sys_run_step==9'h16f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5996[14:0] );

									end
									else
									if((r_sys_run_step==9'h165)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5946[14:0] );

									end
									else
									if((r_sys_run_step==9'h6d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4706[14:0] );

									end
									else
									if((r_sys_run_step==9'he8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5321[14:0] );

									end
									else
									if((r_sys_run_step==9'h44)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4501[14:0] );

									end
									else
									if((r_sys_run_step==9'h13b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5736[14:0] );

									end
									else
									if((r_sys_run_step==9'h12d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5666[14:0] );

									end
									else
									if((r_sys_run_step==9'ha3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4976[14:0] );

									end
									else
									if((r_sys_run_step==9'h136)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5711[14:0] );

									end
									else
									if((r_sys_run_step==9'h129)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5646[14:0] );

									end
									else
									if((r_sys_run_step==9'h173)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp6016[14:0] );

									end
									else
									if((r_sys_run_step==9'h17a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp6051[14:0] );

									end
									else
									if((r_sys_run_step==9'h152)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5851[14:0] );

									end
									else
									if((r_sys_run_step==9'hbb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5096[14:0] );

									end
									else
									if((r_sys_run_step==9'hc0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5121[14:0] );

									end
									else
									if((r_sys_run_step==9'h141)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5766[14:0] );

									end
									else
									if((r_sys_run_step==9'h14e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5831[14:0] );

									end
									else
									if((r_sys_run_step==9'hf6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5391[14:0] );

									end
									else
									if((r_sys_run_step==9'hc5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5146[14:0] );

									end
									else
									if((r_sys_run_step==9'h7b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4776[14:0] );

									end
									else
									if((r_sys_run_step==9'h50)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4561[14:0] );

									end
									else
									if((r_sys_run_step==9'h15b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5896[14:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4278[14:0] );

									end
									else
									if((r_sys_run_step==9'h70)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4721[14:0] );

									end
									else
									if((r_sys_run_step==9'hc2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5131[14:0] );

									end
									else
									if((r_sys_run_step==9'hb0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5041[14:0] );

									end
									else
									if((r_sys_run_step==9'h64)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4661[14:0] );

									end
									else
									if((r_sys_run_step==9'h11d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5586[14:0] );

									end
									else
									if((r_sys_run_step==9'h89)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4846[14:0] );

									end
									else
									if((r_sys_run_step==9'h140)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5761[14:0] );

									end
									else
									if((r_sys_run_step==9'hbf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5116[14:0] );

									end
									else
									if((r_sys_run_step==9'h21)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4326[14:0] );

									end
									else
									if((r_sys_run_step==9'h151)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5846[14:0] );

									end
									else
									if((r_sys_run_step==9'hdf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5276[14:0] );

									end
									else
									if((r_sys_run_step==9'hbc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5101[14:0] );

									end
									else
									if((r_sys_run_step==9'h14b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5816[14:0] );

									end
									else
									if((r_sys_run_step==9'h116)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5551[14:0] );

									end
									else
									if((r_sys_run_step==9'he6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5311[14:0] );

									end
									else
									if((r_sys_run_step==9'h17c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp6061[14:0] );

									end
									else
									if((r_sys_run_step==9'hf7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5396[14:0] );

									end
									else
									if((r_sys_run_step==9'h135)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5706[14:0] );

									end
									else
									if((r_sys_run_step==9'hbe)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5111[14:0] );

									end
									else
									if((r_sys_run_step==9'hfe)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5431[14:0] );

									end
									else
									if((r_sys_run_step==9'h87)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4836[14:0] );

									end
									else
									if((r_sys_run_step==9'h5a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4611[14:0] );

									end
									else
									if((r_sys_run_step==9'h10a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5491[14:0] );

									end
									else
									if((r_sys_run_step==9'h14d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5826[14:0] );

									end
									else
									if((r_sys_run_step==9'h90)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4881[14:0] );

									end
									else
									if((r_sys_run_step==9'he2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5291[14:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4158[14:0] );

									end
									else
									if((r_sys_run_step==9'h15f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5916[14:0] );

									end
									else
									if((r_sys_run_step==9'hdc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5261[14:0] );

									end
									else
									if((r_sys_run_step==9'h119)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5566[14:0] );

									end
									else
									if((r_sys_run_step==9'h168)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5961[14:0] );

									end
									else
									if((r_sys_run_step==9'h72)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4731[14:0] );

									end
									else
									if((r_sys_run_step==9'h109)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5486[14:0] );

									end
									else
									if((r_sys_run_step==9'haf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5036[14:0] );

									end
									else
									if((r_sys_run_step==9'h91)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4886[14:0] );

									end
									else
									if((r_sys_run_step==9'he4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5301[14:0] );

									end
									else
									if((r_sys_run_step==9'h28)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4361[14:0] );

									end
									else
									if((r_sys_run_step==9'h162)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5931[14:0] );

									end
									else
									if((r_sys_run_step==9'h38)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4441[14:0] );

									end
									else
									if((r_sys_run_step==9'hed)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5346[14:0] );

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4536[14:0] );

									end
									else
									if((r_sys_run_step==9'h117)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5556[14:0] );

									end
									else
									if((r_sys_run_step==9'hc4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5141[14:0] );

									end
									else
									if((r_sys_run_step==9'h11b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5576[14:0] );

									end
									else
									if((r_sys_run_step==9'h6f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4716[14:0] );

									end
									else
									if((r_sys_run_step==9'h166)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5951[14:0] );

									end
									else
									if((r_sys_run_step==9'h31)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4406[14:0] );

									end
									else
									if((r_sys_run_step==9'h134)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5701[14:0] );

									end
									else
									if((r_sys_run_step==9'h33)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4416[14:0] );

									end
									else
									if((r_sys_run_step==9'h69)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4686[14:0] );

									end
									else
									if((r_sys_run_step==9'hc8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5161[14:0] );

									end
									else
									if((r_sys_run_step==9'h161)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5926[14:0] );

									end
									else
									if((r_sys_run_step==9'h111)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5526[14:0] );

									end
									else
									if((r_sys_run_step==9'h88)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4841[14:0] );

									end
									else
									if((r_sys_run_step==9'hd6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5231[14:0] );

									end
									else
									if((r_sys_run_step==9'hb9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5086[14:0] );

									end
									else
									if((r_sys_run_step==9'h58)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4601[14:0] );

									end
									else
									if((r_sys_run_step==9'h3a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4451[14:0] );

									end
									else
									if((r_sys_run_step==9'h14c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5821[14:0] );

									end
									else
									if((r_sys_run_step==9'hea)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5331[14:0] );

									end
									else
									if((r_sys_run_step==9'hf0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5361[14:0] );

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4346[14:0] );

									end
									else
									if((r_sys_run_step==9'ha8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5001[14:0] );

									end
									else
									if((r_sys_run_step==9'h121)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5606[14:0] );

									end
									else
									if((r_sys_run_step==9'hd0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5201[14:0] );

									end
									else
									if((r_sys_run_step==9'h2b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4376[14:0] );

									end
									else
									if((r_sys_run_step==9'h110)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5521[14:0] );

									end
									else
									if((r_sys_run_step==9'hd3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5216[14:0] );

									end
									else
									if((r_sys_run_step==9'h4a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4531[14:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4266[14:0] );

									end
									else
									if((r_sys_run_step==9'hd8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5241[14:0] );

									end
									else
									if((r_sys_run_step==9'h9d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4946[14:0] );

									end
									else
									if((r_sys_run_step==9'h13a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5731[14:0] );

									end
									else
									if((r_sys_run_step==9'h3e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4471[14:0] );

									end
									else
									if((r_sys_run_step==9'h125)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5626[14:0] );

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4341[14:0] );

									end
									else
									if((r_sys_run_step==9'h147)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5796[14:0] );

									end
									else
									if((r_sys_run_step==9'h5b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4616[14:0] );

									end
									else
									if((r_sys_run_step==9'h22)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4331[14:0] );

									end
									else
									if((r_sys_run_step==9'h95)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4906[14:0] );

									end
									else
									if((r_sys_run_step==9'hba)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5091[14:0] );

									end
									else
									if((r_sys_run_step==9'h16e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5991[14:0] );

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4541[14:0] );

									end
									else
									if((r_sys_run_step==9'hec)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5341[14:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4164[14:0] );

									end
									else
									if((r_sys_run_step==9'h137)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5716[14:0] );

									end
									else
									if((r_sys_run_step==9'h13f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5756[14:0] );

									end
									else
									if((r_sys_run_step==9'h104)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5461[14:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4296[14:0] );

									end
									else
									if((r_sys_run_step==9'h93)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4896[14:0] );

									end
									else
									if((r_sys_run_step==9'h57)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4596[14:0] );

									end
									else
									if((r_sys_run_step==9'haa)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5011[14:0] );

									end
									else
									if((r_sys_run_step==9'h114)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5541[14:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4302[14:0] );

									end
									else
									if((r_sys_run_step==9'ha0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4961[14:0] );

									end
									else
									if((r_sys_run_step==9'h160)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5921[14:0] );

									end
									else
									if((r_sys_run_step==9'hf5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5386[14:0] );

									end
									else
									if((r_sys_run_step==9'h11f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5596[14:0] );

									end
									else
									if((r_sys_run_step==9'h41)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4486[14:0] );

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4456[14:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4140[14:0] );

									end
									else
									if((r_sys_run_step==9'hf9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5406[14:0] );

									end
									else
									if((r_sys_run_step==9'h7d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4786[14:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4206[14:0] );

									end
									else
									if((r_sys_run_step==9'h15c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5901[14:0] );

									end
									else
									if((r_sys_run_step==9'h138)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5721[14:0] );

									end
									else
									if((r_sys_run_step==9'h15e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5911[14:0] );

									end
									else
									if((r_sys_run_step==9'h139)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5726[14:0] );

									end
									else
									if((r_sys_run_step==9'h124)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5621[14:0] );

									end
									else
									if((r_sys_run_step==9'h81)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4806[14:0] );

									end
									else
									if((r_sys_run_step==9'h154)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5861[14:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4218[14:0] );

									end
									else
									if((r_sys_run_step==9'h177)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp6036[14:0] );

									end
									else
									if((r_sys_run_step==9'h174)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp6021[14:0] );

									end
									else
									if((r_sys_run_step==9'hd7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5236[14:0] );

									end
									else
									if((r_sys_run_step==9'h48)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4521[14:0] );

									end
									else
									if((r_sys_run_step==9'h76)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4751[14:0] );

									end
									else
									if((r_sys_run_step==9'hf2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5371[14:0] );

									end
									else
									if((r_sys_run_step==9'h153)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5856[14:0] );

									end
									else
									if((r_sys_run_step==9'hda)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5251[14:0] );

									end
									else
									if((r_sys_run_step==9'h36)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4431[14:0] );

									end
									else
									if((r_sys_run_step==9'h73)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4736[14:0] );

									end
									else
									if((r_sys_run_step==9'hdd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5266[14:0] );

									end
									else
									if((r_sys_run_step==9'h68)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4681[14:0] );

									end
									else
									if((r_sys_run_step==9'h8a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4851[14:0] );

									end
									else
									if((r_sys_run_step==9'hee)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5351[14:0] );

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4571[14:0] );

									end
									else
									if((r_sys_run_step==9'h159)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5886[14:0] );

									end
									else
									if((r_sys_run_step==9'h146)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5791[14:0] );

									end
									else
									if((r_sys_run_step==9'h7e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4791[14:0] );

									end
									else
									if((r_sys_run_step==9'h10e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5511[14:0] );

									end
									else
									if((r_sys_run_step==9'h175)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp6026[14:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4152[14:0] );

									end
									else
									if((r_sys_run_step==9'he7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp5316[14:0] );

									end
									else
									if((r_sys_run_step==9'h2a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4371[14:0] );

									end
									else
									if((r_sys_run_step==9'h56)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp4591[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp13;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2) || (r_sys_run_step==9'h6) || (r_sys_run_step==9'ha) || (r_sys_run_step==9'he) || (r_sys_run_step==9'h12) || (r_sys_run_step==9'h16) || (r_sys_run_step==9'h1a)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp69;

									end
									else
									if((r_sys_run_step==9'h1) || (r_sys_run_step==9'h3) || (r_sys_run_step==9'h5) || (r_sys_run_step==9'h7) || (r_sys_run_step==9'h9) || (r_sys_run_step==9'hb) || (r_sys_run_step==9'hd) || (r_sys_run_step==9'hf) || (r_sys_run_step==9'h11) || (r_sys_run_step==9'h13) || (r_sys_run_step==9'h15) || (r_sys_run_step==9'h17) || (r_sys_run_step==9'h19) || (r_sys_run_step==9'h1b)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp64;

									end
									else
									if((r_sys_run_step==9'h0) || (r_sys_run_step==9'h4) || (r_sys_run_step==9'h8) || (r_sys_run_step==9'hc) || (r_sys_run_step==9'h10) || (r_sys_run_step==9'h14) || (r_sys_run_step==9'h18)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp60;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==9'h2e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp53_float;

									end
									else
									if((r_sys_run_step==9'h28)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp71_float;

									end
									else
									if((r_sys_run_step==9'h65)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp81_float;

									end
									else
									if((r_sys_run_step==9'h76)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp31_float;

									end
									else
									if((r_sys_run_step==9'h72)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp42_float;

									end
									else
									if((r_sys_run_step==9'h35)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp32_float;

									end
									else
									if((r_sys_run_step==9'h27)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp74_float;

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp50_float;

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp20_float;

									end
									else
									if((r_sys_run_step==9'h3e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==9'h6b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp63_float;

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp80_float;

									end
									else
									if((r_sys_run_step==9'h74)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp37_float;

									end
									else
									if((r_sys_run_step==9'h2d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp56_float;

									end
									else
									if((r_sys_run_step==9'h48)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp72_float;

									end
									else
									if((r_sys_run_step==9'h73)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp39_float;

									end
									else
									if((r_sys_run_step==9'h7e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp7_float;

									end
									else
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h20)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp3470;

									end
									else
									if((r_sys_run_step==9'h55)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp33_float;

									end
									else
									if((r_sys_run_step==9'h80)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==9'h29)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp68_float;

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp64_float;

									end
									else
									if((r_sys_run_step==9'h70)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp48_float;

									end
									else
									if((r_sys_run_step==9'h22)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp89_float;

									end
									else
									if((r_sys_run_step==9'h32)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp41_float;

									end
									else
									if((r_sys_run_step==9'h46)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp79_float;

									end
									else
									if((r_sys_run_step==9'h7c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==9'h71)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp45_float;

									end
									else
									if((r_sys_run_step==9'h43)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp88_float;

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp14_float;

									end
									else
									if((r_sys_run_step==9'h44)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp84_float;

									end
									else
									if((r_sys_run_step==9'h75)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp34_float;

									end
									else
									if((r_sys_run_step==9'h5c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==9'h59)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp22_float;

									end
									else
									if((r_sys_run_step==9'h37)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp26_float;

									end
									else
									if((r_sys_run_step==9'h6f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp51_float;

									end
									else
									if((r_sys_run_step==9'h6e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp54_float;

									end
									else
									if((r_sys_run_step==9'h7a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp19_float;

									end
									else
									if((r_sys_run_step==9'h31)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp44_float;

									end
									else
									if((r_sys_run_step==9'h30)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp47_float;

									end
									else
									if((r_sys_run_step==9'h2a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp65_float;

									end
									else
									if((r_sys_run_step==9'h64)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp85_float;

									end
									else
									if((r_sys_run_step==9'h5f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==9'h56)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp30_float;

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==9'h51)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp46_float;

									end
									else
									if((r_sys_run_step==9'h67)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp76_float;

									end
									else
									if((r_sys_run_step==9'h34)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp35_float;

									end
									else
									if((r_sys_run_step==9'h7d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==9'h5b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==9'h3f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==9'h6c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp60_float;

									end
									else
									if((r_sys_run_step==9'h61)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp92_float;

									end
									else
									if((r_sys_run_step==9'h2c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp59_float;

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==9'h41)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp93_float;

									end
									else
									if((r_sys_run_step==9'h7b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==9'h4a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp67_float;

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp36_float;

									end
									else
									if((r_sys_run_step==9'h38)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp23_float;

									end
									else
									if((r_sys_run_step==9'h26)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp77_float;

									end
									else
									if((r_sys_run_step==9'h6a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp66_float;

									end
									else
									if((r_sys_run_step==9'h6d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp57_float;

									end
									else
									if((r_sys_run_step==9'h68)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp73_float;

									end
									else
									if((r_sys_run_step==9'h49)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp69_float;

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp61_float;

									end
									else
									if((r_sys_run_step==9'h45)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp82_float;

									end
									else
									if((r_sys_run_step==9'h5e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp83_float;

									end
									else
									if((r_sys_run_step==9'h62)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp91_float;

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp43_float;

									end
									else
									if((r_sys_run_step==9'h53)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp40_float;

									end
									else
									if((r_sys_run_step==9'h69)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp70_float;

									end
									else
									if((r_sys_run_step==9'h58)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp25_float;

									end
									else
									if((r_sys_run_step==9'h42)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp90_float;

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp55_float;

									end
									else
									if((r_sys_run_step==9'h50)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp49_float;

									end
									else
									if((r_sys_run_step==9'h7f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==9'h79)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp21_float;

									end
									else
									if((r_sys_run_step==9'h78)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp24_float;

									end
									else
									if((r_sys_run_step==9'h63)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp87_float;

									end
									else
									if((r_sys_run_step==9'h57)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp27_float;

									end
									else
									if((r_sys_run_step==9'h4f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp52_float;

									end
									else
									if((r_sys_run_step==9'h2b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp62_float;

									end
									else
									if((r_sys_run_step==9'h23)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp86_float;

									end
									else
									if((r_sys_run_step==9'h5a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp18_float;

									end
									else
									if((r_sys_run_step==9'h33)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp38_float;

									end
									else
									if((r_sys_run_step==9'h60)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==9'h21) || (r_sys_run_step==9'h40)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp94_float;

									end
									else
									if((r_sys_run_step==9'h3a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==9'h36)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp29_float;

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp75_float;

									end
									else
									if((r_sys_run_step==9'h4d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp58_float;

									end
									else
									if((r_sys_run_step==9'h77)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp28_float;

									end
									else
									if((r_sys_run_step==9'h66)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp78_float;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h82)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp336_float;

									end
									else
									if((r_sys_run_step==9'h174)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp116_float;

									end
									else
									if((r_sys_run_step==9'h140)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp330_float;

									end
									else
									if((r_sys_run_step==9'h16c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp204_float;

									end
									else
									if((r_sys_run_step==9'h12c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp196_float;

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp31_float;

									end
									else
									if((r_sys_run_step==9'h4a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp245_float;

									end
									else
									if((r_sys_run_step==9'h11c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp32_float;

									end
									else
									if((r_sys_run_step==9'h65)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp296_float;

									end
									else
									if((r_sys_run_step==9'h17e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==9'h159)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp63_float;

									end
									else
									if((r_sys_run_step==9'h38)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp80_float;

									end
									else
									if((r_sys_run_step==9'h14c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp205_float;

									end
									else
									if((r_sys_run_step==9'h134)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp112_float;

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp203_float;

									end
									else
									if((r_sys_run_step==9'hae)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp193_float;

									end
									else
									if((r_sys_run_step==9'hdc)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp37_float;

									end
									else
									if((r_sys_run_step==9'h6e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp199_float;

									end
									else
									if((r_sys_run_step==9'ha7)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp266_float;

									end
									else
									if((r_sys_run_step==9'h120)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp331_float;

									end
									else
									if((r_sys_run_step==9'h108)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp257_float;

									end
									else
									if((r_sys_run_step==9'h104)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp302_float;

									end
									else
									if((r_sys_run_step==9'h103)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp312_float;

									end
									else
									if((r_sys_run_step==9'h17a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp45_float;

									end
									else
									if((r_sys_run_step==9'h173)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp128_float;

									end
									else
									if((r_sys_run_step==9'h98)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp88_float;

									end
									else
									if((r_sys_run_step==9'hfe)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp14_float;

									end
									else
									if((r_sys_run_step==9'h109)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp240_float;

									end
									else
									if((r_sys_run_step==9'h7d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp34_float;

									end
									else
									if((r_sys_run_step==9'h48)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp263_float;

									end
									else
									if((r_sys_run_step==9'h15f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp339_float;

									end
									else
									if((r_sys_run_step==9'h13d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==9'h131)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp141_float;

									end
									else
									if((r_sys_run_step==9'h46)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp287_float;

									end
									else
									if((r_sys_run_step==9'hdd)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp26_float;

									end
									else
									if((r_sys_run_step==9'h34)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp129_float;

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp184_float;

									end
									else
									if((r_sys_run_step==9'hee)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp188_float;

									end
									else
									if((r_sys_run_step==9'h84)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp306_float;

									end
									else
									if((r_sys_run_step==9'h12b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp207_float;

									end
									else
									if((r_sys_run_step==9'h135)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp101_float;

									end
									else
									if((r_sys_run_step==9'he6)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp276_float;

									end
									else
									if((r_sys_run_step==9'h127)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp260_float;

									end
									else
									if((r_sys_run_step==9'h106)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp282_float;

									end
									else
									if((r_sys_run_step==9'h66)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp285_float;

									end
									else
									if((r_sys_run_step==9'hbb)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp46_float;

									end
									else
									if((r_sys_run_step==9'h138)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp76_float;

									end
									else
									if((r_sys_run_step==9'h91)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp168_float;

									end
									else
									if((r_sys_run_step==9'hb1)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp157_float;

									end
									else
									if((r_sys_run_step==9'h132)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp130_float;

									end
									else
									if((r_sys_run_step==9'h11e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==9'h5b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp59_float;

									end
									else
									if((r_sys_run_step==9'h44)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp307_float;

									end
									else
									if((r_sys_run_step==9'ha8)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp255_float;

									end
									else
									if((r_sys_run_step==9'h76)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp114_float;

									end
									else
									if((r_sys_run_step==9'h8c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp219_float;

									end
									else
									if((r_sys_run_step==9'hc1)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp334_float;

									end
									else
									if((r_sys_run_step==9'hf6)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp97_float;

									end
									else
									if((r_sys_run_step==9'h147)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp259_float;

									end
									else
									if((r_sys_run_step==9'h11d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp23_float;

									end
									else
									if((r_sys_run_step==9'h83)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp326_float;

									end
									else
									if((r_sys_run_step==9'h8d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp212_float;

									end
									else
									if((r_sys_run_step==9'hc7)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp264_float;

									end
									else
									if((r_sys_run_step==9'h100)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp338_float;

									end
									else
									if((r_sys_run_step==9'h178)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp66_float;

									end
									else
									if((r_sys_run_step==9'h16b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp216_float;

									end
									else
									if((r_sys_run_step==9'h50)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp181_float;

									end
									else
									if((r_sys_run_step==9'h8e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp197_float;

									end
									else
									if((r_sys_run_step==9'hef)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp178_float;

									end
									else
									if((r_sys_run_step==9'h49)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp254_float;

									end
									else
									if((r_sys_run_step==9'h8f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp190_float;

									end
									else
									if((r_sys_run_step==9'hf7)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp83_float;

									end
									else
									if((r_sys_run_step==9'h170)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp160_float;

									end
									else
									if((r_sys_run_step==9'h117)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp91_float;

									end
									else
									if((r_sys_run_step==9'h126)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp270_float;

									end
									else
									if((r_sys_run_step==9'h172)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp138_float;

									end
									else
									if((r_sys_run_step==9'hb9)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp70_float;

									end
									else
									if((r_sys_run_step==9'h12d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp185_float;

									end
									else
									if((r_sys_run_step==9'hfb)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp49_float;

									end
									else
									if((r_sys_run_step==9'h13c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp24_float;

									end
									else
									if((r_sys_run_step==9'hd4)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp125_float;

									end
									else
									if((r_sys_run_step==9'hf3)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp134_float;

									end
									else
									if((r_sys_run_step==9'h23)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp316_float;

									end
									else
									if((r_sys_run_step==9'hc5)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp284_float;

									end
									else
									if((r_sys_run_step==9'hd1)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp158_float;

									end
									else
									if((r_sys_run_step==9'h157)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp86_float;

									end
									else
									if((r_sys_run_step==9'h3e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp18_float;

									end
									else
									if((r_sys_run_step==9'h6f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp187_float;

									end
									else
									if((r_sys_run_step==9'hf5)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp110_float;

									end
									else
									if((r_sys_run_step==9'h156)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp94_float;

									end
									else
									if((r_sys_run_step==9'h60)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==9'h143)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp300_float;

									end
									else
									if((r_sys_run_step==9'h61)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp346_float;

									end
									else
									if((r_sys_run_step==9'h53)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp148_float;

									end
									else
									if((r_sys_run_step==9'hb4)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp127_float;

									end
									else
									if((r_sys_run_step==9'h7b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp58_float;

									end
									else
									if((r_sys_run_step==9'he4)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp303_float;

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp78_float;

									end
									else
									if((r_sys_run_step==9'h9f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==9'h6c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp221_float;

									end
									else
									if((r_sys_run_step==9'h2a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp239_float;

									end
									else
									if((r_sys_run_step==9'h96)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp111_float;

									end
									else
									if((r_sys_run_step==9'h141)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp320_float;

									end
									else
									if((r_sys_run_step==9'h9e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp20_float;

									end
									else
									if((r_sys_run_step==9'h16d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp194_float;

									end
									else
									if((r_sys_run_step==9'h94)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp131_float;

									end
									else
									if((r_sys_run_step==9'h85)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp297_float;

									end
									else
									if((r_sys_run_step==9'h160)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp329_float;

									end
									else
									if((r_sys_run_step==9'hc2)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp324_float;

									end
									else
									if((r_sys_run_step==9'h13b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp39_float;

									end
									else
									if((r_sys_run_step==9'hf4)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp122_float;

									end
									else
									if((r_sys_run_step==9'hbf)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==9'h80)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==9'h9a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp64_float;

									end
									else
									if((r_sys_run_step==9'hd9)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp68_float;

									end
									else
									if((r_sys_run_step==9'h56)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp109_float;

									end
									else
									if((r_sys_run_step==9'hb7)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp89_float;

									end
									else
									if((r_sys_run_step==9'hf1)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp156_float;

									end
									else
									if((r_sys_run_step==9'hca)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp234_float;

									end
									else
									if((r_sys_run_step==9'h145)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp280_float;

									end
									else
									if((r_sys_run_step==9'h67)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp277_float;

									end
									else
									if((r_sys_run_step==9'h74)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp137_float;

									end
									else
									if((r_sys_run_step==9'h27)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp272_float;

									end
									else
									if((r_sys_run_step==9'h17c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp22_float;

									end
									else
									if((r_sys_run_step==9'h15a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp51_float;

									end
									else
									if((r_sys_run_step==9'h33)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp140_float;

									end
									else
									if((r_sys_run_step==9'h21) || (r_sys_run_step==9'h40)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp348_float;

									end
									else
									if((r_sys_run_step==9'hba)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp54_float;

									end
									else
									if((r_sys_run_step==9'hac)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp215_float;

									end
									else
									if((r_sys_run_step==9'h5c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp47_float;

									end
									else
									if((r_sys_run_step==9'h8a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp241_float;

									end
									else
									if((r_sys_run_step==9'ha0)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp344_float;

									end
									else
									if((r_sys_run_step==9'h171)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp150_float;

									end
									else
									if((r_sys_run_step==9'h133)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp119_float;

									end
									else
									if((r_sys_run_step==9'h17d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==9'h130)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp152_float;

									end
									else
									if((r_sys_run_step==9'h105)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp292_float;

									end
									else
									if((r_sys_run_step==9'he0)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp342_float;

									end
									else
									if((r_sys_run_step==9'h26)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp283_float;

									end
									else
									if((r_sys_run_step==9'h162)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp309_float;

									end
									else
									if((r_sys_run_step==9'h43)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp318_float;

									end
									else
									if((r_sys_run_step==9'h111)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp154_float;

									end
									else
									if((r_sys_run_step==9'hd6)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp99_float;

									end
									else
									if((r_sys_run_step==9'h92)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp153_float;

									end
									else
									if((r_sys_run_step==9'h36)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp107_float;

									end
									else
									if((r_sys_run_step==9'h4d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp214_float;

									end
									else
									if((r_sys_run_step==9'h10f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp176_float;

									end
									else
									if((r_sys_run_step==9'hdf)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==9'he5)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp293_float;

									end
									else
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h20)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp4142;

									end
									else
									if((r_sys_run_step==9'hd7)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp93_float;

									end
									else
									if((r_sys_run_step==9'h7f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==9'h32)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp151_float;

									end
									else
									if((r_sys_run_step==9'h10b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp220_float;

									end
									else
									if((r_sys_run_step==9'h73)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp143_float;

									end
									else
									if((r_sys_run_step==9'h11a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp57_float;

									end
									else
									if((r_sys_run_step==9'h10a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp229_float;

									end
									else
									if((r_sys_run_step==9'h5a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp69_float;

									end
									else
									if((r_sys_run_step==9'h78)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp82_float;

									end
									else
									if((r_sys_run_step==9'h13e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==9'hcb)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp224_float;

									end
									else
									if((r_sys_run_step==9'hab)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp223_float;

									end
									else
									if((r_sys_run_step==9'h62)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp337_float;

									end
									else
									if((r_sys_run_step==9'he8)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp251_float;

									end
									else
									if((r_sys_run_step==9'h165)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp279_float;

									end
									else
									if((r_sys_run_step==9'hc6)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp273_float;

									end
									else
									if((r_sys_run_step==9'ha4)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp295_float;

									end
									else
									if((r_sys_run_step==9'h155)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp106_float;

									end
									else
									if((r_sys_run_step==9'h12f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp163_float;

									end
									else
									if((r_sys_run_step==9'h166)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp268_float;

									end
									else
									if((r_sys_run_step==9'h16a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp226_float;

									end
									else
									if((r_sys_run_step==9'haf)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp179_float;

									end
									else
									if((r_sys_run_step==9'hfd)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp27_float;

									end
									else
									if((r_sys_run_step==9'h6b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp230_float;

									end
									else
									if((r_sys_run_step==9'h125)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp281_float;

									end
									else
									if((r_sys_run_step==9'ha2)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp325_float;

									end
									else
									if((r_sys_run_step==9'he7)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp262_float;

									end
									else
									if((r_sys_run_step==9'h142)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp310_float;

									end
									else
									if((r_sys_run_step==9'h81)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp345_float;

									end
									else
									if((r_sys_run_step==9'hbe)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==9'h45)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp298_float;

									end
									else
									if((r_sys_run_step==9'h16f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp172_float;

									end
									else
									if((r_sys_run_step==9'haa)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp236_float;

									end
									else
									if((r_sys_run_step==9'h59)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp75_float;

									end
									else
									if((r_sys_run_step==9'ha5)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp286_float;

									end
									else
									if((r_sys_run_step==9'h101)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp332_float;

									end
									else
									if((r_sys_run_step==9'h10d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp198_float;

									end
									else
									if((r_sys_run_step==9'h7e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp28_float;

									end
									else
									if((r_sys_run_step==9'h9b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp53_float;

									end
									else
									if((r_sys_run_step==9'h13f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp340_float;

									end
									else
									if((r_sys_run_step==9'hcd)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp202_float;

									end
									else
									if((r_sys_run_step==9'h14f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp167_float;

									end
									else
									if((r_sys_run_step==9'hb2)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp149_float;

									end
									else
									if((r_sys_run_step==9'hec)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp210_float;

									end
									else
									if((r_sys_run_step==9'h95)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp121_float;

									end
									else
									if((r_sys_run_step==9'hf8)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp74_float;

									end
									else
									if((r_sys_run_step==9'hbc)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp42_float;

									end
									else
									if((r_sys_run_step==9'hd0)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp169_float;

									end
									else
									if((r_sys_run_step==9'hc4)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp304_float;

									end
									else
									if((r_sys_run_step==9'h136)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp95_float;

									end
									else
									if((r_sys_run_step==9'h179)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp56_float;

									end
									else
									if((r_sys_run_step==9'hc0)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp343_float;

									end
									else
									if((r_sys_run_step==9'h150)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp161_float;

									end
									else
									if((r_sys_run_step==9'h128)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp249_float;

									end
									else
									if((r_sys_run_step==9'ha1)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp335_float;

									end
									else
									if((r_sys_run_step==9'hdb)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp48_float;

									end
									else
									if((r_sys_run_step==9'h9c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp41_float;

									end
									else
									if((r_sys_run_step==9'hf0)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp166_float;

									end
									else
									if((r_sys_run_step==9'h15d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==9'h11f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp341_float;

									end
									else
									if((r_sys_run_step==9'h75)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp126_float;

									end
									else
									if((r_sys_run_step==9'h118)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp84_float;

									end
									else
									if((r_sys_run_step==9'h113)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp132_float;

									end
									else
									if((r_sys_run_step==9'h29)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp250_float;

									end
									else
									if((r_sys_run_step==9'h70)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp177_float;

									end
									else
									if((r_sys_run_step==9'h114)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp120_float;

									end
									else
									if((r_sys_run_step==9'he9)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp242_float;

									end
									else
									if((r_sys_run_step==9'h7a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp65_float;

									end
									else
									if((r_sys_run_step==9'hce)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp191_float;

									end
									else
									if((r_sys_run_step==9'he3)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp313_float;

									end
									else
									if((r_sys_run_step==9'h163)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp299_float;

									end
									else
									if((r_sys_run_step==9'h15e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==9'h99)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp85_float;

									end
									else
									if((r_sys_run_step==9'had)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp201_float;

									end
									else
									if((r_sys_run_step==9'hb5)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp115_float;

									end
									else
									if((r_sys_run_step==9'h41)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp347_float;

									end
									else
									if((r_sys_run_step==9'h124)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp291_float;

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp294_float;

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp225_float;

									end
									else
									if((r_sys_run_step==9'h42)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp328_float;

									end
									else
									if((r_sys_run_step==9'h9d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp35_float;

									end
									else
									if((r_sys_run_step==9'hc8)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp253_float;

									end
									else
									if((r_sys_run_step==9'hde)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==9'h58)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp92_float;

									end
									else
									if((r_sys_run_step==9'h3a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp60_float;

									end
									else
									if((r_sys_run_step==9'h51)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp170_float;

									end
									else
									if((r_sys_run_step==9'h37)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp96_float;

									end
									else
									if((r_sys_run_step==9'hc9)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp244_float;

									end
									else
									if((r_sys_run_step==9'h3f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==9'h158)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp67_float;

									end
									else
									if((r_sys_run_step==9'h31)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp162_float;

									end
									else
									if((r_sys_run_step==9'hb3)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp135_float;

									end
									else
									if((r_sys_run_step==9'hd2)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp147_float;

									end
									else
									if((r_sys_run_step==9'h16e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp182_float;

									end
									else
									if((r_sys_run_step==9'hea)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp231_float;

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp305_float;

									end
									else
									if((r_sys_run_step==9'h72)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp155_float;

									end
									else
									if((r_sys_run_step==9'hcf)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp180_float;

									end
									else
									if((r_sys_run_step==9'h175)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp105_float;

									end
									else
									if((r_sys_run_step==9'hfa)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp61_float;

									end
									else
									if((r_sys_run_step==9'h6a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp243_float;

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp274_float;

									end
									else
									if((r_sys_run_step==9'h68)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp265_float;

									end
									else
									if((r_sys_run_step==9'h176)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp90_float;

									end
									else
									if((r_sys_run_step==9'hc3)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp314_float;

									end
									else
									if((r_sys_run_step==9'h5e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp21_float;

									end
									else
									if((r_sys_run_step==9'h89)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp252_float;

									end
									else
									if((r_sys_run_step==9'h154)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp117_float;

									end
									else
									if((r_sys_run_step==9'hb0)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp171_float;

									end
									else
									if((r_sys_run_step==9'h177)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp87_float;

									end
									else
									if((r_sys_run_step==9'h139)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp62_float;

									end
									else
									if((r_sys_run_step==9'h169)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp237_float;

									end
									else
									if((r_sys_run_step==9'ha9)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp246_float;

									end
									else
									if((r_sys_run_step==9'hb6)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp103_float;

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp159_float;

									end
									else
									if((r_sys_run_step==9'h12e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp174_float;

									end
									else
									if((r_sys_run_step==9'h115)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp108_float;

									end
									else
									if((r_sys_run_step==9'hbd)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp29_float;

									end
									else
									if((r_sys_run_step==9'h2b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp228_float;

									end
									else
									if((r_sys_run_step==9'h164)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp289_float;

									end
									else
									if((r_sys_run_step==9'hf9)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp71_float;

									end
									else
									if((r_sys_run_step==9'h121)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp321_float;

									end
									else
									if((r_sys_run_step==9'h64)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp308_float;

									end
									else
									if((r_sys_run_step==9'h137)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp81_float;

									end
									else
									if((r_sys_run_step==9'h69)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp256_float;

									end
									else
									if((r_sys_run_step==9'h148)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp248_float;

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp133_float;

									end
									else
									if((r_sys_run_step==9'h13a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp50_float;

									end
									else
									if((r_sys_run_step==9'h2d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp206_float;

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp235_float;

									end
									else
									if((r_sys_run_step==9'h107)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp271_float;

									end
									else
									if((r_sys_run_step==9'h77)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp102_float;

									end
									else
									if((r_sys_run_step==9'h153)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp123_float;

									end
									else
									if((r_sys_run_step==9'h79)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp72_float;

									end
									else
									if((r_sys_run_step==9'h167)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp258_float;

									end
									else
									if((r_sys_run_step==9'h17b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp33_float;

									end
									else
									if((r_sys_run_step==9'h14b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp211_float;

									end
									else
									if((r_sys_run_step==9'h116)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp100_float;

									end
									else
									if((r_sys_run_step==9'h63)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp317_float;

									end
									else
									if((r_sys_run_step==9'hd8)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp79_float;

									end
									else
									if((r_sys_run_step==9'ha6)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp275_float;

									end
									else
									if((r_sys_run_step==9'hd5)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp113_float;

									end
									else
									if((r_sys_run_step==9'h10c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp208_float;

									end
									else
									if((r_sys_run_step==9'h97)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp104_float;

									end
									else
									if((r_sys_run_step==9'h110)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp164_float;

									end
									else
									if((r_sys_run_step==9'h123)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp301_float;

									end
									else
									if((r_sys_run_step==9'hed)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp200_float;

									end
									else
									if((r_sys_run_step==9'h5f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp19_float;

									end
									else
									if((r_sys_run_step==9'h12a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp218_float;

									end
									else
									if((r_sys_run_step==9'h11b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp44_float;

									end
									else
									if((r_sys_run_step==9'h55)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp124_float;

									end
									else
									if((r_sys_run_step==9'h22)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp327_float;

									end
									else
									if((r_sys_run_step==9'h146)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp269_float;

									end
									else
									if((r_sys_run_step==9'hd3)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp136_float;

									end
									else
									if((r_sys_run_step==9'h5d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp30_float;

									end
									else
									if((r_sys_run_step==9'h161)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp319_float;

									end
									else
									if((r_sys_run_step==9'h152)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp139_float;

									end
									else
									if((r_sys_run_step==9'h168)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp247_float;

									end
									else
									if((r_sys_run_step==9'h71)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp165_float;

									end
									else
									if((r_sys_run_step==9'h57)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp98_float;

									end
									else
									if((r_sys_run_step==9'h35)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp118_float;

									end
									else
									if((r_sys_run_step==9'h112)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp142_float;

									end
									else
									if((r_sys_run_step==9'hfc)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp36_float;

									end
									else
									if((r_sys_run_step==9'h119)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp77_float;

									end
									else
									if((r_sys_run_step==9'h28)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp261_float;

									end
									else
									if((r_sys_run_step==9'h149)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp238_float;

									end
									else
									if((r_sys_run_step==9'h87)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp278_float;

									end
									else
									if((r_sys_run_step==9'hb8)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp73_float;

									end
									else
									if((r_sys_run_step==9'h102)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp322_float;

									end
									else
									if((r_sys_run_step==9'h88)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp267_float;

									end
									else
									if((r_sys_run_step==9'h10e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp186_float;

									end
									else
									if((r_sys_run_step==9'h14d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp189_float;

									end
									else
									if((r_sys_run_step==9'h4f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp192_float;

									end
									else
									if((r_sys_run_step==9'he1)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp333_float;

									end
									else
									if((r_sys_run_step==9'h90)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp175_float;

									end
									else
									if((r_sys_run_step==9'h14a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp227_float;

									end
									else
									if((r_sys_run_step==9'heb)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp222_float;

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp43_float;

									end
									else
									if((r_sys_run_step==9'h7c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp40_float;

									end
									else
									if((r_sys_run_step==9'h15c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp25_float;

									end
									else
									if((r_sys_run_step==9'h144)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp290_float;

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp55_float;

									end
									else
									if((r_sys_run_step==9'h30)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp173_float;

									end
									else
									if((r_sys_run_step==9'h8b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp232_float;

									end
									else
									if((r_sys_run_step==9'h129)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp233_float;

									end
									else
									if((r_sys_run_step==9'h151)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp145_float;

									end
									else
									if((r_sys_run_step==9'hff)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==9'hda)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp52_float;

									end
									else
									if((r_sys_run_step==9'h14e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp183_float;

									end
									else
									if((r_sys_run_step==9'h15b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp38_float;

									end
									else
									if((r_sys_run_step==9'h2c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp217_float;

									end
									else
									if((r_sys_run_step==9'h93)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp146_float;

									end
									else
									if((r_sys_run_step==9'h6d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp209_float;

									end
									else
									if((r_sys_run_step==9'h86)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp288_float;

									end
									else
									if((r_sys_run_step==9'he2)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp323_float;

									end
									else
									if((r_sys_run_step==9'h2e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp195_float;

									end
									else
									if((r_sys_run_step==9'hcc)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp213_float;

									end
									else
									if((r_sys_run_step==9'hf2)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp144_float;

									end
									else
									if((r_sys_run_step==9'h122)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp311_float;

									end
									else
									if((r_sys_run_step==9'ha3)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp315_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1b)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h86)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h194)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h80)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h17e)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h35: begin
							r_fld_u_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_17 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_17 <= w_sys_tmp5;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_17 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h88)) begin
										r_run_k_17 <= w_sys_tmp1025;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_17 <= w_sys_tmp1026;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h196)) begin
										r_run_k_17 <= w_sys_tmp3461;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_17 <= w_sys_tmp3462;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h80)) begin
										r_run_k_17 <= w_sys_tmp4133;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_17 <= w_sys_tmp4134;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h17e)) begin
										r_run_k_17 <= w_sys_tmp6075;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_j_18 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6)) begin
										r_run_j_18 <= w_sys_tmp14;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_j_18 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0) || (r_sys_run_step==9'h4) || (r_sys_run_step==9'h8) || (r_sys_run_step==9'hc) || (r_sys_run_step==9'h10) || (r_sys_run_step==9'h14) || (r_sys_run_step==9'h18)) begin
										r_run_j_18 <= w_sys_tmp78;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_n_19 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_n_19 <= w_sys_tmp53;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_mx_20 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_my_21 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_nlast_22 <= w_sys_intOne;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy0_j_23 <= r_run_j_18;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3) || (r_sys_run_step==9'h7) || (r_sys_run_step==9'hb) || (r_sys_run_step==9'hf) || (r_sys_run_step==9'h13) || (r_sys_run_step==9'h17) || (r_sys_run_step==9'h1b)) begin
										r_run_copy0_j_23 <= w_sys_tmp75;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy1_j_24 <= r_run_j_18;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2) || (r_sys_run_step==9'h6) || (r_sys_run_step==9'ha) || (r_sys_run_step==9'he) || (r_sys_run_step==9'h12) || (r_sys_run_step==9'h16) || (r_sys_run_step==9'h1a)) begin
										r_run_copy1_j_24 <= w_sys_tmp76;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy2_j_25 <= r_run_j_18;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1) || (r_sys_run_step==9'h5) || (r_sys_run_step==9'h9) || (r_sys_run_step==9'hd) || (r_sys_run_step==9'h11) || (r_sys_run_step==9'h15) || (r_sys_run_step==9'h19)) begin
										r_run_copy2_j_25 <= w_sys_tmp77;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h7: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub09_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub09_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc5)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2202[14:0] );

									end
									else
									if((r_sys_run_step==9'hc4)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2196[14:0] );

									end
									else
									if((r_sys_run_step==9'haf)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2070[14:0] );

									end
									else
									if((r_sys_run_step==9'hc1)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2178[14:0] );

									end
									else
									if((r_sys_run_step==9'hb5)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2106[14:0] );

									end
									else
									if((r_sys_run_step==9'hba)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2136[14:0] );

									end
									else
									if((r_sys_run_step==9'hb6)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2112[14:0] );

									end
									else
									if((r_sys_run_step==9'hab)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2034[14:0] );

									end
									else
									if((r_sys_run_step==9'hc9)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2226[14:0] );

									end
									else
									if((r_sys_run_step==9'hc6)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2208[14:0] );

									end
									else
									if((r_sys_run_step==9'hb7)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2118[14:0] );

									end
									else
									if((r_sys_run_step==9'hc3)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2190[14:0] );

									end
									else
									if((r_sys_run_step==9'hc8)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2220[14:0] );

									end
									else
									if((r_sys_run_step==9'hc7)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2214[14:0] );

									end
									else
									if((r_sys_run_step==9'hb9)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2130[14:0] );

									end
									else
									if((r_sys_run_step==9'hac)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2052[14:0] );

									end
									else
									if((r_sys_run_step==9'hcb)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2238[14:0] );

									end
									else
									if((r_sys_run_step==9'hb2)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2088[14:0] );

									end
									else
									if((r_sys_run_step==9'hc0)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2172[14:0] );

									end
									else
									if((r_sys_run_step==9'hc2)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2184[14:0] );

									end
									else
									if((r_sys_run_step==9'hbc)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2148[14:0] );

									end
									else
									if((r_sys_run_step==9'hb8)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2124[14:0] );

									end
									else
									if((r_sys_run_step==9'hbe)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2160[14:0] );

									end
									else
									if((r_sys_run_step==9'hae)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2064[14:0] );

									end
									else
									if((r_sys_run_step==9'hb0)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2076[14:0] );

									end
									else
									if((r_sys_run_step==9'hbb)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2142[14:0] );

									end
									else
									if((r_sys_run_step==9'hbf)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2166[14:0] );

									end
									else
									if((r_sys_run_step==9'hca)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2232[14:0] );

									end
									else
									if((r_sys_run_step==9'had)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2058[14:0] );

									end
									else
									if((r_sys_run_step==9'haa)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2028[14:0] );

									end
									else
									if((r_sys_run_step==9'hb4)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2100[14:0] );

									end
									else
									if((r_sys_run_step==9'hb1)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2082[14:0] );

									end
									else
									if((r_sys_run_step==9'hb3)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2094[14:0] );

									end
									else
									if((r_sys_run_step==9'hbd)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp2154[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'haa<=r_sys_run_step && r_sys_run_step<=9'hcb)) begin
										r_sub09_u_datain <= w_sys_tmp1034;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'haa<=r_sys_run_step && r_sys_run_step<=9'hcb)) begin
										r_sub09_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub09_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5046[14:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4981[14:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5051[14:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5026[14:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4996[14:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5011[14:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4991[14:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5066[14:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5081[14:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4961[14:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5041[14:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5056[14:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5116[14:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5016[14:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5101[14:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5021[14:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5086[14:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5106[14:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5111[14:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5001[14:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5031[14:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4986[14:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4966[14:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5076[14:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5071[14:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4976[14:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5091[14:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5061[14:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4971[14:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5036[14:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5006[14:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp5096[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1f)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub09_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub08_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub08_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha1)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1986[14:0] );

									end
									else
									if((r_sys_run_step==9'h89)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1842[14:0] );

									end
									else
									if((r_sys_run_step==9'h96)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1920[14:0] );

									end
									else
									if((r_sys_run_step==9'h8d)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1866[14:0] );

									end
									else
									if((r_sys_run_step==9'h99)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1938[14:0] );

									end
									else
									if((r_sys_run_step==9'h94)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1908[14:0] );

									end
									else
									if((r_sys_run_step==9'ha9)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp2034[14:0] );

									end
									else
									if((r_sys_run_step==9'h95)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1914[14:0] );

									end
									else
									if((r_sys_run_step==9'h9b)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1950[14:0] );

									end
									else
									if((r_sys_run_step==9'h8a)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1848[14:0] );

									end
									else
									if((r_sys_run_step==9'ha2)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1992[14:0] );

									end
									else
									if((r_sys_run_step==9'ha5)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp2010[14:0] );

									end
									else
									if((r_sys_run_step==9'h98)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1932[14:0] );

									end
									else
									if((r_sys_run_step==9'h9c)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1956[14:0] );

									end
									else
									if((r_sys_run_step==9'h8c)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1860[14:0] );

									end
									else
									if((r_sys_run_step==9'ha6)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp2016[14:0] );

									end
									else
									if((r_sys_run_step==9'h9d)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1962[14:0] );

									end
									else
									if((r_sys_run_step==9'ha0)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1980[14:0] );

									end
									else
									if((r_sys_run_step==9'h91)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1890[14:0] );

									end
									else
									if((r_sys_run_step==9'h8e)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1872[14:0] );

									end
									else
									if((r_sys_run_step==9'h9f)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1974[14:0] );

									end
									else
									if((r_sys_run_step==9'ha3)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1998[14:0] );

									end
									else
									if((r_sys_run_step==9'h93)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1902[14:0] );

									end
									else
									if((r_sys_run_step==9'ha4)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp2004[14:0] );

									end
									else
									if((r_sys_run_step==9'h92)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1896[14:0] );

									end
									else
									if((r_sys_run_step==9'ha7)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp2022[14:0] );

									end
									else
									if((r_sys_run_step==9'h97)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1926[14:0] );

									end
									else
									if((r_sys_run_step==9'h8f)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1878[14:0] );

									end
									else
									if((r_sys_run_step==9'ha8)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp2028[14:0] );

									end
									else
									if((r_sys_run_step==9'h8b)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1854[14:0] );

									end
									else
									if((r_sys_run_step==9'h9e)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1968[14:0] );

									end
									else
									if((r_sys_run_step==9'h90)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1884[14:0] );

									end
									else
									if((r_sys_run_step==9'h9a)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp1944[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h89<=r_sys_run_step && r_sys_run_step<=9'ha9)) begin
										r_sub08_u_datain <= w_sys_tmp1034;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h89<=r_sys_run_step && r_sys_run_step<=9'ha9)) begin
										r_sub08_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub08_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1e)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4956[14:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4866[14:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4916[14:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4896[14:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4826[14:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4876[14:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4871[14:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4846[14:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4811[14:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4901[14:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4926[14:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4841[14:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4821[14:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4941[14:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4806[14:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4861[14:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4911[14:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4836[14:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4936[14:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4891[14:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4881[14:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4946[14:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4931[14:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4851[14:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4816[14:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4906[14:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4831[14:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4951[14:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4856[14:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4886[14:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4921[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1e)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub08_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h10: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub12_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub12_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11a)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2712[14:0] );

									end
									else
									if((r_sys_run_step==9'h130)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2844[14:0] );

									end
									else
									if((r_sys_run_step==9'h11b)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2718[14:0] );

									end
									else
									if((r_sys_run_step==9'h112)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2664[14:0] );

									end
									else
									if((r_sys_run_step==9'h111)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2658[14:0] );

									end
									else
									if((r_sys_run_step==9'h12d)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2826[14:0] );

									end
									else
									if((r_sys_run_step==9'h125)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2778[14:0] );

									end
									else
									if((r_sys_run_step==9'h12a)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2808[14:0] );

									end
									else
									if((r_sys_run_step==9'h127)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2790[14:0] );

									end
									else
									if((r_sys_run_step==9'h116)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2688[14:0] );

									end
									else
									if((r_sys_run_step==9'h113)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2670[14:0] );

									end
									else
									if((r_sys_run_step==9'h123)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2766[14:0] );

									end
									else
									if((r_sys_run_step==9'h11f)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2742[14:0] );

									end
									else
									if((r_sys_run_step==9'h126)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2784[14:0] );

									end
									else
									if((r_sys_run_step==9'h121)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2754[14:0] );

									end
									else
									if((r_sys_run_step==9'h114)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2676[14:0] );

									end
									else
									if((r_sys_run_step==9'h119)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2706[14:0] );

									end
									else
									if((r_sys_run_step==9'h12b)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2814[14:0] );

									end
									else
									if((r_sys_run_step==9'h124)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2772[14:0] );

									end
									else
									if((r_sys_run_step==9'h12c)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2820[14:0] );

									end
									else
									if((r_sys_run_step==9'h110)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2652[14:0] );

									end
									else
									if((r_sys_run_step==9'h120)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2748[14:0] );

									end
									else
									if((r_sys_run_step==9'h12e)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2832[14:0] );

									end
									else
									if((r_sys_run_step==9'h11c)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2724[14:0] );

									end
									else
									if((r_sys_run_step==9'h129)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2802[14:0] );

									end
									else
									if((r_sys_run_step==9'h118)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2700[14:0] );

									end
									else
									if((r_sys_run_step==9'h115)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2682[14:0] );

									end
									else
									if((r_sys_run_step==9'h122)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2760[14:0] );

									end
									else
									if((r_sys_run_step==9'h12f)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2838[14:0] );

									end
									else
									if((r_sys_run_step==9'h128)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2796[14:0] );

									end
									else
									if((r_sys_run_step==9'h117)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2694[14:0] );

									end
									else
									if((r_sys_run_step==9'h11d)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2730[14:0] );

									end
									else
									if((r_sys_run_step==9'h11e)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp2736[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h110<=r_sys_run_step && r_sys_run_step<=9'h130)) begin
										r_sub12_u_datain <= w_sys_tmp1034;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h110<=r_sys_run_step && r_sys_run_step<=9'h130)) begin
										r_sub12_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub12_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5481[14:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5471[14:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5441[14:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5556[14:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5576[14:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5541[14:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5581[14:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5476[14:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5586[14:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5531[14:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5526[14:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5561[14:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5456[14:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5551[14:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5506[14:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5466[14:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5546[14:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5536[14:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5496[14:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5491[14:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5521[14:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5451[14:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5571[14:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5591[14:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5566[14:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5516[14:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5511[14:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5501[14:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5486[14:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5446[14:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5461[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1e)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub12_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h3: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6f)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp870[14:0] );

									end
									else
									if((r_sys_run_step==9'h6e)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp864[14:0] );

									end
									else
									if((r_sys_run_step==9'h7d)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp954[14:0] );

									end
									else
									if((r_sys_run_step==9'h72)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp888[14:0] );

									end
									else
									if((r_sys_run_step==9'h73)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp894[14:0] );

									end
									else
									if((r_sys_run_step==9'h67)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp810[14:0] );

									end
									else
									if((r_sys_run_step==9'h6c)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp852[14:0] );

									end
									else
									if((r_sys_run_step==9'h75)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp906[14:0] );

									end
									else
									if((r_sys_run_step==9'h82)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp984[14:0] );

									end
									else
									if((r_sys_run_step==9'h7a)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp936[14:0] );

									end
									else
									if((r_sys_run_step==9'h71)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp882[14:0] );

									end
									else
									if((r_sys_run_step==9'h7b)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp942[14:0] );

									end
									else
									if((r_sys_run_step==9'h80)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp972[14:0] );

									end
									else
									if((r_sys_run_step==9'h86)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp1008[14:0] );

									end
									else
									if((r_sys_run_step==9'h70)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp876[14:0] );

									end
									else
									if((r_sys_run_step==9'h6a)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp840[14:0] );

									end
									else
									if((r_sys_run_step==9'h88)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp1020[14:0] );

									end
									else
									if((r_sys_run_step==9'h69)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp834[14:0] );

									end
									else
									if((r_sys_run_step==9'h6b)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp846[14:0] );

									end
									else
									if((r_sys_run_step==9'h87)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp1014[14:0] );

									end
									else
									if((r_sys_run_step==9'h83)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp990[14:0] );

									end
									else
									if((r_sys_run_step==9'h77)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp918[14:0] );

									end
									else
									if((r_sys_run_step==9'h79)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp930[14:0] );

									end
									else
									if((r_sys_run_step==9'h85)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp1002[14:0] );

									end
									else
									if((r_sys_run_step==9'h78)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp924[14:0] );

									end
									else
									if((r_sys_run_step==9'h7e)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp960[14:0] );

									end
									else
									if((r_sys_run_step==9'h81)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp978[14:0] );

									end
									else
									if((r_sys_run_step==9'h6d)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp858[14:0] );

									end
									else
									if((r_sys_run_step==9'h76)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp912[14:0] );

									end
									else
									if((r_sys_run_step==9'h68)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp816[14:0] );

									end
									else
									if((r_sys_run_step==9'h74)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp900[14:0] );

									end
									else
									if((r_sys_run_step==9'h84)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp996[14:0] );

									end
									else
									if((r_sys_run_step==9'h7f)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp966[14:0] );

									end
									else
									if((r_sys_run_step==9'h7c)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp948[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h67<=r_sys_run_step && r_sys_run_step<=9'h88)) begin
										r_sub03_u_datain <= w_sys_tmp218;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h67<=r_sys_run_step && r_sys_run_step<=9'h88)) begin
										r_sub03_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub03_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4014[14:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4084[14:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4039[14:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4004[14:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4059[14:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4119[14:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4124[14:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp3994[14:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp3979[14:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp3984[14:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp3974[14:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4074[14:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4089[14:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4114[14:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4044[14:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4054[14:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4109[14:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4019[14:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4064[14:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp3999[14:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp3989[14:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4094[14:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4034[14:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4079[14:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4029[14:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4099[14:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4129[14:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4049[14:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4009[14:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4104[14:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4024[14:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4069[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1f)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub03_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h2: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4f)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp678[14:0] );

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp672[14:0] );

									end
									else
									if((r_sys_run_step==9'h65)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp810[14:0] );

									end
									else
									if((r_sys_run_step==9'h63)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp798[14:0] );

									end
									else
									if((r_sys_run_step==9'h5f)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp774[14:0] );

									end
									else
									if((r_sys_run_step==9'h5a)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp744[14:0] );

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp708[14:0] );

									end
									else
									if((r_sys_run_step==9'h5b)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp750[14:0] );

									end
									else
									if((r_sys_run_step==9'h48)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp636[14:0] );

									end
									else
									if((r_sys_run_step==9'h57)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp726[14:0] );

									end
									else
									if((r_sys_run_step==9'h5c)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp756[14:0] );

									end
									else
									if((r_sys_run_step==9'h64)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp804[14:0] );

									end
									else
									if((r_sys_run_step==9'h46)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp612[14:0] );

									end
									else
									if((r_sys_run_step==9'h59)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp738[14:0] );

									end
									else
									if((r_sys_run_step==9'h62)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp792[14:0] );

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp654[14:0] );

									end
									else
									if((r_sys_run_step==9'h5e)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp768[14:0] );

									end
									else
									if((r_sys_run_step==9'h55)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp714[14:0] );

									end
									else
									if((r_sys_run_step==9'h4a)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp648[14:0] );

									end
									else
									if((r_sys_run_step==9'h53)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp702[14:0] );

									end
									else
									if((r_sys_run_step==9'h61)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp786[14:0] );

									end
									else
									if((r_sys_run_step==9'h4d)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp666[14:0] );

									end
									else
									if((r_sys_run_step==9'h56)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp720[14:0] );

									end
									else
									if((r_sys_run_step==9'h51)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp690[14:0] );

									end
									else
									if((r_sys_run_step==9'h45)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp606[14:0] );

									end
									else
									if((r_sys_run_step==9'h66)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp816[14:0] );

									end
									else
									if((r_sys_run_step==9'h60)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp780[14:0] );

									end
									else
									if((r_sys_run_step==9'h50)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp684[14:0] );

									end
									else
									if((r_sys_run_step==9'h49)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp642[14:0] );

									end
									else
									if((r_sys_run_step==9'h58)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp732[14:0] );

									end
									else
									if((r_sys_run_step==9'h5d)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp762[14:0] );

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp630[14:0] );

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp660[14:0] );

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp696[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h45<=r_sys_run_step && r_sys_run_step<=9'h66)) begin
										r_sub02_u_datain <= w_sys_tmp218;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h45<=r_sys_run_step && r_sys_run_step<=9'h66)) begin
										r_sub02_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub02_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3934[14:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3889[14:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3844[14:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3924[14:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3834[14:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3874[14:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3909[14:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3944[14:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3854[14:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3914[14:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3959[14:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3839[14:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3964[14:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3894[14:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3949[14:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3859[14:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3829[14:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3869[14:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3864[14:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3969[14:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3879[14:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3819[14:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3814[14:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3884[14:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3904[14:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3939[14:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3929[14:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3899[14:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3849[14:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3954[14:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3824[14:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3919[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1f)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub02_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h9: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub11_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub11_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hff)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2550[14:0] );

									end
									else
									if((r_sys_run_step==9'h100)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2556[14:0] );

									end
									else
									if((r_sys_run_step==9'hf3)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2478[14:0] );

									end
									else
									if((r_sys_run_step==9'hef)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2442[14:0] );

									end
									else
									if((r_sys_run_step==9'hf6)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2496[14:0] );

									end
									else
									if((r_sys_run_step==9'h108)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2604[14:0] );

									end
									else
									if((r_sys_run_step==9'h103)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2574[14:0] );

									end
									else
									if((r_sys_run_step==9'hf1)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2466[14:0] );

									end
									else
									if((r_sys_run_step==9'h10a)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2616[14:0] );

									end
									else
									if((r_sys_run_step==9'h102)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2568[14:0] );

									end
									else
									if((r_sys_run_step==9'hf0)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2460[14:0] );

									end
									else
									if((r_sys_run_step==9'h109)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2610[14:0] );

									end
									else
									if((r_sys_run_step==9'h106)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2592[14:0] );

									end
									else
									if((r_sys_run_step==9'h10e)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2640[14:0] );

									end
									else
									if((r_sys_run_step==9'h10b)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2622[14:0] );

									end
									else
									if((r_sys_run_step==9'h10f)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2646[14:0] );

									end
									else
									if((r_sys_run_step==9'hf5)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2490[14:0] );

									end
									else
									if((r_sys_run_step==9'h10c)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2628[14:0] );

									end
									else
									if((r_sys_run_step==9'hfb)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2526[14:0] );

									end
									else
									if((r_sys_run_step==9'hee)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2436[14:0] );

									end
									else
									if((r_sys_run_step==9'hf8)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2508[14:0] );

									end
									else
									if((r_sys_run_step==9'hf2)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2472[14:0] );

									end
									else
									if((r_sys_run_step==9'hfc)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2532[14:0] );

									end
									else
									if((r_sys_run_step==9'hfd)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2538[14:0] );

									end
									else
									if((r_sys_run_step==9'h107)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2598[14:0] );

									end
									else
									if((r_sys_run_step==9'hf9)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2514[14:0] );

									end
									else
									if((r_sys_run_step==9'hfa)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2520[14:0] );

									end
									else
									if((r_sys_run_step==9'h101)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2562[14:0] );

									end
									else
									if((r_sys_run_step==9'hf7)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2502[14:0] );

									end
									else
									if((r_sys_run_step==9'h105)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2586[14:0] );

									end
									else
									if((r_sys_run_step==9'hf4)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2484[14:0] );

									end
									else
									if((r_sys_run_step==9'h10d)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2634[14:0] );

									end
									else
									if((r_sys_run_step==9'hfe)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2544[14:0] );

									end
									else
									if((r_sys_run_step==9'h104)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp2580[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'hee<=r_sys_run_step && r_sys_run_step<=9'h10f)) begin
										r_sub11_u_datain <= w_sys_tmp1034;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'hee<=r_sys_run_step && r_sys_run_step<=9'h10f)) begin
										r_sub11_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub11_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1a)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5411[14:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5346[14:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5391[14:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5386[14:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5281[14:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5326[14:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5406[14:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5401[14:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5311[14:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5296[14:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5356[14:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5331[14:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5396[14:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5421[14:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5361[14:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5366[14:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5431[14:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5436[14:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5336[14:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5371[14:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5306[14:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5381[14:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5291[14:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5321[14:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5351[14:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5416[14:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5426[14:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5341[14:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5376[14:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5286[14:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5316[14:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5301[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1f)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub11_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'hb: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub14_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub14_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15f)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3126[14:0] );

									end
									else
									if((r_sys_run_step==9'h174)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3252[14:0] );

									end
									else
									if((r_sys_run_step==9'h171)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3234[14:0] );

									end
									else
									if((r_sys_run_step==9'h15e)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3120[14:0] );

									end
									else
									if((r_sys_run_step==9'h155)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3066[14:0] );

									end
									else
									if((r_sys_run_step==9'h154)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3048[14:0] );

									end
									else
									if((r_sys_run_step==9'h15b)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3102[14:0] );

									end
									else
									if((r_sys_run_step==9'h156)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3072[14:0] );

									end
									else
									if((r_sys_run_step==9'h16f)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3222[14:0] );

									end
									else
									if((r_sys_run_step==9'h159)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3090[14:0] );

									end
									else
									if((r_sys_run_step==9'h16a)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3192[14:0] );

									end
									else
									if((r_sys_run_step==9'h170)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3228[14:0] );

									end
									else
									if((r_sys_run_step==9'h15c)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3108[14:0] );

									end
									else
									if((r_sys_run_step==9'h15d)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3114[14:0] );

									end
									else
									if((r_sys_run_step==9'h16e)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3216[14:0] );

									end
									else
									if((r_sys_run_step==9'h163)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3150[14:0] );

									end
									else
									if((r_sys_run_step==9'h167)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3174[14:0] );

									end
									else
									if((r_sys_run_step==9'h161)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3138[14:0] );

									end
									else
									if((r_sys_run_step==9'h160)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3132[14:0] );

									end
									else
									if((r_sys_run_step==9'h157)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3078[14:0] );

									end
									else
									if((r_sys_run_step==9'h166)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3168[14:0] );

									end
									else
									if((r_sys_run_step==9'h165)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3162[14:0] );

									end
									else
									if((r_sys_run_step==9'h16d)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3210[14:0] );

									end
									else
									if((r_sys_run_step==9'h172)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3240[14:0] );

									end
									else
									if((r_sys_run_step==9'h158)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3084[14:0] );

									end
									else
									if((r_sys_run_step==9'h169)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3186[14:0] );

									end
									else
									if((r_sys_run_step==9'h15a)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3096[14:0] );

									end
									else
									if((r_sys_run_step==9'h16c)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3204[14:0] );

									end
									else
									if((r_sys_run_step==9'h164)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3156[14:0] );

									end
									else
									if((r_sys_run_step==9'h162)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3144[14:0] );

									end
									else
									if((r_sys_run_step==9'h16b)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3198[14:0] );

									end
									else
									if((r_sys_run_step==9'h173)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3246[14:0] );

									end
									else
									if((r_sys_run_step==9'h168)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3180[14:0] );

									end
									else
									if((r_sys_run_step==9'h153)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp3042[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h153<=r_sys_run_step && r_sys_run_step<=9'h174)) begin
										r_sub14_u_datain <= w_sys_tmp1034;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h153<=r_sys_run_step && r_sys_run_step<=9'h174)) begin
										r_sub14_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub14_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5766[14:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5891[14:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5831[14:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5896[14:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5806[14:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5866[14:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5906[14:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5761[14:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5776[14:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5846[14:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5816[14:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5841[14:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5901[14:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5786[14:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5821[14:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5911[14:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5861[14:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5836[14:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5876[14:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5826[14:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5871[14:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5856[14:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5881[14:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5796[14:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5886[14:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5771[14:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5791[14:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5811[14:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5801[14:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5781[14:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5756[14:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5851[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1f)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub14_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h32)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp504[14:0] );

									end
									else
									if((r_sys_run_step==9'h35)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp522[14:0] );

									end
									else
									if((r_sys_run_step==9'h42)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp600[14:0] );

									end
									else
									if((r_sys_run_step==9'h2c)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp468[14:0] );

									end
									else
									if((r_sys_run_step==9'h23)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp402[14:0] );

									end
									else
									if((r_sys_run_step==9'h30)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp492[14:0] );

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp426[14:0] );

									end
									else
									if((r_sys_run_step==9'h3f)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp582[14:0] );

									end
									else
									if((r_sys_run_step==9'h40)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp588[14:0] );

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp570[14:0] );

									end
									else
									if((r_sys_run_step==9'h29)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp450[14:0] );

									end
									else
									if((r_sys_run_step==9'h26)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp432[14:0] );

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp486[14:0] );

									end
									else
									if((r_sys_run_step==9'h33)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp510[14:0] );

									end
									else
									if((r_sys_run_step==9'h44)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp612[14:0] );

									end
									else
									if((r_sys_run_step==9'h2a)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp456[14:0] );

									end
									else
									if((r_sys_run_step==9'h37)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp534[14:0] );

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp564[14:0] );

									end
									else
									if((r_sys_run_step==9'h34)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp516[14:0] );

									end
									else
									if((r_sys_run_step==9'h3a)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp552[14:0] );

									end
									else
									if((r_sys_run_step==9'h2e)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp480[14:0] );

									end
									else
									if((r_sys_run_step==9'h3e)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp576[14:0] );

									end
									else
									if((r_sys_run_step==9'h43)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp606[14:0] );

									end
									else
									if((r_sys_run_step==9'h2b)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp462[14:0] );

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp408[14:0] );

									end
									else
									if((r_sys_run_step==9'h28)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp444[14:0] );

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp546[14:0] );

									end
									else
									if((r_sys_run_step==9'h27)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp438[14:0] );

									end
									else
									if((r_sys_run_step==9'h38)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp540[14:0] );

									end
									else
									if((r_sys_run_step==9'h2d)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp474[14:0] );

									end
									else
									if((r_sys_run_step==9'h36)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp528[14:0] );

									end
									else
									if((r_sys_run_step==9'h41)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp594[14:0] );

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp558[14:0] );

									end
									else
									if((r_sys_run_step==9'h31)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp498[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h23<=r_sys_run_step && r_sys_run_step<=9'h44)) begin
										r_sub01_u_datain <= w_sys_tmp218;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h23<=r_sys_run_step && r_sys_run_step<=9'h44)) begin
										r_sub01_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub01_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1e)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3804[14:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3664[14:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3669[14:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3704[14:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3734[14:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3749[14:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3794[14:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3799[14:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3689[14:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3659[14:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3714[14:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3784[14:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3699[14:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3719[14:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3789[14:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3709[14:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3679[14:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3729[14:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3759[14:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3809[14:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3739[14:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3769[14:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3779[14:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3774[14:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3674[14:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3654[14:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3684[14:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3764[14:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3754[14:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3724[14:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3694[14:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3744[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1f)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'ha: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub13_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub13_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14a)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp3000[14:0] );

									end
									else
									if((r_sys_run_step==9'h148)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2988[14:0] );

									end
									else
									if((r_sys_run_step==9'h152)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp3048[14:0] );

									end
									else
									if((r_sys_run_step==9'h138)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2892[14:0] );

									end
									else
									if((r_sys_run_step==9'h13d)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2922[14:0] );

									end
									else
									if((r_sys_run_step==9'h132)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2844[14:0] );

									end
									else
									if((r_sys_run_step==9'h13f)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2934[14:0] );

									end
									else
									if((r_sys_run_step==9'h149)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2994[14:0] );

									end
									else
									if((r_sys_run_step==9'h135)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2874[14:0] );

									end
									else
									if((r_sys_run_step==9'h140)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2940[14:0] );

									end
									else
									if((r_sys_run_step==9'h13c)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2916[14:0] );

									end
									else
									if((r_sys_run_step==9'h150)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp3036[14:0] );

									end
									else
									if((r_sys_run_step==9'h133)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2862[14:0] );

									end
									else
									if((r_sys_run_step==9'h147)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2982[14:0] );

									end
									else
									if((r_sys_run_step==9'h136)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2880[14:0] );

									end
									else
									if((r_sys_run_step==9'h141)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2946[14:0] );

									end
									else
									if((r_sys_run_step==9'h144)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2964[14:0] );

									end
									else
									if((r_sys_run_step==9'h14d)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp3018[14:0] );

									end
									else
									if((r_sys_run_step==9'h139)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2898[14:0] );

									end
									else
									if((r_sys_run_step==9'h134)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2868[14:0] );

									end
									else
									if((r_sys_run_step==9'h142)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2952[14:0] );

									end
									else
									if((r_sys_run_step==9'h14b)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp3006[14:0] );

									end
									else
									if((r_sys_run_step==9'h146)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2976[14:0] );

									end
									else
									if((r_sys_run_step==9'h145)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2970[14:0] );

									end
									else
									if((r_sys_run_step==9'h14f)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp3030[14:0] );

									end
									else
									if((r_sys_run_step==9'h143)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2958[14:0] );

									end
									else
									if((r_sys_run_step==9'h13b)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2910[14:0] );

									end
									else
									if((r_sys_run_step==9'h13e)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2928[14:0] );

									end
									else
									if((r_sys_run_step==9'h14e)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp3024[14:0] );

									end
									else
									if((r_sys_run_step==9'h13a)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2904[14:0] );

									end
									else
									if((r_sys_run_step==9'h137)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2886[14:0] );

									end
									else
									if((r_sys_run_step==9'h131)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp2838[14:0] );

									end
									else
									if((r_sys_run_step==9'h151)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp3042[14:0] );

									end
									else
									if((r_sys_run_step==9'h14c)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp3012[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h131<=r_sys_run_step && r_sys_run_step<=9'h152)) begin
										r_sub13_u_datain <= w_sys_tmp1034;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h131<=r_sys_run_step && r_sys_run_step<=9'h152)) begin
										r_sub13_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub13_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5611[14:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5656[14:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5701[14:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5596[14:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5741[14:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5651[14:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5746[14:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5721[14:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5616[14:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5726[14:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5621[14:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5706[14:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5601[14:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5606[14:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5631[14:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5691[14:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5731[14:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5626[14:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5736[14:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5666[14:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5636[14:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5711[14:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5661[14:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5686[14:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5696[14:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5671[14:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5751[14:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5646[14:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5676[14:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5681[14:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5716[14:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5641[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1f)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub13_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp366[14:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp390[14:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp258[14:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp252[14:0] );

									end
									else
									if((r_sys_run_step==9'h21)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp402[14:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp216[14:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp360[14:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp294[14:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp306[14:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp372[14:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp264[14:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp228[14:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp378[14:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp312[14:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp330[14:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp282[14:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp384[14:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp276[14:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp336[14:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp318[14:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp354[14:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp348[14:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp246[14:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp300[14:0] );

									end
									else
									if((r_sys_run_step==9'h20)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp396[14:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp240[14:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp342[14:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp222[14:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp234[14:0] );

									end
									else
									if((r_sys_run_step==9'h22)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp408[14:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp324[14:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp270[14:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp288[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h22)) begin
										r_sub00_u_datain <= w_sys_tmp218;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h22)) begin
										r_sub00_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub00_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3468[14:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3510[14:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3594[14:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3480[14:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3612[14:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3618[14:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3558[14:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3498[14:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3528[14:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3504[14:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3534[14:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3576[14:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3516[14:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3492[14:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3636[14:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3600[14:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3630[14:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3642[14:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3588[14:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3546[14:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3474[14:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3648[14:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3564[14:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3570[14:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3624[14:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3486[14:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3606[14:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3522[14:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3582[14:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3552[14:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3540[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1e)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h6: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub07_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub07_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h82)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1800[14:0] );

									end
									else
									if((r_sys_run_step==9'h6d)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1674[14:0] );

									end
									else
									if((r_sys_run_step==9'h73)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1710[14:0] );

									end
									else
									if((r_sys_run_step==9'h75)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1722[14:0] );

									end
									else
									if((r_sys_run_step==9'h83)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1806[14:0] );

									end
									else
									if((r_sys_run_step==9'h78)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1740[14:0] );

									end
									else
									if((r_sys_run_step==9'h67)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1626[14:0] );

									end
									else
									if((r_sys_run_step==9'h68)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1632[14:0] );

									end
									else
									if((r_sys_run_step==9'h7e)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1776[14:0] );

									end
									else
									if((r_sys_run_step==9'h6f)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1686[14:0] );

									end
									else
									if((r_sys_run_step==9'h71)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1698[14:0] );

									end
									else
									if((r_sys_run_step==9'h7c)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1764[14:0] );

									end
									else
									if((r_sys_run_step==9'h7a)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1752[14:0] );

									end
									else
									if((r_sys_run_step==9'h7b)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1758[14:0] );

									end
									else
									if((r_sys_run_step==9'h88)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1836[14:0] );

									end
									else
									if((r_sys_run_step==9'h86)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1824[14:0] );

									end
									else
									if((r_sys_run_step==9'h7f)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1782[14:0] );

									end
									else
									if((r_sys_run_step==9'h84)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1812[14:0] );

									end
									else
									if((r_sys_run_step==9'h70)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1692[14:0] );

									end
									else
									if((r_sys_run_step==9'h79)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1746[14:0] );

									end
									else
									if((r_sys_run_step==9'h81)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1794[14:0] );

									end
									else
									if((r_sys_run_step==9'h77)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1734[14:0] );

									end
									else
									if((r_sys_run_step==9'h72)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1704[14:0] );

									end
									else
									if((r_sys_run_step==9'h85)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1818[14:0] );

									end
									else
									if((r_sys_run_step==9'h6c)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1668[14:0] );

									end
									else
									if((r_sys_run_step==9'h87)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1830[14:0] );

									end
									else
									if((r_sys_run_step==9'h6b)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1662[14:0] );

									end
									else
									if((r_sys_run_step==9'h6a)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1656[14:0] );

									end
									else
									if((r_sys_run_step==9'h7d)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1770[14:0] );

									end
									else
									if((r_sys_run_step==9'h80)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1788[14:0] );

									end
									else
									if((r_sys_run_step==9'h6e)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1680[14:0] );

									end
									else
									if((r_sys_run_step==9'h69)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1650[14:0] );

									end
									else
									if((r_sys_run_step==9'h76)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1728[14:0] );

									end
									else
									if((r_sys_run_step==9'h74)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1716[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h67<=r_sys_run_step && r_sys_run_step<=9'h88)) begin
										r_sub07_u_datain <= w_sys_tmp1034;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h67<=r_sys_run_step && r_sys_run_step<=9'h88)) begin
										r_sub07_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub07_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4781[14:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4666[14:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4746[14:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4776[14:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4741[14:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4716[14:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4721[14:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4661[14:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4651[14:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4676[14:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4711[14:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4801[14:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4691[14:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4756[14:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4686[14:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4766[14:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4786[14:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4646[14:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4761[14:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4771[14:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4751[14:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4796[14:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4696[14:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4726[14:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4671[14:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4706[14:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4736[14:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4681[14:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4701[14:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4791[14:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4656[14:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4731[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1f)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub07_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h5: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub06_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub06_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5e)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1584[14:0] );

									end
									else
									if((r_sys_run_step==9'h4f)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1494[14:0] );

									end
									else
									if((r_sys_run_step==9'h65)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1626[14:0] );

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1470[14:0] );

									end
									else
									if((r_sys_run_step==9'h66)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1632[14:0] );

									end
									else
									if((r_sys_run_step==9'h61)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1602[14:0] );

									end
									else
									if((r_sys_run_step==9'h55)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1530[14:0] );

									end
									else
									if((r_sys_run_step==9'h58)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1548[14:0] );

									end
									else
									if((r_sys_run_step==9'h63)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1614[14:0] );

									end
									else
									if((r_sys_run_step==9'h56)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1536[14:0] );

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1524[14:0] );

									end
									else
									if((r_sys_run_step==9'h64)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1620[14:0] );

									end
									else
									if((r_sys_run_step==9'h57)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1542[14:0] );

									end
									else
									if((r_sys_run_step==9'h51)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1506[14:0] );

									end
									else
									if((r_sys_run_step==9'h5f)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1590[14:0] );

									end
									else
									if((r_sys_run_step==9'h53)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1518[14:0] );

									end
									else
									if((r_sys_run_step==9'h49)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1458[14:0] );

									end
									else
									if((r_sys_run_step==9'h46)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1428[14:0] );

									end
									else
									if((r_sys_run_step==9'h62)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1608[14:0] );

									end
									else
									if((r_sys_run_step==9'h4a)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1464[14:0] );

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1446[14:0] );

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1488[14:0] );

									end
									else
									if((r_sys_run_step==9'h4d)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1482[14:0] );

									end
									else
									if((r_sys_run_step==9'h5c)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1572[14:0] );

									end
									else
									if((r_sys_run_step==9'h50)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1500[14:0] );

									end
									else
									if((r_sys_run_step==9'h59)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1554[14:0] );

									end
									else
									if((r_sys_run_step==9'h5d)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1578[14:0] );

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1476[14:0] );

									end
									else
									if((r_sys_run_step==9'h60)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1596[14:0] );

									end
									else
									if((r_sys_run_step==9'h45)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1422[14:0] );

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1512[14:0] );

									end
									else
									if((r_sys_run_step==9'h48)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1452[14:0] );

									end
									else
									if((r_sys_run_step==9'h5a)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1560[14:0] );

									end
									else
									if((r_sys_run_step==9'h5b)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1566[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h45<=r_sys_run_step && r_sys_run_step<=9'h66)) begin
										r_sub06_u_datain <= w_sys_tmp1034;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h45<=r_sys_run_step && r_sys_run_step<=9'h66)) begin
										r_sub06_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub06_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4536[14:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4626[14:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4491[14:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4566[14:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4596[14:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4496[14:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4561[14:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4551[14:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4631[14:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4576[14:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4526[14:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4506[14:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4636[14:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4606[14:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4486[14:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4546[14:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4601[14:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4581[14:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4641[14:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4621[14:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4611[14:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4556[14:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4521[14:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4531[14:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4511[14:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4586[14:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4501[14:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4571[14:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4616[14:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4516[14:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4541[14:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4591[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1f)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub06_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'hc: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub15_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub15_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h176)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3252[14:0] );

									end
									else
									if((r_sys_run_step==9'h188)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3372[14:0] );

									end
									else
									if((r_sys_run_step==9'h193)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3438[14:0] );

									end
									else
									if((r_sys_run_step==9'h192)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3432[14:0] );

									end
									else
									if((r_sys_run_step==9'h17c)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3300[14:0] );

									end
									else
									if((r_sys_run_step==9'h179)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3282[14:0] );

									end
									else
									if((r_sys_run_step==9'h186)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3360[14:0] );

									end
									else
									if((r_sys_run_step==9'h177)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3270[14:0] );

									end
									else
									if((r_sys_run_step==9'h194)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3444[14:0] );

									end
									else
									if((r_sys_run_step==9'h182)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3336[14:0] );

									end
									else
									if((r_sys_run_step==9'h18b)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3390[14:0] );

									end
									else
									if((r_sys_run_step==9'h18e)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3408[14:0] );

									end
									else
									if((r_sys_run_step==9'h18d)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3402[14:0] );

									end
									else
									if((r_sys_run_step==9'h18a)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3384[14:0] );

									end
									else
									if((r_sys_run_step==9'h18f)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3414[14:0] );

									end
									else
									if((r_sys_run_step==9'h195)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3450[14:0] );

									end
									else
									if((r_sys_run_step==9'h183)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3342[14:0] );

									end
									else
									if((r_sys_run_step==9'h187)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3366[14:0] );

									end
									else
									if((r_sys_run_step==9'h178)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3276[14:0] );

									end
									else
									if((r_sys_run_step==9'h17a)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3288[14:0] );

									end
									else
									if((r_sys_run_step==9'h196)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3456[14:0] );

									end
									else
									if((r_sys_run_step==9'h17d)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3306[14:0] );

									end
									else
									if((r_sys_run_step==9'h17f)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3318[14:0] );

									end
									else
									if((r_sys_run_step==9'h181)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3330[14:0] );

									end
									else
									if((r_sys_run_step==9'h185)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3354[14:0] );

									end
									else
									if((r_sys_run_step==9'h180)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3324[14:0] );

									end
									else
									if((r_sys_run_step==9'h17b)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3294[14:0] );

									end
									else
									if((r_sys_run_step==9'h17e)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3312[14:0] );

									end
									else
									if((r_sys_run_step==9'h18c)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3396[14:0] );

									end
									else
									if((r_sys_run_step==9'h190)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3420[14:0] );

									end
									else
									if((r_sys_run_step==9'h175)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3246[14:0] );

									end
									else
									if((r_sys_run_step==9'h184)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3348[14:0] );

									end
									else
									if((r_sys_run_step==9'h191)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3426[14:0] );

									end
									else
									if((r_sys_run_step==9'h189)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp3378[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h175<=r_sys_run_step && r_sys_run_step<=9'h196)) begin
										r_sub15_u_datain <= w_sys_tmp1034;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h175<=r_sys_run_step && r_sys_run_step<=9'h196)) begin
										r_sub15_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub15_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp5981[14:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp6031[14:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp5931[14:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp6001[14:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp5966[14:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp5971[14:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp5951[14:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp5921[14:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp6056[14:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp6066[14:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp6041[14:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp5926[14:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp6061[14:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp5956[14:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp6006[14:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp6011[14:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp6036[14:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp6021[14:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp6046[14:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp5986[14:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp6071[14:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp5946[14:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp5996[14:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp5916[14:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp5976[14:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp5941[14:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp5961[14:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp5936[14:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp5991[14:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp6026[14:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp6016[14:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp6051[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1f)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub15_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h4: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub05_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub05_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2a)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1272[14:0] );

									end
									else
									if((r_sys_run_step==9'h37)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1350[14:0] );

									end
									else
									if((r_sys_run_step==9'h28)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1260[14:0] );

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1302[14:0] );

									end
									else
									if((r_sys_run_step==9'h3a)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1368[14:0] );

									end
									else
									if((r_sys_run_step==9'h2c)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1284[14:0] );

									end
									else
									if((r_sys_run_step==9'h29)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1266[14:0] );

									end
									else
									if((r_sys_run_step==9'h35)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1338[14:0] );

									end
									else
									if((r_sys_run_step==9'h32)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1320[14:0] );

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1224[14:0] );

									end
									else
									if((r_sys_run_step==9'h2b)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1278[14:0] );

									end
									else
									if((r_sys_run_step==9'h34)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1332[14:0] );

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1242[14:0] );

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1386[14:0] );

									end
									else
									if((r_sys_run_step==9'h3e)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1392[14:0] );

									end
									else
									if((r_sys_run_step==9'h2d)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1290[14:0] );

									end
									else
									if((r_sys_run_step==9'h26)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1248[14:0] );

									end
									else
									if((r_sys_run_step==9'h27)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1254[14:0] );

									end
									else
									if((r_sys_run_step==9'h31)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1314[14:0] );

									end
									else
									if((r_sys_run_step==9'h42)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1416[14:0] );

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1374[14:0] );

									end
									else
									if((r_sys_run_step==9'h33)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1326[14:0] );

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1362[14:0] );

									end
									else
									if((r_sys_run_step==9'h23)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1218[14:0] );

									end
									else
									if((r_sys_run_step==9'h44)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1428[14:0] );

									end
									else
									if((r_sys_run_step==9'h36)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1344[14:0] );

									end
									else
									if((r_sys_run_step==9'h30)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1308[14:0] );

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1380[14:0] );

									end
									else
									if((r_sys_run_step==9'h41)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1410[14:0] );

									end
									else
									if((r_sys_run_step==9'h40)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1404[14:0] );

									end
									else
									if((r_sys_run_step==9'h43)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1422[14:0] );

									end
									else
									if((r_sys_run_step==9'h3f)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1398[14:0] );

									end
									else
									if((r_sys_run_step==9'h38)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1356[14:0] );

									end
									else
									if((r_sys_run_step==9'h2e)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1296[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h23<=r_sys_run_step && r_sys_run_step<=9'h44)) begin
										r_sub05_u_datain <= w_sys_tmp1034;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h23<=r_sys_run_step && r_sys_run_step<=9'h44)) begin
										r_sub05_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub05_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4446[14:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4441[14:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4351[14:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4336[14:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4406[14:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4416[14:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4466[14:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4386[14:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4456[14:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4326[14:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4476[14:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4391[14:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4451[14:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4366[14:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4346[14:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4381[14:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4426[14:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4396[14:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4376[14:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4401[14:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4421[14:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4431[14:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4471[14:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4356[14:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4341[14:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4411[14:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4331[14:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4481[14:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4461[14:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4436[14:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4371[14:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4361[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1f)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub05_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'he: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub04_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub04_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1182[14:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1170[14:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1068[14:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1164[14:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1206[14:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1050[14:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1110[14:0] );

									end
									else
									if((r_sys_run_step==9'h22)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1224[14:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1140[14:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1032[14:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1062[14:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1038[14:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1128[14:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1074[14:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1188[14:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1086[14:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1104[14:0] );

									end
									else
									if((r_sys_run_step==9'h20)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1212[14:0] );

									end
									else
									if((r_sys_run_step==9'h21)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1218[14:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1134[14:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1158[14:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1098[14:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1122[14:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1080[14:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1176[14:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1200[14:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1044[14:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1092[14:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1056[14:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1146[14:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1116[14:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1194[14:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1152[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h22)) begin
										r_sub04_u_datain <= w_sys_tmp1034;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h22)) begin
										r_sub04_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub04_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1a)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4296[14:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4200[14:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4284[14:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4236[14:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4314[14:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4302[14:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4254[14:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4278[14:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4308[14:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4230[14:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4290[14:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4224[14:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4140[14:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4206[14:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4320[14:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4248[14:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4260[14:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4218[14:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4146[14:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4176[14:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4266[14:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4242[14:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4272[14:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4158[14:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4170[14:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4182[14:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4212[14:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4194[14:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4188[14:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4164[14:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4152[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1e)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub04_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h8: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub10_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub10_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hed)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2442[14:0] );

									end
									else
									if((r_sys_run_step==9'he4)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2388[14:0] );

									end
									else
									if((r_sys_run_step==9'he7)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2406[14:0] );

									end
									else
									if((r_sys_run_step==9'heb)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2430[14:0] );

									end
									else
									if((r_sys_run_step==9'hda)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2328[14:0] );

									end
									else
									if((r_sys_run_step==9'hcf)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2262[14:0] );

									end
									else
									if((r_sys_run_step==9'hd5)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2298[14:0] );

									end
									else
									if((r_sys_run_step==9'he8)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2412[14:0] );

									end
									else
									if((r_sys_run_step==9'hd0)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2268[14:0] );

									end
									else
									if((r_sys_run_step==9'hd8)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2316[14:0] );

									end
									else
									if((r_sys_run_step==9'hdb)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2334[14:0] );

									end
									else
									if((r_sys_run_step==9'he9)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2418[14:0] );

									end
									else
									if((r_sys_run_step==9'hdc)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2340[14:0] );

									end
									else
									if((r_sys_run_step==9'hd9)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2322[14:0] );

									end
									else
									if((r_sys_run_step==9'he0)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2364[14:0] );

									end
									else
									if((r_sys_run_step==9'hdf)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2358[14:0] );

									end
									else
									if((r_sys_run_step==9'hd2)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2280[14:0] );

									end
									else
									if((r_sys_run_step==9'he5)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2394[14:0] );

									end
									else
									if((r_sys_run_step==9'hd6)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2304[14:0] );

									end
									else
									if((r_sys_run_step==9'hcd)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2238[14:0] );

									end
									else
									if((r_sys_run_step==9'hce)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2256[14:0] );

									end
									else
									if((r_sys_run_step==9'hde)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2352[14:0] );

									end
									else
									if((r_sys_run_step==9'hd1)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2274[14:0] );

									end
									else
									if((r_sys_run_step==9'he6)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2400[14:0] );

									end
									else
									if((r_sys_run_step==9'hea)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2424[14:0] );

									end
									else
									if((r_sys_run_step==9'hd3)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2286[14:0] );

									end
									else
									if((r_sys_run_step==9'hec)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2436[14:0] );

									end
									else
									if((r_sys_run_step==9'he2)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2376[14:0] );

									end
									else
									if((r_sys_run_step==9'hcc)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2232[14:0] );

									end
									else
									if((r_sys_run_step==9'hd7)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2310[14:0] );

									end
									else
									if((r_sys_run_step==9'hd4)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2292[14:0] );

									end
									else
									if((r_sys_run_step==9'he1)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2370[14:0] );

									end
									else
									if((r_sys_run_step==9'he3)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2382[14:0] );

									end
									else
									if((r_sys_run_step==9'hdd)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp2346[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'hcc<=r_sys_run_step && r_sys_run_step<=9'hed)) begin
										r_sub10_u_datain <= w_sys_tmp1034;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'hcc<=r_sys_run_step && r_sys_run_step<=9'hed)) begin
										r_sub10_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub10_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5121[14:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5156[14:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5271[14:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5126[14:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5141[14:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5256[14:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5146[14:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5171[14:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5196[14:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5131[14:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5181[14:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5161[14:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5136[14:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5191[14:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5276[14:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5206[14:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5231[14:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5226[14:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5236[14:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5211[14:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5201[14:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5216[14:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5241[14:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5176[14:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5186[14:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5251[14:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5246[14:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5151[14:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5266[14:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5261[14:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5221[14:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp5166[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1f)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub10_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h21)) begin
										r_sys_tmp0_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h21)) begin
										r_sys_tmp0_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h21)) begin
										r_sys_tmp1_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h21)) begin
										r_sys_tmp1_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h20)) begin
										r_sys_tmp2_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h21)) begin
										r_sys_tmp2_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h20)) begin
										r_sys_tmp3_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h21)) begin
										r_sys_tmp3_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h20)) begin
										r_sys_tmp4_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h21)) begin
										r_sys_tmp4_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1f)) begin
										r_sys_tmp5_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h21)) begin
										r_sys_tmp5_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1f)) begin
										r_sys_tmp6_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h21)) begin
										r_sys_tmp6_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1f)) begin
										r_sys_tmp7_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h21)) begin
										r_sys_tmp7_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1e)) begin
										r_sys_tmp8_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h20)) begin
										r_sys_tmp8_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1e)) begin
										r_sys_tmp9_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h20)) begin
										r_sys_tmp9_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1e)) begin
										r_sys_tmp10_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h20)) begin
										r_sys_tmp10_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1d)) begin
										r_sys_tmp11_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h20)) begin
										r_sys_tmp11_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1d)) begin
										r_sys_tmp12_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h20)) begin
										r_sys_tmp12_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1d)) begin
										r_sys_tmp13_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h20)) begin
										r_sys_tmp13_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1c)) begin
										r_sys_tmp14_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h20)) begin
										r_sys_tmp14_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1c)) begin
										r_sys_tmp15_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h20)) begin
										r_sys_tmp15_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1c)) begin
										r_sys_tmp16_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h20)) begin
										r_sys_tmp16_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sys_tmp17_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h20)) begin
										r_sys_tmp17_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sys_tmp18_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1f)) begin
										r_sys_tmp18_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sys_tmp19_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h20)) begin
										r_sys_tmp19_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1a)) begin
										r_sys_tmp20_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1f)) begin
										r_sys_tmp20_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1a)) begin
										r_sys_tmp21_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1f)) begin
										r_sys_tmp21_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1a)) begin
										r_sys_tmp22_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1f)) begin
										r_sys_tmp22_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h19)) begin
										r_sys_tmp23_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1f)) begin
										r_sys_tmp23_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h19)) begin
										r_sys_tmp24_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1f)) begin
										r_sys_tmp24_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h19)) begin
										r_sys_tmp25_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1f)) begin
										r_sys_tmp25_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_tmp26_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1f)) begin
										r_sys_tmp26_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_tmp27_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1f)) begin
										r_sys_tmp27_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_tmp28_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1f)) begin
										r_sys_tmp28_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h17)) begin
										r_sys_tmp29_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1f)) begin
										r_sys_tmp29_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h17)) begin
										r_sys_tmp30_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1e)) begin
										r_sys_tmp30_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h17)) begin
										r_sys_tmp31_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1e)) begin
										r_sys_tmp31_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h16)) begin
										r_sys_tmp32_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1e)) begin
										r_sys_tmp32_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h16)) begin
										r_sys_tmp33_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1e)) begin
										r_sys_tmp33_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h16)) begin
										r_sys_tmp34_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1e)) begin
										r_sys_tmp34_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp35_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1e)) begin
										r_sys_tmp35_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp36_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1e)) begin
										r_sys_tmp36_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp37_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1e)) begin
										r_sys_tmp37_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp38_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1e)) begin
										r_sys_tmp38_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp39_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1e)) begin
										r_sys_tmp39_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp40_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1d)) begin
										r_sys_tmp40_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp41_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1d)) begin
										r_sys_tmp41_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp42_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1e)) begin
										r_sys_tmp42_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp43_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1d)) begin
										r_sys_tmp43_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp44_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1d)) begin
										r_sys_tmp44_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp45_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1d)) begin
										r_sys_tmp45_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp46_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1d)) begin
										r_sys_tmp46_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp47_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1d)) begin
										r_sys_tmp47_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp48_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1d)) begin
										r_sys_tmp48_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp49_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1d)) begin
										r_sys_tmp49_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp50_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1d)) begin
										r_sys_tmp50_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp51_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1d)) begin
										r_sys_tmp51_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp52_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1c)) begin
										r_sys_tmp52_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp53_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1c)) begin
										r_sys_tmp53_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp54_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1c)) begin
										r_sys_tmp54_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp55_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1c)) begin
										r_sys_tmp55_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp56_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1c)) begin
										r_sys_tmp56_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp57_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1c)) begin
										r_sys_tmp57_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp58_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1c)) begin
										r_sys_tmp58_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp59_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1c)) begin
										r_sys_tmp59_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp60_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sys_tmp60_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp61_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1c)) begin
										r_sys_tmp61_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp62_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1c)) begin
										r_sys_tmp62_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp63_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1c)) begin
										r_sys_tmp63_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp64_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sys_tmp64_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp65_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sys_tmp65_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp66_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sys_tmp66_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp67_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sys_tmp67_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp68_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sys_tmp68_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp69_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sys_tmp69_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp70_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sys_tmp70_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp71_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sys_tmp71_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp72_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1a)) begin
										r_sys_tmp72_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp73_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1a)) begin
										r_sys_tmp73_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp74_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1a)) begin
										r_sys_tmp74_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp75_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1a)) begin
										r_sys_tmp75_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp76_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sys_tmp76_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp77_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sys_tmp77_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp78_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1a)) begin
										r_sys_tmp78_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp79_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1a)) begin
										r_sys_tmp79_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp80_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h19)) begin
										r_sys_tmp80_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp81_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1a)) begin
										r_sys_tmp81_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp82_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h19)) begin
										r_sys_tmp82_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp83_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h19)) begin
										r_sys_tmp83_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp84_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1a)) begin
										r_sys_tmp84_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp85_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1a)) begin
										r_sys_tmp85_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp86_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1a)) begin
										r_sys_tmp86_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp87_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1a)) begin
										r_sys_tmp87_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp88_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h19)) begin
										r_sys_tmp88_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp89_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h19)) begin
										r_sys_tmp89_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp90_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h19)) begin
										r_sys_tmp90_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp91_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h19)) begin
										r_sys_tmp91_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp92_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h19)) begin
										r_sys_tmp92_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp93_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h19)) begin
										r_sys_tmp93_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2) || (r_sys_run_step==9'h21)) begin
										r_sys_tmp94_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h19)) begin
										r_sys_tmp94_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h19)) begin
										r_sys_tmp95_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_tmp96_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_tmp97_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_tmp98_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_tmp99_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_tmp100_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_tmp101_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_tmp102_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_tmp103_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_tmp104_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_tmp105_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_tmp106_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h17)) begin
										r_sys_tmp107_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h17)) begin
										r_sys_tmp108_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h17)) begin
										r_sys_tmp109_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h17)) begin
										r_sys_tmp110_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h17)) begin
										r_sys_tmp111_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h17)) begin
										r_sys_tmp112_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h17)) begin
										r_sys_tmp113_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h17)) begin
										r_sys_tmp114_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h17)) begin
										r_sys_tmp115_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h17)) begin
										r_sys_tmp116_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h17)) begin
										r_sys_tmp117_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h16)) begin
										r_sys_tmp118_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h16)) begin
										r_sys_tmp119_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h16)) begin
										r_sys_tmp120_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h16)) begin
										r_sys_tmp121_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h16)) begin
										r_sys_tmp122_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h16)) begin
										r_sys_tmp123_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h16)) begin
										r_sys_tmp124_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h16)) begin
										r_sys_tmp125_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h16)) begin
										r_sys_tmp126_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h16)) begin
										r_sys_tmp127_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h16)) begin
										r_sys_tmp128_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp129_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp130_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp131_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp132_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp133_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp134_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp135_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp136_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp137_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp138_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp139_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp140_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp141_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp142_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp143_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp144_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp145_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp146_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp147_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp148_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp149_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp150_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp151_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp152_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp153_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp154_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp155_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp156_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp157_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp158_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp159_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp160_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp161_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp162_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp163_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp164_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp165_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp166_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp167_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp168_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp169_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp170_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp171_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp172_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp173_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp174_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp175_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp176_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp177_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp178_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp179_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp180_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp181_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp182_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp183_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp184_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp185_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp186_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp187_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp188_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp189_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp190_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp191_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp192_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp193_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp194_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp195_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp196_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp197_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp198_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp199_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp200_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp201_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp202_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp203_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp204_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp205_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp206_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp207_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp208_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp209_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp210_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp211_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp212_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp213_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp214_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp215_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp216_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp217_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp218_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp219_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp220_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp221_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp222_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp223_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp224_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp225_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp226_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp227_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp228_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp229_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp230_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp231_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp232_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp233_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp234_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp235_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp236_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp237_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp238_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp239_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp240_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp241_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp242_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp243_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp244_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp245_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp246_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp247_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp248_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp249_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp250_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp251_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp252_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp253_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp254_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp255_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp256_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp257_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp258_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp259_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp260_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp261_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp262_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp263_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp264_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp265_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp266_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp267_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp268_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp269_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp270_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp271_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp272_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp273_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp274_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp275_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp276_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp277_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp278_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp279_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp280_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp281_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp282_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp283_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp284_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp285_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp286_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp287_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp288_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp289_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp290_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp291_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp292_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp293_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp294_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp295_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp296_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp297_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp298_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp299_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp300_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp301_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp302_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp303_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp304_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp305_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp306_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp307_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp308_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp309_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp310_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp311_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp312_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp313_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp314_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp315_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp316_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp317_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp318_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp319_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp320_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp321_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp322_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp323_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp324_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp325_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp326_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp327_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp328_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp329_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp330_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp331_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp332_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp333_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp334_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp335_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp336_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp337_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp338_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp339_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp340_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp341_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp342_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp343_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp344_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp345_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp346_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp347_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2) || (r_sys_run_step==9'h21)) begin
										r_sys_tmp348_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
