/*
TimeStamp:	2016/6/3		7:21
*/


module c1_test03(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy	
);

	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 5:0] r_sys_run_phase;
	reg         [ 4:0] r_sys_run_stage;
	reg         [ 6:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 4:0] w_sys_run_stage_p1;
	wire        [ 6:0] w_sys_run_step_p1;
	wire signed [ 8:0] w_fld_u_0_addr_0;
	wire        [31:0] w_fld_u_0_datain_0;
	wire        [31:0] w_fld_u_0_dataout_0;
	wire               w_fld_u_0_r_w_0;
	wire               w_fld_u_0_ce_0;
	reg  signed [ 8:0] r_fld_u_0_addr_1;
	reg         [31:0] r_fld_u_0_datain_1;
	wire        [31:0] w_fld_u_0_dataout_1;
	reg                r_fld_u_0_r_w_1;
	wire               w_fld_u_0_ce_1;
	wire signed [ 8:0] w_fld_uu_1_addr_0;
	wire        [31:0] w_fld_uu_1_datain_0;
	wire        [31:0] w_fld_uu_1_dataout_0;
	wire               w_fld_uu_1_r_w_0;
	wire               w_fld_uu_1_ce_0;
	reg  signed [ 8:0] r_fld_uu_1_addr_1;
	reg         [31:0] r_fld_uu_1_datain_1;
	wire        [31:0] w_fld_uu_1_dataout_1;
	reg                r_fld_uu_1_r_w_1;
	wire               w_fld_uu_1_ce_1;
	reg  signed [31:0] r_run_k_27;
	reg  signed [31:0] r_run_j_28;
	reg  signed [31:0] r_run_n_29;
	reg  signed [31:0] r_run_mx_30;
	reg  signed [31:0] r_run_my_31;
	reg  signed [31:0] r_run_nlast_32;
	reg         [31:0] r_run_dx_33;
	reg         [31:0] r_run_dy_34;
	reg  signed [31:0] r_run_copy0_j_35;
	reg  signed [31:0] r_run_copy0_j_36;
	reg  signed [31:0] r_run_copy1_j_37;
	reg  signed [31:0] r_run_copy2_j_38;
	reg                r_sub19_run_req;
	wire               w_sub19_run_busy;
	wire signed [ 8:0] w_sub19_u_addr;
	reg  signed [ 8:0] r_sub19_u_addr;
	wire        [31:0] w_sub19_u_datain;
	reg         [31:0] r_sub19_u_datain;
	wire        [31:0] w_sub19_u_dataout;
	wire               w_sub19_u_r_w;
	reg                r_sub19_u_r_w;
	wire signed [ 8:0] w_sub19_result_addr;
	reg  signed [ 8:0] r_sub19_result_addr;
	wire        [31:0] w_sub19_result_datain;
	reg         [31:0] r_sub19_result_datain;
	wire        [31:0] w_sub19_result_dataout;
	wire               w_sub19_result_r_w;
	reg                r_sub19_result_r_w;
	reg                r_sub09_run_req;
	wire               w_sub09_run_busy;
	wire signed [ 8:0] w_sub09_u_addr;
	reg  signed [ 8:0] r_sub09_u_addr;
	wire        [31:0] w_sub09_u_datain;
	reg         [31:0] r_sub09_u_datain;
	wire        [31:0] w_sub09_u_dataout;
	wire               w_sub09_u_r_w;
	reg                r_sub09_u_r_w;
	wire signed [ 8:0] w_sub09_result_addr;
	reg  signed [ 8:0] r_sub09_result_addr;
	wire        [31:0] w_sub09_result_datain;
	reg         [31:0] r_sub09_result_datain;
	wire        [31:0] w_sub09_result_dataout;
	wire               w_sub09_result_r_w;
	reg                r_sub09_result_r_w;
	reg                r_sub08_run_req;
	wire               w_sub08_run_busy;
	wire signed [ 8:0] w_sub08_u_addr;
	reg  signed [ 8:0] r_sub08_u_addr;
	wire        [31:0] w_sub08_u_datain;
	reg         [31:0] r_sub08_u_datain;
	wire        [31:0] w_sub08_u_dataout;
	wire               w_sub08_u_r_w;
	reg                r_sub08_u_r_w;
	wire signed [ 8:0] w_sub08_result_addr;
	reg  signed [ 8:0] r_sub08_result_addr;
	wire        [31:0] w_sub08_result_datain;
	reg         [31:0] r_sub08_result_datain;
	wire        [31:0] w_sub08_result_dataout;
	wire               w_sub08_result_r_w;
	reg                r_sub08_result_r_w;
	reg                r_sub24_run_req;
	wire               w_sub24_run_busy;
	wire signed [ 8:0] w_sub24_u_addr;
	reg  signed [ 8:0] r_sub24_u_addr;
	wire        [31:0] w_sub24_u_datain;
	reg         [31:0] r_sub24_u_datain;
	wire        [31:0] w_sub24_u_dataout;
	wire               w_sub24_u_r_w;
	reg                r_sub24_u_r_w;
	wire signed [ 8:0] w_sub24_result_addr;
	reg  signed [ 8:0] r_sub24_result_addr;
	wire        [31:0] w_sub24_result_datain;
	reg         [31:0] r_sub24_result_datain;
	wire        [31:0] w_sub24_result_dataout;
	wire               w_sub24_result_r_w;
	reg                r_sub24_result_r_w;
	reg                r_sub22_run_req;
	wire               w_sub22_run_busy;
	wire signed [ 8:0] w_sub22_u_addr;
	reg  signed [ 8:0] r_sub22_u_addr;
	wire        [31:0] w_sub22_u_datain;
	reg         [31:0] r_sub22_u_datain;
	wire        [31:0] w_sub22_u_dataout;
	wire               w_sub22_u_r_w;
	reg                r_sub22_u_r_w;
	wire signed [ 8:0] w_sub22_result_addr;
	reg  signed [ 8:0] r_sub22_result_addr;
	wire        [31:0] w_sub22_result_datain;
	reg         [31:0] r_sub22_result_datain;
	wire        [31:0] w_sub22_result_dataout;
	wire               w_sub22_result_r_w;
	reg                r_sub22_result_r_w;
	reg                r_sub23_run_req;
	wire               w_sub23_run_busy;
	wire signed [ 8:0] w_sub23_u_addr;
	reg  signed [ 8:0] r_sub23_u_addr;
	wire        [31:0] w_sub23_u_datain;
	reg         [31:0] r_sub23_u_datain;
	wire        [31:0] w_sub23_u_dataout;
	wire               w_sub23_u_r_w;
	reg                r_sub23_u_r_w;
	wire signed [ 8:0] w_sub23_result_addr;
	reg  signed [ 8:0] r_sub23_result_addr;
	wire        [31:0] w_sub23_result_datain;
	reg         [31:0] r_sub23_result_datain;
	wire        [31:0] w_sub23_result_dataout;
	wire               w_sub23_result_r_w;
	reg                r_sub23_result_r_w;
	reg                r_sub12_run_req;
	wire               w_sub12_run_busy;
	wire signed [ 8:0] w_sub12_u_addr;
	reg  signed [ 8:0] r_sub12_u_addr;
	wire        [31:0] w_sub12_u_datain;
	reg         [31:0] r_sub12_u_datain;
	wire        [31:0] w_sub12_u_dataout;
	wire               w_sub12_u_r_w;
	reg                r_sub12_u_r_w;
	wire signed [ 8:0] w_sub12_result_addr;
	reg  signed [ 8:0] r_sub12_result_addr;
	wire        [31:0] w_sub12_result_datain;
	reg         [31:0] r_sub12_result_datain;
	wire        [31:0] w_sub12_result_dataout;
	wire               w_sub12_result_r_w;
	reg                r_sub12_result_r_w;
	reg                r_sub03_run_req;
	wire               w_sub03_run_busy;
	wire signed [ 8:0] w_sub03_u_addr;
	reg  signed [ 8:0] r_sub03_u_addr;
	wire        [31:0] w_sub03_u_datain;
	reg         [31:0] r_sub03_u_datain;
	wire        [31:0] w_sub03_u_dataout;
	wire               w_sub03_u_r_w;
	reg                r_sub03_u_r_w;
	wire signed [ 8:0] w_sub03_result_addr;
	reg  signed [ 8:0] r_sub03_result_addr;
	wire        [31:0] w_sub03_result_datain;
	reg         [31:0] r_sub03_result_datain;
	wire        [31:0] w_sub03_result_dataout;
	wire               w_sub03_result_r_w;
	reg                r_sub03_result_r_w;
	reg                r_sub02_run_req;
	wire               w_sub02_run_busy;
	wire signed [ 8:0] w_sub02_u_addr;
	reg  signed [ 8:0] r_sub02_u_addr;
	wire        [31:0] w_sub02_u_datain;
	reg         [31:0] r_sub02_u_datain;
	wire        [31:0] w_sub02_u_dataout;
	wire               w_sub02_u_r_w;
	reg                r_sub02_u_r_w;
	wire signed [ 8:0] w_sub02_result_addr;
	reg  signed [ 8:0] r_sub02_result_addr;
	wire        [31:0] w_sub02_result_datain;
	reg         [31:0] r_sub02_result_datain;
	wire        [31:0] w_sub02_result_dataout;
	wire               w_sub02_result_r_w;
	reg                r_sub02_result_r_w;
	reg                r_sub11_run_req;
	wire               w_sub11_run_busy;
	wire signed [ 8:0] w_sub11_u_addr;
	reg  signed [ 8:0] r_sub11_u_addr;
	wire        [31:0] w_sub11_u_datain;
	reg         [31:0] r_sub11_u_datain;
	wire        [31:0] w_sub11_u_dataout;
	wire               w_sub11_u_r_w;
	reg                r_sub11_u_r_w;
	wire signed [ 8:0] w_sub11_result_addr;
	reg  signed [ 8:0] r_sub11_result_addr;
	wire        [31:0] w_sub11_result_datain;
	reg         [31:0] r_sub11_result_datain;
	wire        [31:0] w_sub11_result_dataout;
	wire               w_sub11_result_r_w;
	reg                r_sub11_result_r_w;
	reg                r_sub14_run_req;
	wire               w_sub14_run_busy;
	wire signed [ 8:0] w_sub14_u_addr;
	reg  signed [ 8:0] r_sub14_u_addr;
	wire        [31:0] w_sub14_u_datain;
	reg         [31:0] r_sub14_u_datain;
	wire        [31:0] w_sub14_u_dataout;
	wire               w_sub14_u_r_w;
	reg                r_sub14_u_r_w;
	wire signed [ 8:0] w_sub14_result_addr;
	reg  signed [ 8:0] r_sub14_result_addr;
	wire        [31:0] w_sub14_result_datain;
	reg         [31:0] r_sub14_result_datain;
	wire        [31:0] w_sub14_result_dataout;
	wire               w_sub14_result_r_w;
	reg                r_sub14_result_r_w;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [ 8:0] w_sub01_u_addr;
	reg  signed [ 8:0] r_sub01_u_addr;
	wire        [31:0] w_sub01_u_datain;
	reg         [31:0] r_sub01_u_datain;
	wire        [31:0] w_sub01_u_dataout;
	wire               w_sub01_u_r_w;
	reg                r_sub01_u_r_w;
	wire signed [ 8:0] w_sub01_result_addr;
	reg  signed [ 8:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [ 8:0] w_sub00_u_addr;
	reg  signed [ 8:0] r_sub00_u_addr;
	wire        [31:0] w_sub00_u_datain;
	reg         [31:0] r_sub00_u_datain;
	wire        [31:0] w_sub00_u_dataout;
	wire               w_sub00_u_r_w;
	reg                r_sub00_u_r_w;
	wire signed [ 8:0] w_sub00_result_addr;
	reg  signed [ 8:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	reg                r_sub13_run_req;
	wire               w_sub13_run_busy;
	wire signed [ 8:0] w_sub13_u_addr;
	reg  signed [ 8:0] r_sub13_u_addr;
	wire        [31:0] w_sub13_u_datain;
	reg         [31:0] r_sub13_u_datain;
	wire        [31:0] w_sub13_u_dataout;
	wire               w_sub13_u_r_w;
	reg                r_sub13_u_r_w;
	wire signed [ 8:0] w_sub13_result_addr;
	reg  signed [ 8:0] r_sub13_result_addr;
	wire        [31:0] w_sub13_result_datain;
	reg         [31:0] r_sub13_result_datain;
	wire        [31:0] w_sub13_result_dataout;
	wire               w_sub13_result_r_w;
	reg                r_sub13_result_r_w;
	reg                r_sub07_run_req;
	wire               w_sub07_run_busy;
	wire signed [ 8:0] w_sub07_u_addr;
	reg  signed [ 8:0] r_sub07_u_addr;
	wire        [31:0] w_sub07_u_datain;
	reg         [31:0] r_sub07_u_datain;
	wire        [31:0] w_sub07_u_dataout;
	wire               w_sub07_u_r_w;
	reg                r_sub07_u_r_w;
	wire signed [ 8:0] w_sub07_result_addr;
	reg  signed [ 8:0] r_sub07_result_addr;
	wire        [31:0] w_sub07_result_datain;
	reg         [31:0] r_sub07_result_datain;
	wire        [31:0] w_sub07_result_dataout;
	wire               w_sub07_result_r_w;
	reg                r_sub07_result_r_w;
	reg                r_sub16_run_req;
	wire               w_sub16_run_busy;
	wire signed [ 8:0] w_sub16_u_addr;
	reg  signed [ 8:0] r_sub16_u_addr;
	wire        [31:0] w_sub16_u_datain;
	reg         [31:0] r_sub16_u_datain;
	wire        [31:0] w_sub16_u_dataout;
	wire               w_sub16_u_r_w;
	reg                r_sub16_u_r_w;
	wire signed [ 8:0] w_sub16_result_addr;
	reg  signed [ 8:0] r_sub16_result_addr;
	wire        [31:0] w_sub16_result_datain;
	reg         [31:0] r_sub16_result_datain;
	wire        [31:0] w_sub16_result_dataout;
	wire               w_sub16_result_r_w;
	reg                r_sub16_result_r_w;
	reg                r_sub06_run_req;
	wire               w_sub06_run_busy;
	wire signed [ 8:0] w_sub06_u_addr;
	reg  signed [ 8:0] r_sub06_u_addr;
	wire        [31:0] w_sub06_u_datain;
	reg         [31:0] r_sub06_u_datain;
	wire        [31:0] w_sub06_u_dataout;
	wire               w_sub06_u_r_w;
	reg                r_sub06_u_r_w;
	wire signed [ 8:0] w_sub06_result_addr;
	reg  signed [ 8:0] r_sub06_result_addr;
	wire        [31:0] w_sub06_result_datain;
	reg         [31:0] r_sub06_result_datain;
	wire        [31:0] w_sub06_result_dataout;
	wire               w_sub06_result_r_w;
	reg                r_sub06_result_r_w;
	reg                r_sub15_run_req;
	wire               w_sub15_run_busy;
	wire signed [ 8:0] w_sub15_u_addr;
	reg  signed [ 8:0] r_sub15_u_addr;
	wire        [31:0] w_sub15_u_datain;
	reg         [31:0] r_sub15_u_datain;
	wire        [31:0] w_sub15_u_dataout;
	wire               w_sub15_u_r_w;
	reg                r_sub15_u_r_w;
	wire signed [ 8:0] w_sub15_result_addr;
	reg  signed [ 8:0] r_sub15_result_addr;
	wire        [31:0] w_sub15_result_datain;
	reg         [31:0] r_sub15_result_datain;
	wire        [31:0] w_sub15_result_dataout;
	wire               w_sub15_result_r_w;
	reg                r_sub15_result_r_w;
	reg                r_sub05_run_req;
	wire               w_sub05_run_busy;
	wire signed [ 8:0] w_sub05_u_addr;
	reg  signed [ 8:0] r_sub05_u_addr;
	wire        [31:0] w_sub05_u_datain;
	reg         [31:0] r_sub05_u_datain;
	wire        [31:0] w_sub05_u_dataout;
	wire               w_sub05_u_r_w;
	reg                r_sub05_u_r_w;
	wire signed [ 8:0] w_sub05_q_addr;
	reg  signed [ 8:0] r_sub05_q_addr;
	wire        [31:0] w_sub05_q_datain;
	reg         [31:0] r_sub05_q_datain;
	wire        [31:0] w_sub05_q_dataout;
	wire               w_sub05_q_r_w;
	reg                r_sub05_q_r_w;
	wire signed [ 8:0] w_sub05_result_addr;
	reg  signed [ 8:0] r_sub05_result_addr;
	wire        [31:0] w_sub05_result_datain;
	reg         [31:0] r_sub05_result_datain;
	wire        [31:0] w_sub05_result_dataout;
	wire               w_sub05_result_r_w;
	reg                r_sub05_result_r_w;
	reg                r_sub18_run_req;
	wire               w_sub18_run_busy;
	wire signed [ 8:0] w_sub18_u_addr;
	reg  signed [ 8:0] r_sub18_u_addr;
	wire        [31:0] w_sub18_u_datain;
	reg         [31:0] r_sub18_u_datain;
	wire        [31:0] w_sub18_u_dataout;
	wire               w_sub18_u_r_w;
	reg                r_sub18_u_r_w;
	wire signed [ 8:0] w_sub18_result_addr;
	reg  signed [ 8:0] r_sub18_result_addr;
	wire        [31:0] w_sub18_result_datain;
	reg         [31:0] r_sub18_result_datain;
	wire        [31:0] w_sub18_result_dataout;
	wire               w_sub18_result_r_w;
	reg                r_sub18_result_r_w;
	reg                r_sub04_run_req;
	wire               w_sub04_run_busy;
	wire signed [ 8:0] w_sub04_u_addr;
	reg  signed [ 8:0] r_sub04_u_addr;
	wire        [31:0] w_sub04_u_datain;
	reg         [31:0] r_sub04_u_datain;
	wire        [31:0] w_sub04_u_dataout;
	wire               w_sub04_u_r_w;
	reg                r_sub04_u_r_w;
	wire signed [ 8:0] w_sub04_result_addr;
	reg  signed [ 8:0] r_sub04_result_addr;
	wire        [31:0] w_sub04_result_datain;
	reg         [31:0] r_sub04_result_datain;
	wire        [31:0] w_sub04_result_dataout;
	wire               w_sub04_result_r_w;
	reg                r_sub04_result_r_w;
	reg                r_sub17_run_req;
	wire               w_sub17_run_busy;
	wire signed [ 8:0] w_sub17_u_addr;
	reg  signed [ 8:0] r_sub17_u_addr;
	wire        [31:0] w_sub17_u_datain;
	reg         [31:0] r_sub17_u_datain;
	wire        [31:0] w_sub17_u_dataout;
	wire               w_sub17_u_r_w;
	reg                r_sub17_u_r_w;
	wire signed [ 8:0] w_sub17_result_addr;
	reg  signed [ 8:0] r_sub17_result_addr;
	wire        [31:0] w_sub17_result_datain;
	reg         [31:0] r_sub17_result_datain;
	wire        [31:0] w_sub17_result_dataout;
	wire               w_sub17_result_r_w;
	reg                r_sub17_result_r_w;
	reg                r_sub10_run_req;
	wire               w_sub10_run_busy;
	wire signed [ 8:0] w_sub10_u_addr;
	reg  signed [ 8:0] r_sub10_u_addr;
	wire        [31:0] w_sub10_u_datain;
	reg         [31:0] r_sub10_u_datain;
	wire        [31:0] w_sub10_u_dataout;
	wire               w_sub10_u_r_w;
	reg                r_sub10_u_r_w;
	wire signed [ 8:0] w_sub10_result_addr;
	reg  signed [ 8:0] r_sub10_result_addr;
	wire        [31:0] w_sub10_result_datain;
	reg         [31:0] r_sub10_result_datain;
	wire        [31:0] w_sub10_result_dataout;
	wire               w_sub10_result_r_w;
	reg                r_sub10_result_r_w;
	reg                r_sub20_run_req;
	wire               w_sub20_run_busy;
	wire signed [ 8:0] w_sub20_u_addr;
	reg  signed [ 8:0] r_sub20_u_addr;
	wire        [31:0] w_sub20_u_datain;
	reg         [31:0] r_sub20_u_datain;
	wire        [31:0] w_sub20_u_dataout;
	wire               w_sub20_u_r_w;
	reg                r_sub20_u_r_w;
	wire signed [ 8:0] w_sub20_result_addr;
	reg  signed [ 8:0] r_sub20_result_addr;
	wire        [31:0] w_sub20_result_datain;
	reg         [31:0] r_sub20_result_datain;
	wire        [31:0] w_sub20_result_dataout;
	wire               w_sub20_result_r_w;
	reg                r_sub20_result_r_w;
	reg                r_sub21_run_req;
	wire               w_sub21_run_busy;
	wire signed [ 8:0] w_sub21_u_addr;
	reg  signed [ 8:0] r_sub21_u_addr;
	wire        [31:0] w_sub21_u_datain;
	reg         [31:0] r_sub21_u_datain;
	wire        [31:0] w_sub21_u_dataout;
	wire               w_sub21_u_r_w;
	reg                r_sub21_u_r_w;
	wire signed [ 8:0] w_sub21_q_addr;
	reg  signed [ 8:0] r_sub21_q_addr;
	wire        [31:0] w_sub21_q_datain;
	reg         [31:0] r_sub21_q_datain;
	wire        [31:0] w_sub21_q_dataout;
	wire               w_sub21_q_r_w;
	reg                r_sub21_q_r_w;
	wire signed [ 8:0] w_sub21_result_addr;
	reg  signed [ 8:0] r_sub21_result_addr;
	wire        [31:0] w_sub21_result_datain;
	reg         [31:0] r_sub21_result_datain;
	wire        [31:0] w_sub21_result_dataout;
	wire               w_sub21_result_r_w;
	reg                r_sub21_result_r_w;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg         [31:0] r_sys_tmp4_float;
	reg         [31:0] r_sys_tmp5_float;
	reg         [31:0] r_sys_tmp6_float;
	reg         [31:0] r_sys_tmp7_float;
	reg         [31:0] r_sys_tmp8_float;
	reg         [31:0] r_sys_tmp9_float;
	reg         [31:0] r_sys_tmp10_float;
	reg         [31:0] r_sys_tmp11_float;
	reg         [31:0] r_sys_tmp12_float;
	reg         [31:0] r_sys_tmp13_float;
	reg         [31:0] r_sys_tmp14_float;
	reg         [31:0] r_sys_tmp15_float;
	reg         [31:0] r_sys_tmp16_float;
	reg         [31:0] r_sys_tmp17_float;
	reg         [31:0] r_sys_tmp18_float;
	reg         [31:0] r_sys_tmp19_float;
	reg         [31:0] r_sys_tmp20_float;
	reg         [31:0] r_sys_tmp21_float;
	reg         [31:0] r_sys_tmp22_float;
	reg         [31:0] r_sys_tmp23_float;
	reg         [31:0] r_sys_tmp24_float;
	reg         [31:0] r_sys_tmp25_float;
	reg         [31:0] r_sys_tmp26_float;
	reg         [31:0] r_sys_tmp27_float;
	reg         [31:0] r_sys_tmp28_float;
	reg         [31:0] r_sys_tmp29_float;
	reg         [31:0] r_sys_tmp30_float;
	reg         [31:0] r_sys_tmp31_float;
	reg         [31:0] r_sys_tmp32_float;
	reg         [31:0] r_sys_tmp33_float;
	reg         [31:0] r_sys_tmp34_float;
	reg         [31:0] r_sys_tmp35_float;
	reg         [31:0] r_sys_tmp36_float;
	reg         [31:0] r_sys_tmp37_float;
	reg         [31:0] r_sys_tmp38_float;
	reg         [31:0] r_sys_tmp39_float;
	reg         [31:0] r_sys_tmp40_float;
	reg         [31:0] r_sys_tmp41_float;
	reg         [31:0] r_sys_tmp42_float;
	reg         [31:0] r_sys_tmp43_float;
	reg         [31:0] r_sys_tmp44_float;
	reg         [31:0] r_sys_tmp45_float;
	reg         [31:0] r_sys_tmp46_float;
	reg         [31:0] r_sys_tmp47_float;
	reg         [31:0] r_sys_tmp48_float;
	reg         [31:0] r_sys_tmp49_float;
	reg         [31:0] r_sys_tmp50_float;
	reg         [31:0] r_sys_tmp51_float;
	reg         [31:0] r_sys_tmp52_float;
	wire signed [31:0] w_sys_tmp1;
	wire        [31:0] w_sys_tmp3;
	wire signed [31:0] w_sys_tmp5;
	wire               w_sys_tmp6;
	wire               w_sys_tmp7;
	wire signed [31:0] w_sys_tmp8;
	wire               w_sys_tmp9;
	wire               w_sys_tmp10;
	wire signed [31:0] w_sys_tmp13;
	wire signed [31:0] w_sys_tmp14;
	wire signed [31:0] w_sys_tmp15;
	wire        [31:0] w_sys_tmp16;
	wire signed [31:0] w_sys_tmp18;
	wire signed [31:0] w_sys_tmp19;
	wire signed [31:0] w_sys_tmp22;
	wire signed [31:0] w_sys_tmp23;
	wire               w_sys_tmp96;
	wire               w_sys_tmp97;
	wire signed [31:0] w_sys_tmp98;
	wire               w_sys_tmp99;
	wire               w_sys_tmp100;
	wire signed [31:0] w_sys_tmp103;
	wire signed [31:0] w_sys_tmp104;
	wire        [31:0] w_sys_tmp105;
	wire signed [31:0] w_sys_tmp107;
	wire signed [31:0] w_sys_tmp108;
	wire        [31:0] w_sys_tmp110;
	wire signed [31:0] w_sys_tmp112;
	wire signed [31:0] w_sys_tmp113;
	wire        [31:0] w_sys_tmp115;
	wire signed [31:0] w_sys_tmp117;
	wire signed [31:0] w_sys_tmp118;
	wire signed [31:0] w_sys_tmp121;
	wire signed [31:0] w_sys_tmp122;
	wire signed [31:0] w_sys_tmp123;
	wire signed [31:0] w_sys_tmp124;
	wire               w_sys_tmp263;
	wire               w_sys_tmp264;
	wire signed [31:0] w_sys_tmp265;
	wire signed [31:0] w_sys_tmp268;
	wire signed [31:0] w_sys_tmp269;
	wire        [31:0] w_sys_tmp270;
	wire signed [31:0] w_sys_tmp274;
	wire signed [31:0] w_sys_tmp275;
	wire signed [31:0] w_sys_tmp280;
	wire signed [31:0] w_sys_tmp281;
	wire signed [31:0] w_sys_tmp286;
	wire signed [31:0] w_sys_tmp287;
	wire signed [31:0] w_sys_tmp292;
	wire signed [31:0] w_sys_tmp293;
	wire signed [31:0] w_sys_tmp310;
	wire signed [31:0] w_sys_tmp311;
	wire signed [31:0] w_sys_tmp316;
	wire signed [31:0] w_sys_tmp317;
	wire signed [31:0] w_sys_tmp322;
	wire signed [31:0] w_sys_tmp323;
	wire signed [31:0] w_sys_tmp328;
	wire signed [31:0] w_sys_tmp329;
	wire signed [31:0] w_sys_tmp346;
	wire signed [31:0] w_sys_tmp347;
	wire signed [31:0] w_sys_tmp352;
	wire signed [31:0] w_sys_tmp353;
	wire signed [31:0] w_sys_tmp358;
	wire signed [31:0] w_sys_tmp359;
	wire signed [31:0] w_sys_tmp364;
	wire signed [31:0] w_sys_tmp365;
	wire signed [31:0] w_sys_tmp382;
	wire signed [31:0] w_sys_tmp383;
	wire signed [31:0] w_sys_tmp388;
	wire signed [31:0] w_sys_tmp389;
	wire signed [31:0] w_sys_tmp394;
	wire signed [31:0] w_sys_tmp395;
	wire signed [31:0] w_sys_tmp400;
	wire signed [31:0] w_sys_tmp401;
	wire signed [31:0] w_sys_tmp418;
	wire signed [31:0] w_sys_tmp419;
	wire signed [31:0] w_sys_tmp424;
	wire signed [31:0] w_sys_tmp425;
	wire signed [31:0] w_sys_tmp430;
	wire signed [31:0] w_sys_tmp431;
	wire signed [31:0] w_sys_tmp436;
	wire signed [31:0] w_sys_tmp437;
	wire signed [31:0] w_sys_tmp441;
	wire signed [31:0] w_sys_tmp442;
	wire               w_sys_tmp443;
	wire               w_sys_tmp444;
	wire signed [31:0] w_sys_tmp445;
	wire signed [31:0] w_sys_tmp448;
	wire signed [31:0] w_sys_tmp449;
	wire        [31:0] w_sys_tmp450;
	wire signed [31:0] w_sys_tmp454;
	wire signed [31:0] w_sys_tmp455;
	wire signed [31:0] w_sys_tmp460;
	wire signed [31:0] w_sys_tmp461;
	wire signed [31:0] w_sys_tmp466;
	wire signed [31:0] w_sys_tmp467;
	wire signed [31:0] w_sys_tmp472;
	wire signed [31:0] w_sys_tmp473;
	wire signed [31:0] w_sys_tmp490;
	wire signed [31:0] w_sys_tmp491;
	wire signed [31:0] w_sys_tmp496;
	wire signed [31:0] w_sys_tmp497;
	wire signed [31:0] w_sys_tmp502;
	wire signed [31:0] w_sys_tmp503;
	wire signed [31:0] w_sys_tmp508;
	wire signed [31:0] w_sys_tmp509;
	wire signed [31:0] w_sys_tmp526;
	wire signed [31:0] w_sys_tmp527;
	wire signed [31:0] w_sys_tmp532;
	wire signed [31:0] w_sys_tmp533;
	wire signed [31:0] w_sys_tmp538;
	wire signed [31:0] w_sys_tmp539;
	wire signed [31:0] w_sys_tmp544;
	wire signed [31:0] w_sys_tmp545;
	wire signed [31:0] w_sys_tmp562;
	wire signed [31:0] w_sys_tmp563;
	wire signed [31:0] w_sys_tmp568;
	wire signed [31:0] w_sys_tmp569;
	wire signed [31:0] w_sys_tmp574;
	wire signed [31:0] w_sys_tmp575;
	wire signed [31:0] w_sys_tmp580;
	wire signed [31:0] w_sys_tmp581;
	wire signed [31:0] w_sys_tmp598;
	wire signed [31:0] w_sys_tmp599;
	wire signed [31:0] w_sys_tmp604;
	wire signed [31:0] w_sys_tmp605;
	wire signed [31:0] w_sys_tmp610;
	wire signed [31:0] w_sys_tmp611;
	wire signed [31:0] w_sys_tmp616;
	wire signed [31:0] w_sys_tmp617;
	wire signed [31:0] w_sys_tmp622;
	wire signed [31:0] w_sys_tmp623;
	wire signed [31:0] w_sys_tmp628;
	wire signed [31:0] w_sys_tmp629;
	wire signed [31:0] w_sys_tmp634;
	wire signed [31:0] w_sys_tmp635;
	wire signed [31:0] w_sys_tmp640;
	wire signed [31:0] w_sys_tmp641;
	wire signed [31:0] w_sys_tmp646;
	wire signed [31:0] w_sys_tmp647;
	wire signed [31:0] w_sys_tmp664;
	wire signed [31:0] w_sys_tmp665;
	wire signed [31:0] w_sys_tmp670;
	wire signed [31:0] w_sys_tmp671;
	wire signed [31:0] w_sys_tmp676;
	wire signed [31:0] w_sys_tmp677;
	wire signed [31:0] w_sys_tmp682;
	wire signed [31:0] w_sys_tmp683;
	wire signed [31:0] w_sys_tmp700;
	wire signed [31:0] w_sys_tmp701;
	wire signed [31:0] w_sys_tmp706;
	wire signed [31:0] w_sys_tmp707;
	wire signed [31:0] w_sys_tmp712;
	wire signed [31:0] w_sys_tmp713;
	wire signed [31:0] w_sys_tmp718;
	wire signed [31:0] w_sys_tmp719;
	wire signed [31:0] w_sys_tmp736;
	wire signed [31:0] w_sys_tmp737;
	wire signed [31:0] w_sys_tmp742;
	wire signed [31:0] w_sys_tmp743;
	wire signed [31:0] w_sys_tmp748;
	wire signed [31:0] w_sys_tmp749;
	wire signed [31:0] w_sys_tmp754;
	wire signed [31:0] w_sys_tmp755;
	wire signed [31:0] w_sys_tmp772;
	wire signed [31:0] w_sys_tmp773;
	wire signed [31:0] w_sys_tmp778;
	wire signed [31:0] w_sys_tmp779;
	wire signed [31:0] w_sys_tmp784;
	wire signed [31:0] w_sys_tmp785;
	wire signed [31:0] w_sys_tmp790;
	wire signed [31:0] w_sys_tmp791;
	wire signed [31:0] w_sys_tmp796;
	wire signed [31:0] w_sys_tmp797;
	wire signed [31:0] w_sys_tmp802;
	wire signed [31:0] w_sys_tmp803;
	wire signed [31:0] w_sys_tmp808;
	wire signed [31:0] w_sys_tmp809;
	wire signed [31:0] w_sys_tmp814;
	wire signed [31:0] w_sys_tmp815;
	wire signed [31:0] w_sys_tmp820;
	wire signed [31:0] w_sys_tmp821;
	wire signed [31:0] w_sys_tmp838;
	wire signed [31:0] w_sys_tmp839;
	wire signed [31:0] w_sys_tmp844;
	wire signed [31:0] w_sys_tmp845;
	wire signed [31:0] w_sys_tmp850;
	wire signed [31:0] w_sys_tmp851;
	wire signed [31:0] w_sys_tmp856;
	wire signed [31:0] w_sys_tmp857;
	wire signed [31:0] w_sys_tmp874;
	wire signed [31:0] w_sys_tmp875;
	wire signed [31:0] w_sys_tmp880;
	wire signed [31:0] w_sys_tmp881;
	wire signed [31:0] w_sys_tmp886;
	wire signed [31:0] w_sys_tmp887;
	wire signed [31:0] w_sys_tmp892;
	wire signed [31:0] w_sys_tmp893;
	wire signed [31:0] w_sys_tmp910;
	wire signed [31:0] w_sys_tmp911;
	wire signed [31:0] w_sys_tmp916;
	wire signed [31:0] w_sys_tmp917;
	wire signed [31:0] w_sys_tmp922;
	wire signed [31:0] w_sys_tmp923;
	wire signed [31:0] w_sys_tmp928;
	wire signed [31:0] w_sys_tmp929;
	wire signed [31:0] w_sys_tmp946;
	wire signed [31:0] w_sys_tmp947;
	wire signed [31:0] w_sys_tmp952;
	wire signed [31:0] w_sys_tmp953;
	wire signed [31:0] w_sys_tmp958;
	wire signed [31:0] w_sys_tmp959;
	wire signed [31:0] w_sys_tmp964;
	wire signed [31:0] w_sys_tmp965;
	wire signed [31:0] w_sys_tmp970;
	wire signed [31:0] w_sys_tmp971;
	wire signed [31:0] w_sys_tmp976;
	wire signed [31:0] w_sys_tmp977;
	wire signed [31:0] w_sys_tmp982;
	wire signed [31:0] w_sys_tmp983;
	wire signed [31:0] w_sys_tmp988;
	wire signed [31:0] w_sys_tmp989;
	wire signed [31:0] w_sys_tmp994;
	wire signed [31:0] w_sys_tmp995;
	wire signed [31:0] w_sys_tmp1012;
	wire signed [31:0] w_sys_tmp1013;
	wire signed [31:0] w_sys_tmp1018;
	wire signed [31:0] w_sys_tmp1019;
	wire signed [31:0] w_sys_tmp1024;
	wire signed [31:0] w_sys_tmp1025;
	wire signed [31:0] w_sys_tmp1030;
	wire signed [31:0] w_sys_tmp1031;
	wire signed [31:0] w_sys_tmp1048;
	wire signed [31:0] w_sys_tmp1049;
	wire signed [31:0] w_sys_tmp1054;
	wire signed [31:0] w_sys_tmp1055;
	wire signed [31:0] w_sys_tmp1060;
	wire signed [31:0] w_sys_tmp1061;
	wire signed [31:0] w_sys_tmp1066;
	wire signed [31:0] w_sys_tmp1067;
	wire signed [31:0] w_sys_tmp1084;
	wire signed [31:0] w_sys_tmp1085;
	wire signed [31:0] w_sys_tmp1090;
	wire signed [31:0] w_sys_tmp1091;
	wire signed [31:0] w_sys_tmp1096;
	wire signed [31:0] w_sys_tmp1097;
	wire signed [31:0] w_sys_tmp1102;
	wire signed [31:0] w_sys_tmp1103;
	wire signed [31:0] w_sys_tmp1120;
	wire signed [31:0] w_sys_tmp1121;
	wire signed [31:0] w_sys_tmp1126;
	wire signed [31:0] w_sys_tmp1127;
	wire signed [31:0] w_sys_tmp1132;
	wire signed [31:0] w_sys_tmp1133;
	wire signed [31:0] w_sys_tmp1138;
	wire signed [31:0] w_sys_tmp1139;
	wire signed [31:0] w_sys_tmp1143;
	wire signed [31:0] w_sys_tmp1144;
	wire               w_sys_tmp1145;
	wire               w_sys_tmp1146;
	wire signed [31:0] w_sys_tmp1147;
	wire signed [31:0] w_sys_tmp1150;
	wire signed [31:0] w_sys_tmp1151;
	wire        [31:0] w_sys_tmp1152;
	wire signed [31:0] w_sys_tmp1156;
	wire signed [31:0] w_sys_tmp1157;
	wire signed [31:0] w_sys_tmp1162;
	wire signed [31:0] w_sys_tmp1163;
	wire signed [31:0] w_sys_tmp1168;
	wire signed [31:0] w_sys_tmp1169;
	wire signed [31:0] w_sys_tmp1173;
	wire signed [31:0] w_sys_tmp1174;
	wire signed [31:0] w_sys_tmp1178;
	wire signed [31:0] w_sys_tmp1179;
	wire signed [31:0] w_sys_tmp1183;
	wire signed [31:0] w_sys_tmp1184;
	wire signed [31:0] w_sys_tmp1188;
	wire signed [31:0] w_sys_tmp1189;
	wire signed [31:0] w_sys_tmp1193;
	wire signed [31:0] w_sys_tmp1194;
	wire signed [31:0] w_sys_tmp1198;
	wire signed [31:0] w_sys_tmp1199;
	wire signed [31:0] w_sys_tmp1203;
	wire signed [31:0] w_sys_tmp1204;
	wire signed [31:0] w_sys_tmp1208;
	wire signed [31:0] w_sys_tmp1209;
	wire signed [31:0] w_sys_tmp1213;
	wire signed [31:0] w_sys_tmp1214;
	wire signed [31:0] w_sys_tmp1218;
	wire signed [31:0] w_sys_tmp1219;
	wire signed [31:0] w_sys_tmp1223;
	wire signed [31:0] w_sys_tmp1224;
	wire signed [31:0] w_sys_tmp1228;
	wire signed [31:0] w_sys_tmp1229;
	wire signed [31:0] w_sys_tmp1233;
	wire signed [31:0] w_sys_tmp1234;
	wire signed [31:0] w_sys_tmp1238;
	wire signed [31:0] w_sys_tmp1239;
	wire signed [31:0] w_sys_tmp1243;
	wire signed [31:0] w_sys_tmp1244;
	wire signed [31:0] w_sys_tmp1247;
	wire signed [31:0] w_sys_tmp1248;
	wire               w_sys_tmp1249;
	wire               w_sys_tmp1250;
	wire signed [31:0] w_sys_tmp1251;
	wire signed [31:0] w_sys_tmp1254;
	wire signed [31:0] w_sys_tmp1255;
	wire        [31:0] w_sys_tmp1256;
	wire signed [31:0] w_sys_tmp1260;
	wire signed [31:0] w_sys_tmp1261;
	wire signed [31:0] w_sys_tmp1266;
	wire signed [31:0] w_sys_tmp1267;
	wire signed [31:0] w_sys_tmp1272;
	wire signed [31:0] w_sys_tmp1273;
	wire signed [31:0] w_sys_tmp1277;
	wire signed [31:0] w_sys_tmp1278;
	wire signed [31:0] w_sys_tmp1282;
	wire signed [31:0] w_sys_tmp1283;
	wire signed [31:0] w_sys_tmp1287;
	wire signed [31:0] w_sys_tmp1288;
	wire signed [31:0] w_sys_tmp1292;
	wire signed [31:0] w_sys_tmp1293;
	wire signed [31:0] w_sys_tmp1297;
	wire signed [31:0] w_sys_tmp1298;
	wire signed [31:0] w_sys_tmp1302;
	wire signed [31:0] w_sys_tmp1303;
	wire signed [31:0] w_sys_tmp1307;
	wire signed [31:0] w_sys_tmp1308;
	wire signed [31:0] w_sys_tmp1312;
	wire signed [31:0] w_sys_tmp1313;
	wire signed [31:0] w_sys_tmp1317;
	wire signed [31:0] w_sys_tmp1318;
	wire signed [31:0] w_sys_tmp1322;
	wire signed [31:0] w_sys_tmp1323;
	wire signed [31:0] w_sys_tmp1327;
	wire signed [31:0] w_sys_tmp1328;
	wire signed [31:0] w_sys_tmp1332;
	wire signed [31:0] w_sys_tmp1333;
	wire signed [31:0] w_sys_tmp1337;
	wire signed [31:0] w_sys_tmp1338;
	wire signed [31:0] w_sys_tmp1342;
	wire signed [31:0] w_sys_tmp1343;
	wire signed [31:0] w_sys_tmp1347;
	wire signed [31:0] w_sys_tmp1348;
	wire signed [31:0] w_sys_tmp1351;
	wire signed [31:0] w_sys_tmp1352;
	wire               w_sys_tmp1353;
	wire               w_sys_tmp1354;
	wire signed [31:0] w_sys_tmp1355;
	wire signed [31:0] w_sys_tmp1358;
	wire signed [31:0] w_sys_tmp1359;
	wire        [31:0] w_sys_tmp1360;
	wire signed [31:0] w_sys_tmp1364;
	wire signed [31:0] w_sys_tmp1365;
	wire signed [31:0] w_sys_tmp1370;
	wire signed [31:0] w_sys_tmp1371;
	wire signed [31:0] w_sys_tmp1376;
	wire signed [31:0] w_sys_tmp1377;
	wire signed [31:0] w_sys_tmp1381;
	wire signed [31:0] w_sys_tmp1382;
	wire signed [31:0] w_sys_tmp1386;
	wire signed [31:0] w_sys_tmp1387;
	wire signed [31:0] w_sys_tmp1391;
	wire signed [31:0] w_sys_tmp1392;
	wire signed [31:0] w_sys_tmp1396;
	wire signed [31:0] w_sys_tmp1397;
	wire signed [31:0] w_sys_tmp1401;
	wire signed [31:0] w_sys_tmp1402;
	wire signed [31:0] w_sys_tmp1406;
	wire signed [31:0] w_sys_tmp1407;
	wire signed [31:0] w_sys_tmp1411;
	wire signed [31:0] w_sys_tmp1412;
	wire signed [31:0] w_sys_tmp1416;
	wire signed [31:0] w_sys_tmp1417;
	wire signed [31:0] w_sys_tmp1421;
	wire signed [31:0] w_sys_tmp1422;
	wire signed [31:0] w_sys_tmp1426;
	wire signed [31:0] w_sys_tmp1427;
	wire signed [31:0] w_sys_tmp1431;
	wire signed [31:0] w_sys_tmp1432;
	wire signed [31:0] w_sys_tmp1436;
	wire signed [31:0] w_sys_tmp1437;
	wire signed [31:0] w_sys_tmp1441;
	wire signed [31:0] w_sys_tmp1442;
	wire signed [31:0] w_sys_tmp1446;
	wire signed [31:0] w_sys_tmp1447;
	wire signed [31:0] w_sys_tmp1451;
	wire signed [31:0] w_sys_tmp1452;
	wire signed [31:0] w_sys_tmp1456;
	wire signed [31:0] w_sys_tmp1457;
	wire signed [31:0] w_sys_tmp1461;
	wire signed [31:0] w_sys_tmp1462;
	wire signed [31:0] w_sys_tmp1466;
	wire signed [31:0] w_sys_tmp1467;
	wire signed [31:0] w_sys_tmp1471;
	wire signed [31:0] w_sys_tmp1472;
	wire signed [31:0] w_sys_tmp1476;
	wire signed [31:0] w_sys_tmp1477;
	wire signed [31:0] w_sys_tmp1481;
	wire signed [31:0] w_sys_tmp1482;
	wire signed [31:0] w_sys_tmp1486;
	wire signed [31:0] w_sys_tmp1487;
	wire signed [31:0] w_sys_tmp1491;
	wire signed [31:0] w_sys_tmp1492;
	wire signed [31:0] w_sys_tmp1496;
	wire signed [31:0] w_sys_tmp1497;
	wire signed [31:0] w_sys_tmp1501;
	wire signed [31:0] w_sys_tmp1502;
	wire signed [31:0] w_sys_tmp1506;
	wire signed [31:0] w_sys_tmp1507;
	wire signed [31:0] w_sys_tmp1511;
	wire signed [31:0] w_sys_tmp1512;
	wire signed [31:0] w_sys_tmp1516;
	wire signed [31:0] w_sys_tmp1517;
	wire signed [31:0] w_sys_tmp1521;
	wire signed [31:0] w_sys_tmp1522;
	wire signed [31:0] w_sys_tmp1526;
	wire signed [31:0] w_sys_tmp1527;
	wire signed [31:0] w_sys_tmp1531;
	wire signed [31:0] w_sys_tmp1532;
	wire signed [31:0] w_sys_tmp1536;
	wire signed [31:0] w_sys_tmp1537;
	wire signed [31:0] w_sys_tmp1541;
	wire signed [31:0] w_sys_tmp1542;
	wire signed [31:0] w_sys_tmp1546;
	wire signed [31:0] w_sys_tmp1547;
	wire signed [31:0] w_sys_tmp1551;
	wire signed [31:0] w_sys_tmp1552;
	wire signed [31:0] w_sys_tmp1556;
	wire signed [31:0] w_sys_tmp1557;
	wire signed [31:0] w_sys_tmp1561;
	wire signed [31:0] w_sys_tmp1562;
	wire signed [31:0] w_sys_tmp1566;
	wire signed [31:0] w_sys_tmp1567;
	wire signed [31:0] w_sys_tmp1571;
	wire signed [31:0] w_sys_tmp1572;
	wire signed [31:0] w_sys_tmp1576;
	wire signed [31:0] w_sys_tmp1577;
	wire signed [31:0] w_sys_tmp1581;
	wire signed [31:0] w_sys_tmp1582;
	wire signed [31:0] w_sys_tmp1586;
	wire signed [31:0] w_sys_tmp1587;
	wire signed [31:0] w_sys_tmp1591;
	wire signed [31:0] w_sys_tmp1592;
	wire signed [31:0] w_sys_tmp1596;
	wire signed [31:0] w_sys_tmp1597;
	wire signed [31:0] w_sys_tmp1601;
	wire signed [31:0] w_sys_tmp1602;
	wire signed [31:0] w_sys_tmp1606;
	wire signed [31:0] w_sys_tmp1607;
	wire signed [31:0] w_sys_tmp1611;
	wire signed [31:0] w_sys_tmp1612;
	wire signed [31:0] w_sys_tmp1616;
	wire signed [31:0] w_sys_tmp1617;
	wire signed [31:0] w_sys_tmp1621;
	wire signed [31:0] w_sys_tmp1622;
	wire signed [31:0] w_sys_tmp1626;
	wire signed [31:0] w_sys_tmp1627;
	wire signed [31:0] w_sys_tmp1631;
	wire signed [31:0] w_sys_tmp1632;
	wire signed [31:0] w_sys_tmp1636;
	wire signed [31:0] w_sys_tmp1637;
	wire signed [31:0] w_sys_tmp1641;
	wire signed [31:0] w_sys_tmp1642;
	wire signed [31:0] w_sys_tmp1645;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 5'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 7'h1);
	assign w_fld_u_0_addr_0 = 9'sh0;
	assign w_fld_u_0_datain_0 = 32'h0;
	assign w_fld_u_0_r_w_0 = 1'h0;
	assign w_fld_u_0_ce_0 = w_sys_ce;
	assign w_fld_u_0_ce_1 = w_sys_ce;
	assign w_fld_uu_1_addr_0 = 9'sh0;
	assign w_fld_uu_1_datain_0 = 32'h0;
	assign w_fld_uu_1_r_w_0 = 1'h0;
	assign w_fld_uu_1_ce_0 = w_sys_ce;
	assign w_fld_uu_1_ce_1 = w_sys_ce;
	assign w_sub19_u_addr = ( (|r_sys_processing_methodID) ? r_sub19_u_addr : 9'sh0 ) ;
	assign w_sub19_u_datain = ( (|r_sys_processing_methodID) ? r_sub19_u_datain : 32'h0 ) ;
	assign w_sub19_u_r_w = ( (|r_sys_processing_methodID) ? r_sub19_u_r_w : 1'h0 ) ;
	assign w_sub19_result_addr = ( (|r_sys_processing_methodID) ? r_sub19_result_addr : 9'sh0 ) ;
	assign w_sub19_result_datain = ( (|r_sys_processing_methodID) ? r_sub19_result_datain : 32'h0 ) ;
	assign w_sub19_result_r_w = ( (|r_sys_processing_methodID) ? r_sub19_result_r_w : 1'h0 ) ;
	assign w_sub09_u_addr = ( (|r_sys_processing_methodID) ? r_sub09_u_addr : 9'sh0 ) ;
	assign w_sub09_u_datain = ( (|r_sys_processing_methodID) ? r_sub09_u_datain : 32'h0 ) ;
	assign w_sub09_u_r_w = ( (|r_sys_processing_methodID) ? r_sub09_u_r_w : 1'h0 ) ;
	assign w_sub09_result_addr = ( (|r_sys_processing_methodID) ? r_sub09_result_addr : 9'sh0 ) ;
	assign w_sub09_result_datain = ( (|r_sys_processing_methodID) ? r_sub09_result_datain : 32'h0 ) ;
	assign w_sub09_result_r_w = ( (|r_sys_processing_methodID) ? r_sub09_result_r_w : 1'h0 ) ;
	assign w_sub08_u_addr = ( (|r_sys_processing_methodID) ? r_sub08_u_addr : 9'sh0 ) ;
	assign w_sub08_u_datain = ( (|r_sys_processing_methodID) ? r_sub08_u_datain : 32'h0 ) ;
	assign w_sub08_u_r_w = ( (|r_sys_processing_methodID) ? r_sub08_u_r_w : 1'h0 ) ;
	assign w_sub08_result_addr = ( (|r_sys_processing_methodID) ? r_sub08_result_addr : 9'sh0 ) ;
	assign w_sub08_result_datain = ( (|r_sys_processing_methodID) ? r_sub08_result_datain : 32'h0 ) ;
	assign w_sub08_result_r_w = ( (|r_sys_processing_methodID) ? r_sub08_result_r_w : 1'h0 ) ;
	assign w_sub24_u_addr = ( (|r_sys_processing_methodID) ? r_sub24_u_addr : 9'sh0 ) ;
	assign w_sub24_u_datain = ( (|r_sys_processing_methodID) ? r_sub24_u_datain : 32'h0 ) ;
	assign w_sub24_u_r_w = ( (|r_sys_processing_methodID) ? r_sub24_u_r_w : 1'h0 ) ;
	assign w_sub24_result_addr = ( (|r_sys_processing_methodID) ? r_sub24_result_addr : 9'sh0 ) ;
	assign w_sub24_result_datain = ( (|r_sys_processing_methodID) ? r_sub24_result_datain : 32'h0 ) ;
	assign w_sub24_result_r_w = ( (|r_sys_processing_methodID) ? r_sub24_result_r_w : 1'h0 ) ;
	assign w_sub22_u_addr = ( (|r_sys_processing_methodID) ? r_sub22_u_addr : 9'sh0 ) ;
	assign w_sub22_u_datain = ( (|r_sys_processing_methodID) ? r_sub22_u_datain : 32'h0 ) ;
	assign w_sub22_u_r_w = ( (|r_sys_processing_methodID) ? r_sub22_u_r_w : 1'h0 ) ;
	assign w_sub22_result_addr = ( (|r_sys_processing_methodID) ? r_sub22_result_addr : 9'sh0 ) ;
	assign w_sub22_result_datain = ( (|r_sys_processing_methodID) ? r_sub22_result_datain : 32'h0 ) ;
	assign w_sub22_result_r_w = ( (|r_sys_processing_methodID) ? r_sub22_result_r_w : 1'h0 ) ;
	assign w_sub23_u_addr = ( (|r_sys_processing_methodID) ? r_sub23_u_addr : 9'sh0 ) ;
	assign w_sub23_u_datain = ( (|r_sys_processing_methodID) ? r_sub23_u_datain : 32'h0 ) ;
	assign w_sub23_u_r_w = ( (|r_sys_processing_methodID) ? r_sub23_u_r_w : 1'h0 ) ;
	assign w_sub23_result_addr = ( (|r_sys_processing_methodID) ? r_sub23_result_addr : 9'sh0 ) ;
	assign w_sub23_result_datain = ( (|r_sys_processing_methodID) ? r_sub23_result_datain : 32'h0 ) ;
	assign w_sub23_result_r_w = ( (|r_sys_processing_methodID) ? r_sub23_result_r_w : 1'h0 ) ;
	assign w_sub12_u_addr = ( (|r_sys_processing_methodID) ? r_sub12_u_addr : 9'sh0 ) ;
	assign w_sub12_u_datain = ( (|r_sys_processing_methodID) ? r_sub12_u_datain : 32'h0 ) ;
	assign w_sub12_u_r_w = ( (|r_sys_processing_methodID) ? r_sub12_u_r_w : 1'h0 ) ;
	assign w_sub12_result_addr = ( (|r_sys_processing_methodID) ? r_sub12_result_addr : 9'sh0 ) ;
	assign w_sub12_result_datain = ( (|r_sys_processing_methodID) ? r_sub12_result_datain : 32'h0 ) ;
	assign w_sub12_result_r_w = ( (|r_sys_processing_methodID) ? r_sub12_result_r_w : 1'h0 ) ;
	assign w_sub03_u_addr = ( (|r_sys_processing_methodID) ? r_sub03_u_addr : 9'sh0 ) ;
	assign w_sub03_u_datain = ( (|r_sys_processing_methodID) ? r_sub03_u_datain : 32'h0 ) ;
	assign w_sub03_u_r_w = ( (|r_sys_processing_methodID) ? r_sub03_u_r_w : 1'h0 ) ;
	assign w_sub03_result_addr = ( (|r_sys_processing_methodID) ? r_sub03_result_addr : 9'sh0 ) ;
	assign w_sub03_result_datain = ( (|r_sys_processing_methodID) ? r_sub03_result_datain : 32'h0 ) ;
	assign w_sub03_result_r_w = ( (|r_sys_processing_methodID) ? r_sub03_result_r_w : 1'h0 ) ;
	assign w_sub02_u_addr = ( (|r_sys_processing_methodID) ? r_sub02_u_addr : 9'sh0 ) ;
	assign w_sub02_u_datain = ( (|r_sys_processing_methodID) ? r_sub02_u_datain : 32'h0 ) ;
	assign w_sub02_u_r_w = ( (|r_sys_processing_methodID) ? r_sub02_u_r_w : 1'h0 ) ;
	assign w_sub02_result_addr = ( (|r_sys_processing_methodID) ? r_sub02_result_addr : 9'sh0 ) ;
	assign w_sub02_result_datain = ( (|r_sys_processing_methodID) ? r_sub02_result_datain : 32'h0 ) ;
	assign w_sub02_result_r_w = ( (|r_sys_processing_methodID) ? r_sub02_result_r_w : 1'h0 ) ;
	assign w_sub11_u_addr = ( (|r_sys_processing_methodID) ? r_sub11_u_addr : 9'sh0 ) ;
	assign w_sub11_u_datain = ( (|r_sys_processing_methodID) ? r_sub11_u_datain : 32'h0 ) ;
	assign w_sub11_u_r_w = ( (|r_sys_processing_methodID) ? r_sub11_u_r_w : 1'h0 ) ;
	assign w_sub11_result_addr = ( (|r_sys_processing_methodID) ? r_sub11_result_addr : 9'sh0 ) ;
	assign w_sub11_result_datain = ( (|r_sys_processing_methodID) ? r_sub11_result_datain : 32'h0 ) ;
	assign w_sub11_result_r_w = ( (|r_sys_processing_methodID) ? r_sub11_result_r_w : 1'h0 ) ;
	assign w_sub14_u_addr = ( (|r_sys_processing_methodID) ? r_sub14_u_addr : 9'sh0 ) ;
	assign w_sub14_u_datain = ( (|r_sys_processing_methodID) ? r_sub14_u_datain : 32'h0 ) ;
	assign w_sub14_u_r_w = ( (|r_sys_processing_methodID) ? r_sub14_u_r_w : 1'h0 ) ;
	assign w_sub14_result_addr = ( (|r_sys_processing_methodID) ? r_sub14_result_addr : 9'sh0 ) ;
	assign w_sub14_result_datain = ( (|r_sys_processing_methodID) ? r_sub14_result_datain : 32'h0 ) ;
	assign w_sub14_result_r_w = ( (|r_sys_processing_methodID) ? r_sub14_result_r_w : 1'h0 ) ;
	assign w_sub01_u_addr = ( (|r_sys_processing_methodID) ? r_sub01_u_addr : 9'sh0 ) ;
	assign w_sub01_u_datain = ( (|r_sys_processing_methodID) ? r_sub01_u_datain : 32'h0 ) ;
	assign w_sub01_u_r_w = ( (|r_sys_processing_methodID) ? r_sub01_u_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 9'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub00_u_addr = ( (|r_sys_processing_methodID) ? r_sub00_u_addr : 9'sh0 ) ;
	assign w_sub00_u_datain = ( (|r_sys_processing_methodID) ? r_sub00_u_datain : 32'h0 ) ;
	assign w_sub00_u_r_w = ( (|r_sys_processing_methodID) ? r_sub00_u_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 9'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sub13_u_addr = ( (|r_sys_processing_methodID) ? r_sub13_u_addr : 9'sh0 ) ;
	assign w_sub13_u_datain = ( (|r_sys_processing_methodID) ? r_sub13_u_datain : 32'h0 ) ;
	assign w_sub13_u_r_w = ( (|r_sys_processing_methodID) ? r_sub13_u_r_w : 1'h0 ) ;
	assign w_sub13_result_addr = ( (|r_sys_processing_methodID) ? r_sub13_result_addr : 9'sh0 ) ;
	assign w_sub13_result_datain = ( (|r_sys_processing_methodID) ? r_sub13_result_datain : 32'h0 ) ;
	assign w_sub13_result_r_w = ( (|r_sys_processing_methodID) ? r_sub13_result_r_w : 1'h0 ) ;
	assign w_sub07_u_addr = ( (|r_sys_processing_methodID) ? r_sub07_u_addr : 9'sh0 ) ;
	assign w_sub07_u_datain = ( (|r_sys_processing_methodID) ? r_sub07_u_datain : 32'h0 ) ;
	assign w_sub07_u_r_w = ( (|r_sys_processing_methodID) ? r_sub07_u_r_w : 1'h0 ) ;
	assign w_sub07_result_addr = ( (|r_sys_processing_methodID) ? r_sub07_result_addr : 9'sh0 ) ;
	assign w_sub07_result_datain = ( (|r_sys_processing_methodID) ? r_sub07_result_datain : 32'h0 ) ;
	assign w_sub07_result_r_w = ( (|r_sys_processing_methodID) ? r_sub07_result_r_w : 1'h0 ) ;
	assign w_sub16_u_addr = ( (|r_sys_processing_methodID) ? r_sub16_u_addr : 9'sh0 ) ;
	assign w_sub16_u_datain = ( (|r_sys_processing_methodID) ? r_sub16_u_datain : 32'h0 ) ;
	assign w_sub16_u_r_w = ( (|r_sys_processing_methodID) ? r_sub16_u_r_w : 1'h0 ) ;
	assign w_sub16_result_addr = ( (|r_sys_processing_methodID) ? r_sub16_result_addr : 9'sh0 ) ;
	assign w_sub16_result_datain = ( (|r_sys_processing_methodID) ? r_sub16_result_datain : 32'h0 ) ;
	assign w_sub16_result_r_w = ( (|r_sys_processing_methodID) ? r_sub16_result_r_w : 1'h0 ) ;
	assign w_sub06_u_addr = ( (|r_sys_processing_methodID) ? r_sub06_u_addr : 9'sh0 ) ;
	assign w_sub06_u_datain = ( (|r_sys_processing_methodID) ? r_sub06_u_datain : 32'h0 ) ;
	assign w_sub06_u_r_w = ( (|r_sys_processing_methodID) ? r_sub06_u_r_w : 1'h0 ) ;
	assign w_sub06_result_addr = ( (|r_sys_processing_methodID) ? r_sub06_result_addr : 9'sh0 ) ;
	assign w_sub06_result_datain = ( (|r_sys_processing_methodID) ? r_sub06_result_datain : 32'h0 ) ;
	assign w_sub06_result_r_w = ( (|r_sys_processing_methodID) ? r_sub06_result_r_w : 1'h0 ) ;
	assign w_sub15_u_addr = ( (|r_sys_processing_methodID) ? r_sub15_u_addr : 9'sh0 ) ;
	assign w_sub15_u_datain = ( (|r_sys_processing_methodID) ? r_sub15_u_datain : 32'h0 ) ;
	assign w_sub15_u_r_w = ( (|r_sys_processing_methodID) ? r_sub15_u_r_w : 1'h0 ) ;
	assign w_sub15_result_addr = ( (|r_sys_processing_methodID) ? r_sub15_result_addr : 9'sh0 ) ;
	assign w_sub15_result_datain = ( (|r_sys_processing_methodID) ? r_sub15_result_datain : 32'h0 ) ;
	assign w_sub15_result_r_w = ( (|r_sys_processing_methodID) ? r_sub15_result_r_w : 1'h0 ) ;
	assign w_sub05_u_addr = ( (|r_sys_processing_methodID) ? r_sub05_u_addr : 9'sh0 ) ;
	assign w_sub05_u_datain = ( (|r_sys_processing_methodID) ? r_sub05_u_datain : 32'h0 ) ;
	assign w_sub05_u_r_w = ( (|r_sys_processing_methodID) ? r_sub05_u_r_w : 1'h0 ) ;
	assign w_sub05_q_addr = ( (|r_sys_processing_methodID) ? r_sub05_q_addr : 9'sh0 ) ;
	assign w_sub05_q_datain = ( (|r_sys_processing_methodID) ? r_sub05_q_datain : 32'h0 ) ;
	assign w_sub05_q_r_w = ( (|r_sys_processing_methodID) ? r_sub05_q_r_w : 1'h0 ) ;
	assign w_sub05_result_addr = ( (|r_sys_processing_methodID) ? r_sub05_result_addr : 9'sh0 ) ;
	assign w_sub05_result_datain = ( (|r_sys_processing_methodID) ? r_sub05_result_datain : 32'h0 ) ;
	assign w_sub05_result_r_w = ( (|r_sys_processing_methodID) ? r_sub05_result_r_w : 1'h0 ) ;
	assign w_sub18_u_addr = ( (|r_sys_processing_methodID) ? r_sub18_u_addr : 9'sh0 ) ;
	assign w_sub18_u_datain = ( (|r_sys_processing_methodID) ? r_sub18_u_datain : 32'h0 ) ;
	assign w_sub18_u_r_w = ( (|r_sys_processing_methodID) ? r_sub18_u_r_w : 1'h0 ) ;
	assign w_sub18_result_addr = ( (|r_sys_processing_methodID) ? r_sub18_result_addr : 9'sh0 ) ;
	assign w_sub18_result_datain = ( (|r_sys_processing_methodID) ? r_sub18_result_datain : 32'h0 ) ;
	assign w_sub18_result_r_w = ( (|r_sys_processing_methodID) ? r_sub18_result_r_w : 1'h0 ) ;
	assign w_sub04_u_addr = ( (|r_sys_processing_methodID) ? r_sub04_u_addr : 9'sh0 ) ;
	assign w_sub04_u_datain = ( (|r_sys_processing_methodID) ? r_sub04_u_datain : 32'h0 ) ;
	assign w_sub04_u_r_w = ( (|r_sys_processing_methodID) ? r_sub04_u_r_w : 1'h0 ) ;
	assign w_sub04_result_addr = ( (|r_sys_processing_methodID) ? r_sub04_result_addr : 9'sh0 ) ;
	assign w_sub04_result_datain = ( (|r_sys_processing_methodID) ? r_sub04_result_datain : 32'h0 ) ;
	assign w_sub04_result_r_w = ( (|r_sys_processing_methodID) ? r_sub04_result_r_w : 1'h0 ) ;
	assign w_sub17_u_addr = ( (|r_sys_processing_methodID) ? r_sub17_u_addr : 9'sh0 ) ;
	assign w_sub17_u_datain = ( (|r_sys_processing_methodID) ? r_sub17_u_datain : 32'h0 ) ;
	assign w_sub17_u_r_w = ( (|r_sys_processing_methodID) ? r_sub17_u_r_w : 1'h0 ) ;
	assign w_sub17_result_addr = ( (|r_sys_processing_methodID) ? r_sub17_result_addr : 9'sh0 ) ;
	assign w_sub17_result_datain = ( (|r_sys_processing_methodID) ? r_sub17_result_datain : 32'h0 ) ;
	assign w_sub17_result_r_w = ( (|r_sys_processing_methodID) ? r_sub17_result_r_w : 1'h0 ) ;
	assign w_sub10_u_addr = ( (|r_sys_processing_methodID) ? r_sub10_u_addr : 9'sh0 ) ;
	assign w_sub10_u_datain = ( (|r_sys_processing_methodID) ? r_sub10_u_datain : 32'h0 ) ;
	assign w_sub10_u_r_w = ( (|r_sys_processing_methodID) ? r_sub10_u_r_w : 1'h0 ) ;
	assign w_sub10_result_addr = ( (|r_sys_processing_methodID) ? r_sub10_result_addr : 9'sh0 ) ;
	assign w_sub10_result_datain = ( (|r_sys_processing_methodID) ? r_sub10_result_datain : 32'h0 ) ;
	assign w_sub10_result_r_w = ( (|r_sys_processing_methodID) ? r_sub10_result_r_w : 1'h0 ) ;
	assign w_sub20_u_addr = ( (|r_sys_processing_methodID) ? r_sub20_u_addr : 9'sh0 ) ;
	assign w_sub20_u_datain = ( (|r_sys_processing_methodID) ? r_sub20_u_datain : 32'h0 ) ;
	assign w_sub20_u_r_w = ( (|r_sys_processing_methodID) ? r_sub20_u_r_w : 1'h0 ) ;
	assign w_sub20_result_addr = ( (|r_sys_processing_methodID) ? r_sub20_result_addr : 9'sh0 ) ;
	assign w_sub20_result_datain = ( (|r_sys_processing_methodID) ? r_sub20_result_datain : 32'h0 ) ;
	assign w_sub20_result_r_w = ( (|r_sys_processing_methodID) ? r_sub20_result_r_w : 1'h0 ) ;
	assign w_sub21_u_addr = ( (|r_sys_processing_methodID) ? r_sub21_u_addr : 9'sh0 ) ;
	assign w_sub21_u_datain = ( (|r_sys_processing_methodID) ? r_sub21_u_datain : 32'h0 ) ;
	assign w_sub21_u_r_w = ( (|r_sys_processing_methodID) ? r_sub21_u_r_w : 1'h0 ) ;
	assign w_sub21_q_addr = ( (|r_sys_processing_methodID) ? r_sub21_q_addr : 9'sh0 ) ;
	assign w_sub21_q_datain = ( (|r_sys_processing_methodID) ? r_sub21_q_datain : 32'h0 ) ;
	assign w_sub21_q_r_w = ( (|r_sys_processing_methodID) ? r_sub21_q_r_w : 1'h0 ) ;
	assign w_sub21_result_addr = ( (|r_sys_processing_methodID) ? r_sub21_result_addr : 9'sh0 ) ;
	assign w_sub21_result_datain = ( (|r_sys_processing_methodID) ? r_sub21_result_datain : 32'h0 ) ;
	assign w_sub21_result_r_w = ( (|r_sys_processing_methodID) ? r_sub21_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh00000015;
	assign w_sys_tmp3 = 32'h3d4ccccd;
	assign w_sys_tmp5 = 32'sh00000002;
	assign w_sys_tmp6 = ( !w_sys_tmp7 );
	assign w_sys_tmp7 = (r_run_my_31 < r_run_k_27);
	assign w_sys_tmp8 = (r_run_k_27 + w_sys_intOne);
	assign w_sys_tmp9 = ( !w_sys_tmp10 );
	assign w_sys_tmp10 = (r_run_mx_30 < r_run_j_28);
	assign w_sys_tmp13 = (w_sys_tmp14 + r_run_k_27);
	assign w_sys_tmp14 = (r_run_j_28 * w_sys_tmp15);
	assign w_sys_tmp15 = 32'sh00000015;
	assign w_sys_tmp16 = 32'h0;
	assign w_sys_tmp18 = (w_sys_tmp19 + r_run_k_27);
	assign w_sys_tmp19 = (r_run_copy0_j_35 * w_sys_tmp15);
	assign w_sys_tmp22 = (r_run_copy0_j_35 + w_sys_intOne);
	assign w_sys_tmp23 = (r_run_j_28 + w_sys_intOne);
	assign w_sys_tmp96 = ( !w_sys_tmp97 );
	assign w_sys_tmp97 = (r_run_nlast_32 < r_run_n_29);
	assign w_sys_tmp98 = (r_run_n_29 + w_sys_intOne);
	assign w_sys_tmp99 = ( !w_sys_tmp100 );
	assign w_sys_tmp100 = (r_run_my_31 < r_run_j_28);
	assign w_sys_tmp103 = (w_sys_tmp104 + r_run_j_28);
	assign w_sys_tmp104 = 32'sh00000015;
	assign w_sys_tmp105 = 32'h3f000000;
	assign w_sys_tmp107 = (w_sys_tmp108 + r_run_copy2_j_38);
	assign w_sys_tmp108 = (r_run_mx_30 * w_sys_tmp104);
	assign w_sys_tmp110 = 32'h0;
	assign w_sys_tmp112 = (w_sys_tmp113 + w_sys_intOne);
	assign w_sys_tmp113 = (r_run_copy1_j_37 * w_sys_tmp104);
	assign w_sys_tmp115 = 32'h3f800000;
	assign w_sys_tmp117 = (w_sys_tmp118 + r_run_my_31);
	assign w_sys_tmp118 = (r_run_copy0_j_36 * w_sys_tmp104);
	assign w_sys_tmp121 = (r_run_copy0_j_36 + w_sys_intOne);
	assign w_sys_tmp122 = (r_run_copy1_j_37 + w_sys_intOne);
	assign w_sys_tmp123 = (r_run_copy2_j_38 + w_sys_intOne);
	assign w_sys_tmp124 = (r_run_j_28 + w_sys_intOne);
	assign w_sys_tmp263 = ( !w_sys_tmp264 );
	assign w_sys_tmp264 = (w_sys_tmp265 < r_run_k_27);
	assign w_sys_tmp265 = 32'sh00000005;
	assign w_sys_tmp268 = (w_sys_tmp269 + r_run_k_27);
	assign w_sys_tmp269 = 32'sh00000015;
	assign w_sys_tmp270 = w_fld_u_0_dataout_1;
	assign w_sys_tmp274 = (w_sys_tmp275 + r_run_k_27);
	assign w_sys_tmp275 = 32'sh0000002a;
	assign w_sys_tmp280 = (w_sys_tmp281 + r_run_k_27);
	assign w_sys_tmp281 = 32'sh0000003f;
	assign w_sys_tmp286 = (w_sys_tmp287 + r_run_k_27);
	assign w_sys_tmp287 = 32'sh00000054;
	assign w_sys_tmp292 = (w_sys_tmp293 + r_run_k_27);
	assign w_sys_tmp293 = 32'sh00000069;
	assign w_sys_tmp310 = (w_sys_tmp311 + r_run_k_27);
	assign w_sys_tmp311 = 32'sh0000007e;
	assign w_sys_tmp316 = (w_sys_tmp317 + r_run_k_27);
	assign w_sys_tmp317 = 32'sh00000093;
	assign w_sys_tmp322 = (w_sys_tmp323 + r_run_k_27);
	assign w_sys_tmp323 = 32'sh000000a8;
	assign w_sys_tmp328 = (w_sys_tmp329 + r_run_k_27);
	assign w_sys_tmp329 = 32'sh000000bd;
	assign w_sys_tmp346 = (w_sys_tmp347 + r_run_k_27);
	assign w_sys_tmp347 = 32'sh000000d2;
	assign w_sys_tmp352 = (w_sys_tmp353 + r_run_k_27);
	assign w_sys_tmp353 = 32'sh000000e7;
	assign w_sys_tmp358 = (w_sys_tmp359 + r_run_k_27);
	assign w_sys_tmp359 = 32'sh000000fc;
	assign w_sys_tmp364 = (w_sys_tmp365 + r_run_k_27);
	assign w_sys_tmp365 = 32'sh00000111;
	assign w_sys_tmp382 = (w_sys_tmp383 + r_run_k_27);
	assign w_sys_tmp383 = 32'sh00000126;
	assign w_sys_tmp388 = (w_sys_tmp389 + r_run_k_27);
	assign w_sys_tmp389 = 32'sh0000013b;
	assign w_sys_tmp394 = (w_sys_tmp395 + r_run_k_27);
	assign w_sys_tmp395 = 32'sh00000150;
	assign w_sys_tmp400 = (w_sys_tmp401 + r_run_k_27);
	assign w_sys_tmp401 = 32'sh00000165;
	assign w_sys_tmp418 = (w_sys_tmp419 + r_run_k_27);
	assign w_sys_tmp419 = 32'sh0000017a;
	assign w_sys_tmp424 = (w_sys_tmp425 + r_run_k_27);
	assign w_sys_tmp425 = 32'sh0000018f;
	assign w_sys_tmp430 = (w_sys_tmp431 + r_run_k_27);
	assign w_sys_tmp431 = 32'sh000001a4;
	assign w_sys_tmp436 = (w_sys_tmp437 + r_run_k_27);
	assign w_sys_tmp437 = 32'sh000001b9;
	assign w_sys_tmp441 = (r_run_k_27 + w_sys_intOne);
	assign w_sys_tmp442 = 32'sh00000004;
	assign w_sys_tmp443 = ( !w_sys_tmp444 );
	assign w_sys_tmp444 = (w_sys_tmp445 < r_run_k_27);
	assign w_sys_tmp445 = 32'sh00000009;
	assign w_sys_tmp448 = (w_sys_tmp449 + r_run_k_27);
	assign w_sys_tmp449 = 32'sh00000015;
	assign w_sys_tmp450 = w_fld_u_0_dataout_1;
	assign w_sys_tmp454 = (w_sys_tmp455 + r_run_k_27);
	assign w_sys_tmp455 = 32'sh0000002a;
	assign w_sys_tmp460 = (w_sys_tmp461 + r_run_k_27);
	assign w_sys_tmp461 = 32'sh0000003f;
	assign w_sys_tmp466 = (w_sys_tmp467 + r_run_k_27);
	assign w_sys_tmp467 = 32'sh00000054;
	assign w_sys_tmp472 = (w_sys_tmp473 + r_run_k_27);
	assign w_sys_tmp473 = 32'sh00000069;
	assign w_sys_tmp490 = (w_sys_tmp491 + r_run_k_27);
	assign w_sys_tmp491 = 32'sh0000007e;
	assign w_sys_tmp496 = (w_sys_tmp497 + r_run_k_27);
	assign w_sys_tmp497 = 32'sh00000093;
	assign w_sys_tmp502 = (w_sys_tmp503 + r_run_k_27);
	assign w_sys_tmp503 = 32'sh000000a8;
	assign w_sys_tmp508 = (w_sys_tmp509 + r_run_k_27);
	assign w_sys_tmp509 = 32'sh000000bd;
	assign w_sys_tmp526 = (w_sys_tmp527 + r_run_k_27);
	assign w_sys_tmp527 = 32'sh000000d2;
	assign w_sys_tmp532 = (w_sys_tmp533 + r_run_k_27);
	assign w_sys_tmp533 = 32'sh000000e7;
	assign w_sys_tmp538 = (w_sys_tmp539 + r_run_k_27);
	assign w_sys_tmp539 = 32'sh000000fc;
	assign w_sys_tmp544 = (w_sys_tmp545 + r_run_k_27);
	assign w_sys_tmp545 = 32'sh00000111;
	assign w_sys_tmp562 = (w_sys_tmp563 + r_run_k_27);
	assign w_sys_tmp563 = 32'sh00000126;
	assign w_sys_tmp568 = (w_sys_tmp569 + r_run_k_27);
	assign w_sys_tmp569 = 32'sh0000013b;
	assign w_sys_tmp574 = (w_sys_tmp575 + r_run_k_27);
	assign w_sys_tmp575 = 32'sh00000150;
	assign w_sys_tmp580 = (w_sys_tmp581 + r_run_k_27);
	assign w_sys_tmp581 = 32'sh00000165;
	assign w_sys_tmp598 = (w_sys_tmp599 + r_run_k_27);
	assign w_sys_tmp599 = 32'sh0000017a;
	assign w_sys_tmp604 = (w_sys_tmp605 + r_run_k_27);
	assign w_sys_tmp605 = 32'sh0000018f;
	assign w_sys_tmp610 = (w_sys_tmp611 + r_run_k_27);
	assign w_sys_tmp611 = 32'sh000001a4;
	assign w_sys_tmp616 = (w_sys_tmp617 + r_run_k_27);
	assign w_sys_tmp617 = 32'sh000001b9;
	assign w_sys_tmp622 = (w_sys_tmp623 + r_run_k_27);
	assign w_sys_tmp623 = 32'sh00000019;
	assign w_sys_tmp628 = (w_sys_tmp629 + r_run_k_27);
	assign w_sys_tmp629 = 32'sh0000002e;
	assign w_sys_tmp634 = (w_sys_tmp635 + r_run_k_27);
	assign w_sys_tmp635 = 32'sh00000043;
	assign w_sys_tmp640 = (w_sys_tmp641 + r_run_k_27);
	assign w_sys_tmp641 = 32'sh00000058;
	assign w_sys_tmp646 = (w_sys_tmp647 + r_run_k_27);
	assign w_sys_tmp647 = 32'sh0000006d;
	assign w_sys_tmp664 = (w_sys_tmp665 + r_run_k_27);
	assign w_sys_tmp665 = 32'sh00000082;
	assign w_sys_tmp670 = (w_sys_tmp671 + r_run_k_27);
	assign w_sys_tmp671 = 32'sh00000097;
	assign w_sys_tmp676 = (w_sys_tmp677 + r_run_k_27);
	assign w_sys_tmp677 = 32'sh000000ac;
	assign w_sys_tmp682 = (w_sys_tmp683 + r_run_k_27);
	assign w_sys_tmp683 = 32'sh000000c1;
	assign w_sys_tmp700 = (w_sys_tmp701 + r_run_k_27);
	assign w_sys_tmp701 = 32'sh000000d6;
	assign w_sys_tmp706 = (w_sys_tmp707 + r_run_k_27);
	assign w_sys_tmp707 = 32'sh000000eb;
	assign w_sys_tmp712 = (w_sys_tmp713 + r_run_k_27);
	assign w_sys_tmp713 = 32'sh00000100;
	assign w_sys_tmp718 = (w_sys_tmp719 + r_run_k_27);
	assign w_sys_tmp719 = 32'sh00000115;
	assign w_sys_tmp736 = (w_sys_tmp737 + r_run_k_27);
	assign w_sys_tmp737 = 32'sh0000012a;
	assign w_sys_tmp742 = (w_sys_tmp743 + r_run_k_27);
	assign w_sys_tmp743 = 32'sh0000013f;
	assign w_sys_tmp748 = (w_sys_tmp749 + r_run_k_27);
	assign w_sys_tmp749 = 32'sh00000154;
	assign w_sys_tmp754 = (w_sys_tmp755 + r_run_k_27);
	assign w_sys_tmp755 = 32'sh00000169;
	assign w_sys_tmp772 = (w_sys_tmp773 + r_run_k_27);
	assign w_sys_tmp773 = 32'sh0000017e;
	assign w_sys_tmp778 = (w_sys_tmp779 + r_run_k_27);
	assign w_sys_tmp779 = 32'sh00000193;
	assign w_sys_tmp784 = (w_sys_tmp785 + r_run_k_27);
	assign w_sys_tmp785 = 32'sh000001a8;
	assign w_sys_tmp790 = (w_sys_tmp791 + r_run_k_27);
	assign w_sys_tmp791 = 32'sh000001bd;
	assign w_sys_tmp796 = (w_sys_tmp797 + r_run_k_27);
	assign w_sys_tmp797 = 32'sh0000001d;
	assign w_sys_tmp802 = (w_sys_tmp803 + r_run_k_27);
	assign w_sys_tmp803 = 32'sh00000032;
	assign w_sys_tmp808 = (w_sys_tmp809 + r_run_k_27);
	assign w_sys_tmp809 = 32'sh00000047;
	assign w_sys_tmp814 = (w_sys_tmp815 + r_run_k_27);
	assign w_sys_tmp815 = 32'sh0000005c;
	assign w_sys_tmp820 = (w_sys_tmp821 + r_run_k_27);
	assign w_sys_tmp821 = 32'sh00000071;
	assign w_sys_tmp838 = (w_sys_tmp839 + r_run_k_27);
	assign w_sys_tmp839 = 32'sh00000086;
	assign w_sys_tmp844 = (w_sys_tmp845 + r_run_k_27);
	assign w_sys_tmp845 = 32'sh0000009b;
	assign w_sys_tmp850 = (w_sys_tmp851 + r_run_k_27);
	assign w_sys_tmp851 = 32'sh000000b0;
	assign w_sys_tmp856 = (w_sys_tmp857 + r_run_k_27);
	assign w_sys_tmp857 = 32'sh000000c5;
	assign w_sys_tmp874 = (w_sys_tmp875 + r_run_k_27);
	assign w_sys_tmp875 = 32'sh000000da;
	assign w_sys_tmp880 = (w_sys_tmp881 + r_run_k_27);
	assign w_sys_tmp881 = 32'sh000000ef;
	assign w_sys_tmp886 = (w_sys_tmp887 + r_run_k_27);
	assign w_sys_tmp887 = 32'sh00000104;
	assign w_sys_tmp892 = (w_sys_tmp893 + r_run_k_27);
	assign w_sys_tmp893 = 32'sh00000119;
	assign w_sys_tmp910 = (w_sys_tmp911 + r_run_k_27);
	assign w_sys_tmp911 = 32'sh0000012e;
	assign w_sys_tmp916 = (w_sys_tmp917 + r_run_k_27);
	assign w_sys_tmp917 = 32'sh00000143;
	assign w_sys_tmp922 = (w_sys_tmp923 + r_run_k_27);
	assign w_sys_tmp923 = 32'sh00000158;
	assign w_sys_tmp928 = (w_sys_tmp929 + r_run_k_27);
	assign w_sys_tmp929 = 32'sh0000016d;
	assign w_sys_tmp946 = (w_sys_tmp947 + r_run_k_27);
	assign w_sys_tmp947 = 32'sh00000182;
	assign w_sys_tmp952 = (w_sys_tmp953 + r_run_k_27);
	assign w_sys_tmp953 = 32'sh00000197;
	assign w_sys_tmp958 = (w_sys_tmp959 + r_run_k_27);
	assign w_sys_tmp959 = 32'sh000001ac;
	assign w_sys_tmp964 = (w_sys_tmp965 + r_run_k_27);
	assign w_sys_tmp965 = 32'sh000001c1;
	assign w_sys_tmp970 = (w_sys_tmp971 + r_run_k_27);
	assign w_sys_tmp971 = 32'sh00000021;
	assign w_sys_tmp976 = (w_sys_tmp977 + r_run_k_27);
	assign w_sys_tmp977 = 32'sh00000036;
	assign w_sys_tmp982 = (w_sys_tmp983 + r_run_k_27);
	assign w_sys_tmp983 = 32'sh0000004b;
	assign w_sys_tmp988 = (w_sys_tmp989 + r_run_k_27);
	assign w_sys_tmp989 = 32'sh00000060;
	assign w_sys_tmp994 = (w_sys_tmp995 + r_run_k_27);
	assign w_sys_tmp995 = 32'sh00000075;
	assign w_sys_tmp1012 = (w_sys_tmp1013 + r_run_k_27);
	assign w_sys_tmp1013 = 32'sh0000008a;
	assign w_sys_tmp1018 = (w_sys_tmp1019 + r_run_k_27);
	assign w_sys_tmp1019 = 32'sh0000009f;
	assign w_sys_tmp1024 = (w_sys_tmp1025 + r_run_k_27);
	assign w_sys_tmp1025 = 32'sh000000b4;
	assign w_sys_tmp1030 = (w_sys_tmp1031 + r_run_k_27);
	assign w_sys_tmp1031 = 32'sh000000c9;
	assign w_sys_tmp1048 = (w_sys_tmp1049 + r_run_k_27);
	assign w_sys_tmp1049 = 32'sh000000de;
	assign w_sys_tmp1054 = (w_sys_tmp1055 + r_run_k_27);
	assign w_sys_tmp1055 = 32'sh000000f3;
	assign w_sys_tmp1060 = (w_sys_tmp1061 + r_run_k_27);
	assign w_sys_tmp1061 = 32'sh00000108;
	assign w_sys_tmp1066 = (w_sys_tmp1067 + r_run_k_27);
	assign w_sys_tmp1067 = 32'sh0000011d;
	assign w_sys_tmp1084 = (w_sys_tmp1085 + r_run_k_27);
	assign w_sys_tmp1085 = 32'sh00000132;
	assign w_sys_tmp1090 = (w_sys_tmp1091 + r_run_k_27);
	assign w_sys_tmp1091 = 32'sh00000147;
	assign w_sys_tmp1096 = (w_sys_tmp1097 + r_run_k_27);
	assign w_sys_tmp1097 = 32'sh0000015c;
	assign w_sys_tmp1102 = (w_sys_tmp1103 + r_run_k_27);
	assign w_sys_tmp1103 = 32'sh00000171;
	assign w_sys_tmp1120 = (w_sys_tmp1121 + r_run_k_27);
	assign w_sys_tmp1121 = 32'sh00000186;
	assign w_sys_tmp1126 = (w_sys_tmp1127 + r_run_k_27);
	assign w_sys_tmp1127 = 32'sh0000019b;
	assign w_sys_tmp1132 = (w_sys_tmp1133 + r_run_k_27);
	assign w_sys_tmp1133 = 32'sh000001b0;
	assign w_sys_tmp1138 = (w_sys_tmp1139 + r_run_k_27);
	assign w_sys_tmp1139 = 32'sh000001c5;
	assign w_sys_tmp1143 = (r_run_k_27 + w_sys_intOne);
	assign w_sys_tmp1144 = 32'sh00000002;
	assign w_sys_tmp1145 = ( !w_sys_tmp1146 );
	assign w_sys_tmp1146 = (w_sys_tmp1147 < r_run_k_27);
	assign w_sys_tmp1147 = 32'sh00000004;
	assign w_sys_tmp1150 = (w_sys_tmp1151 + r_run_k_27);
	assign w_sys_tmp1151 = 32'sh0000002a;
	assign w_sys_tmp1152 = w_sub00_result_dataout;
	assign w_sys_tmp1156 = (w_sys_tmp1157 + r_run_k_27);
	assign w_sys_tmp1157 = 32'sh0000003f;
	assign w_sys_tmp1162 = (w_sys_tmp1163 + r_run_k_27);
	assign w_sys_tmp1163 = 32'sh00000054;
	assign w_sys_tmp1168 = (w_sys_tmp1169 + r_run_k_27);
	assign w_sys_tmp1169 = 32'sh00000069;
	assign w_sys_tmp1173 = (w_sys_tmp1174 + r_run_k_27);
	assign w_sys_tmp1174 = 32'sh0000007e;
	assign w_sys_tmp1178 = (w_sys_tmp1179 + r_run_k_27);
	assign w_sys_tmp1179 = 32'sh00000093;
	assign w_sys_tmp1183 = (w_sys_tmp1184 + r_run_k_27);
	assign w_sys_tmp1184 = 32'sh000000a8;
	assign w_sys_tmp1188 = (w_sys_tmp1189 + r_run_k_27);
	assign w_sys_tmp1189 = 32'sh000000bd;
	assign w_sys_tmp1193 = (w_sys_tmp1194 + r_run_k_27);
	assign w_sys_tmp1194 = 32'sh000000d2;
	assign w_sys_tmp1198 = (w_sys_tmp1199 + r_run_k_27);
	assign w_sys_tmp1199 = 32'sh000000e7;
	assign w_sys_tmp1203 = (w_sys_tmp1204 + r_run_k_27);
	assign w_sys_tmp1204 = 32'sh000000fc;
	assign w_sys_tmp1208 = (w_sys_tmp1209 + r_run_k_27);
	assign w_sys_tmp1209 = 32'sh00000111;
	assign w_sys_tmp1213 = (w_sys_tmp1214 + r_run_k_27);
	assign w_sys_tmp1214 = 32'sh00000126;
	assign w_sys_tmp1218 = (w_sys_tmp1219 + r_run_k_27);
	assign w_sys_tmp1219 = 32'sh0000013b;
	assign w_sys_tmp1223 = (w_sys_tmp1224 + r_run_k_27);
	assign w_sys_tmp1224 = 32'sh00000150;
	assign w_sys_tmp1228 = (w_sys_tmp1229 + r_run_k_27);
	assign w_sys_tmp1229 = 32'sh00000165;
	assign w_sys_tmp1233 = (w_sys_tmp1234 + r_run_k_27);
	assign w_sys_tmp1234 = 32'sh0000017a;
	assign w_sys_tmp1238 = (w_sys_tmp1239 + r_run_k_27);
	assign w_sys_tmp1239 = 32'sh0000018f;
	assign w_sys_tmp1243 = (w_sys_tmp1244 + r_run_k_27);
	assign w_sys_tmp1244 = 32'sh000001a4;
	assign w_sys_tmp1247 = (r_run_k_27 + w_sys_intOne);
	assign w_sys_tmp1248 = 32'sh00000005;
	assign w_sys_tmp1249 = ( !w_sys_tmp1250 );
	assign w_sys_tmp1250 = (w_sys_tmp1251 < r_run_k_27);
	assign w_sys_tmp1251 = 32'sh00000008;
	assign w_sys_tmp1254 = (w_sys_tmp1255 + r_run_k_27);
	assign w_sys_tmp1255 = 32'sh0000002a;
	assign w_sys_tmp1256 = w_sub05_result_dataout;
	assign w_sys_tmp1260 = (w_sys_tmp1261 + r_run_k_27);
	assign w_sys_tmp1261 = 32'sh0000003f;
	assign w_sys_tmp1266 = (w_sys_tmp1267 + r_run_k_27);
	assign w_sys_tmp1267 = 32'sh00000054;
	assign w_sys_tmp1272 = (w_sys_tmp1273 + r_run_k_27);
	assign w_sys_tmp1273 = 32'sh00000069;
	assign w_sys_tmp1277 = (w_sys_tmp1278 + r_run_k_27);
	assign w_sys_tmp1278 = 32'sh0000007e;
	assign w_sys_tmp1282 = (w_sys_tmp1283 + r_run_k_27);
	assign w_sys_tmp1283 = 32'sh00000093;
	assign w_sys_tmp1287 = (w_sys_tmp1288 + r_run_k_27);
	assign w_sys_tmp1288 = 32'sh000000a8;
	assign w_sys_tmp1292 = (w_sys_tmp1293 + r_run_k_27);
	assign w_sys_tmp1293 = 32'sh000000bd;
	assign w_sys_tmp1297 = (w_sys_tmp1298 + r_run_k_27);
	assign w_sys_tmp1298 = 32'sh000000d2;
	assign w_sys_tmp1302 = (w_sys_tmp1303 + r_run_k_27);
	assign w_sys_tmp1303 = 32'sh000000e7;
	assign w_sys_tmp1307 = (w_sys_tmp1308 + r_run_k_27);
	assign w_sys_tmp1308 = 32'sh000000fc;
	assign w_sys_tmp1312 = (w_sys_tmp1313 + r_run_k_27);
	assign w_sys_tmp1313 = 32'sh00000111;
	assign w_sys_tmp1317 = (w_sys_tmp1318 + r_run_k_27);
	assign w_sys_tmp1318 = 32'sh00000126;
	assign w_sys_tmp1322 = (w_sys_tmp1323 + r_run_k_27);
	assign w_sys_tmp1323 = 32'sh0000013b;
	assign w_sys_tmp1327 = (w_sys_tmp1328 + r_run_k_27);
	assign w_sys_tmp1328 = 32'sh00000150;
	assign w_sys_tmp1332 = (w_sys_tmp1333 + r_run_k_27);
	assign w_sys_tmp1333 = 32'sh00000165;
	assign w_sys_tmp1337 = (w_sys_tmp1338 + r_run_k_27);
	assign w_sys_tmp1338 = 32'sh0000017a;
	assign w_sys_tmp1342 = (w_sys_tmp1343 + r_run_k_27);
	assign w_sys_tmp1343 = 32'sh0000018f;
	assign w_sys_tmp1347 = (w_sys_tmp1348 + r_run_k_27);
	assign w_sys_tmp1348 = 32'sh000001a4;
	assign w_sys_tmp1351 = (r_run_k_27 + w_sys_intOne);
	assign w_sys_tmp1352 = 32'sh00000009;
	assign w_sys_tmp1353 = ( !w_sys_tmp1354 );
	assign w_sys_tmp1354 = (w_sys_tmp1355 < r_run_k_27);
	assign w_sys_tmp1355 = 32'sh0000000c;
	assign w_sys_tmp1358 = (w_sys_tmp1359 + r_run_k_27);
	assign w_sys_tmp1359 = 32'sh0000002e;
	assign w_sys_tmp1360 = w_sub10_result_dataout;
	assign w_sys_tmp1364 = (w_sys_tmp1365 + r_run_k_27);
	assign w_sys_tmp1365 = 32'sh00000043;
	assign w_sys_tmp1370 = (w_sys_tmp1371 + r_run_k_27);
	assign w_sys_tmp1371 = 32'sh00000058;
	assign w_sys_tmp1376 = (w_sys_tmp1377 + r_run_k_27);
	assign w_sys_tmp1377 = 32'sh0000006d;
	assign w_sys_tmp1381 = (w_sys_tmp1382 + r_run_k_27);
	assign w_sys_tmp1382 = 32'sh00000082;
	assign w_sys_tmp1386 = (w_sys_tmp1387 + r_run_k_27);
	assign w_sys_tmp1387 = 32'sh00000097;
	assign w_sys_tmp1391 = (w_sys_tmp1392 + r_run_k_27);
	assign w_sys_tmp1392 = 32'sh000000ac;
	assign w_sys_tmp1396 = (w_sys_tmp1397 + r_run_k_27);
	assign w_sys_tmp1397 = 32'sh000000c1;
	assign w_sys_tmp1401 = (w_sys_tmp1402 + r_run_k_27);
	assign w_sys_tmp1402 = 32'sh000000d6;
	assign w_sys_tmp1406 = (w_sys_tmp1407 + r_run_k_27);
	assign w_sys_tmp1407 = 32'sh000000eb;
	assign w_sys_tmp1411 = (w_sys_tmp1412 + r_run_k_27);
	assign w_sys_tmp1412 = 32'sh00000100;
	assign w_sys_tmp1416 = (w_sys_tmp1417 + r_run_k_27);
	assign w_sys_tmp1417 = 32'sh00000115;
	assign w_sys_tmp1421 = (w_sys_tmp1422 + r_run_k_27);
	assign w_sys_tmp1422 = 32'sh0000012a;
	assign w_sys_tmp1426 = (w_sys_tmp1427 + r_run_k_27);
	assign w_sys_tmp1427 = 32'sh0000013f;
	assign w_sys_tmp1431 = (w_sys_tmp1432 + r_run_k_27);
	assign w_sys_tmp1432 = 32'sh00000154;
	assign w_sys_tmp1436 = (w_sys_tmp1437 + r_run_k_27);
	assign w_sys_tmp1437 = 32'sh00000169;
	assign w_sys_tmp1441 = (w_sys_tmp1442 + r_run_k_27);
	assign w_sys_tmp1442 = 32'sh0000017e;
	assign w_sys_tmp1446 = (w_sys_tmp1447 + r_run_k_27);
	assign w_sys_tmp1447 = 32'sh00000193;
	assign w_sys_tmp1451 = (w_sys_tmp1452 + r_run_k_27);
	assign w_sys_tmp1452 = 32'sh000001a8;
	assign w_sys_tmp1456 = (w_sys_tmp1457 + r_run_k_27);
	assign w_sys_tmp1457 = 32'sh00000032;
	assign w_sys_tmp1461 = (w_sys_tmp1462 + r_run_k_27);
	assign w_sys_tmp1462 = 32'sh00000047;
	assign w_sys_tmp1466 = (w_sys_tmp1467 + r_run_k_27);
	assign w_sys_tmp1467 = 32'sh0000005c;
	assign w_sys_tmp1471 = (w_sys_tmp1472 + r_run_k_27);
	assign w_sys_tmp1472 = 32'sh00000071;
	assign w_sys_tmp1476 = (w_sys_tmp1477 + r_run_k_27);
	assign w_sys_tmp1477 = 32'sh00000086;
	assign w_sys_tmp1481 = (w_sys_tmp1482 + r_run_k_27);
	assign w_sys_tmp1482 = 32'sh0000009b;
	assign w_sys_tmp1486 = (w_sys_tmp1487 + r_run_k_27);
	assign w_sys_tmp1487 = 32'sh000000b0;
	assign w_sys_tmp1491 = (w_sys_tmp1492 + r_run_k_27);
	assign w_sys_tmp1492 = 32'sh000000c5;
	assign w_sys_tmp1496 = (w_sys_tmp1497 + r_run_k_27);
	assign w_sys_tmp1497 = 32'sh000000da;
	assign w_sys_tmp1501 = (w_sys_tmp1502 + r_run_k_27);
	assign w_sys_tmp1502 = 32'sh000000ef;
	assign w_sys_tmp1506 = (w_sys_tmp1507 + r_run_k_27);
	assign w_sys_tmp1507 = 32'sh00000104;
	assign w_sys_tmp1511 = (w_sys_tmp1512 + r_run_k_27);
	assign w_sys_tmp1512 = 32'sh00000119;
	assign w_sys_tmp1516 = (w_sys_tmp1517 + r_run_k_27);
	assign w_sys_tmp1517 = 32'sh0000012e;
	assign w_sys_tmp1521 = (w_sys_tmp1522 + r_run_k_27);
	assign w_sys_tmp1522 = 32'sh00000143;
	assign w_sys_tmp1526 = (w_sys_tmp1527 + r_run_k_27);
	assign w_sys_tmp1527 = 32'sh00000158;
	assign w_sys_tmp1531 = (w_sys_tmp1532 + r_run_k_27);
	assign w_sys_tmp1532 = 32'sh0000016d;
	assign w_sys_tmp1536 = (w_sys_tmp1537 + r_run_k_27);
	assign w_sys_tmp1537 = 32'sh00000182;
	assign w_sys_tmp1541 = (w_sys_tmp1542 + r_run_k_27);
	assign w_sys_tmp1542 = 32'sh00000197;
	assign w_sys_tmp1546 = (w_sys_tmp1547 + r_run_k_27);
	assign w_sys_tmp1547 = 32'sh000001ac;
	assign w_sys_tmp1551 = (w_sys_tmp1552 + r_run_k_27);
	assign w_sys_tmp1552 = 32'sh00000036;
	assign w_sys_tmp1556 = (w_sys_tmp1557 + r_run_k_27);
	assign w_sys_tmp1557 = 32'sh0000004b;
	assign w_sys_tmp1561 = (w_sys_tmp1562 + r_run_k_27);
	assign w_sys_tmp1562 = 32'sh00000060;
	assign w_sys_tmp1566 = (w_sys_tmp1567 + r_run_k_27);
	assign w_sys_tmp1567 = 32'sh00000075;
	assign w_sys_tmp1571 = (w_sys_tmp1572 + r_run_k_27);
	assign w_sys_tmp1572 = 32'sh0000008a;
	assign w_sys_tmp1576 = (w_sys_tmp1577 + r_run_k_27);
	assign w_sys_tmp1577 = 32'sh0000009f;
	assign w_sys_tmp1581 = (w_sys_tmp1582 + r_run_k_27);
	assign w_sys_tmp1582 = 32'sh000000b4;
	assign w_sys_tmp1586 = (w_sys_tmp1587 + r_run_k_27);
	assign w_sys_tmp1587 = 32'sh000000c9;
	assign w_sys_tmp1591 = (w_sys_tmp1592 + r_run_k_27);
	assign w_sys_tmp1592 = 32'sh000000de;
	assign w_sys_tmp1596 = (w_sys_tmp1597 + r_run_k_27);
	assign w_sys_tmp1597 = 32'sh000000f3;
	assign w_sys_tmp1601 = (w_sys_tmp1602 + r_run_k_27);
	assign w_sys_tmp1602 = 32'sh00000108;
	assign w_sys_tmp1606 = (w_sys_tmp1607 + r_run_k_27);
	assign w_sys_tmp1607 = 32'sh0000011d;
	assign w_sys_tmp1611 = (w_sys_tmp1612 + r_run_k_27);
	assign w_sys_tmp1612 = 32'sh00000132;
	assign w_sys_tmp1616 = (w_sys_tmp1617 + r_run_k_27);
	assign w_sys_tmp1617 = 32'sh00000147;
	assign w_sys_tmp1621 = (w_sys_tmp1622 + r_run_k_27);
	assign w_sys_tmp1622 = 32'sh0000015c;
	assign w_sys_tmp1626 = (w_sys_tmp1627 + r_run_k_27);
	assign w_sys_tmp1627 = 32'sh00000171;
	assign w_sys_tmp1631 = (w_sys_tmp1632 + r_run_k_27);
	assign w_sys_tmp1632 = 32'sh00000186;
	assign w_sys_tmp1636 = (w_sys_tmp1637 + r_run_k_27);
	assign w_sys_tmp1637 = 32'sh0000019b;
	assign w_sys_tmp1641 = (w_sys_tmp1642 + r_run_k_27);
	assign w_sys_tmp1642 = 32'sh000001b0;
	assign w_sys_tmp1645 = (r_run_k_27 + w_sys_intOne);


	sub19
		sub19_inst(
			.i_fld_result_1_addr_0 (w_sub19_result_addr),
			.i_fld_result_1_datain_0 (w_sub19_result_datain),
			.o_fld_result_1_dataout_0 (w_sub19_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub19_result_r_w),
			.i_fld_u_0_addr_0 (w_sub19_u_addr),
			.i_fld_u_0_datain_0 (w_sub19_u_datain),
			.o_fld_u_0_dataout_0 (w_sub19_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub19_u_r_w),
			.o_run_busy (w_sub19_run_busy),
			.i_run_req (r_sub19_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub09
		sub09_inst(
			.i_fld_result_1_addr_0 (w_sub09_result_addr),
			.i_fld_result_1_datain_0 (w_sub09_result_datain),
			.o_fld_result_1_dataout_0 (w_sub09_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub09_result_r_w),
			.i_fld_u_0_addr_0 (w_sub09_u_addr),
			.i_fld_u_0_datain_0 (w_sub09_u_datain),
			.o_fld_u_0_dataout_0 (w_sub09_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub09_u_r_w),
			.o_run_busy (w_sub09_run_busy),
			.i_run_req (r_sub09_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub08
		sub08_inst(
			.i_fld_result_1_addr_0 (w_sub08_result_addr),
			.i_fld_result_1_datain_0 (w_sub08_result_datain),
			.o_fld_result_1_dataout_0 (w_sub08_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub08_result_r_w),
			.i_fld_u_0_addr_0 (w_sub08_u_addr),
			.i_fld_u_0_datain_0 (w_sub08_u_datain),
			.o_fld_u_0_dataout_0 (w_sub08_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub08_u_r_w),
			.o_run_busy (w_sub08_run_busy),
			.i_run_req (r_sub08_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub24
		sub24_inst(
			.i_fld_result_1_addr_0 (w_sub24_result_addr),
			.i_fld_result_1_datain_0 (w_sub24_result_datain),
			.o_fld_result_1_dataout_0 (w_sub24_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub24_result_r_w),
			.i_fld_u_0_addr_0 (w_sub24_u_addr),
			.i_fld_u_0_datain_0 (w_sub24_u_datain),
			.o_fld_u_0_dataout_0 (w_sub24_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub24_u_r_w),
			.o_run_busy (w_sub24_run_busy),
			.i_run_req (r_sub24_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub22
		sub22_inst(
			.i_fld_result_1_addr_0 (w_sub22_result_addr),
			.i_fld_result_1_datain_0 (w_sub22_result_datain),
			.o_fld_result_1_dataout_0 (w_sub22_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub22_result_r_w),
			.i_fld_u_0_addr_0 (w_sub22_u_addr),
			.i_fld_u_0_datain_0 (w_sub22_u_datain),
			.o_fld_u_0_dataout_0 (w_sub22_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub22_u_r_w),
			.o_run_busy (w_sub22_run_busy),
			.i_run_req (r_sub22_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub23
		sub23_inst(
			.i_fld_result_1_addr_0 (w_sub23_result_addr),
			.i_fld_result_1_datain_0 (w_sub23_result_datain),
			.o_fld_result_1_dataout_0 (w_sub23_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub23_result_r_w),
			.i_fld_u_0_addr_0 (w_sub23_u_addr),
			.i_fld_u_0_datain_0 (w_sub23_u_datain),
			.o_fld_u_0_dataout_0 (w_sub23_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub23_u_r_w),
			.o_run_busy (w_sub23_run_busy),
			.i_run_req (r_sub23_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub12
		sub12_inst(
			.i_fld_result_1_addr_0 (w_sub12_result_addr),
			.i_fld_result_1_datain_0 (w_sub12_result_datain),
			.o_fld_result_1_dataout_0 (w_sub12_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub12_result_r_w),
			.i_fld_u_0_addr_0 (w_sub12_u_addr),
			.i_fld_u_0_datain_0 (w_sub12_u_datain),
			.o_fld_u_0_dataout_0 (w_sub12_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub12_u_r_w),
			.o_run_busy (w_sub12_run_busy),
			.i_run_req (r_sub12_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub03
		sub03_inst(
			.i_fld_result_1_addr_0 (w_sub03_result_addr),
			.i_fld_result_1_datain_0 (w_sub03_result_datain),
			.o_fld_result_1_dataout_0 (w_sub03_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub03_result_r_w),
			.i_fld_u_0_addr_0 (w_sub03_u_addr),
			.i_fld_u_0_datain_0 (w_sub03_u_datain),
			.o_fld_u_0_dataout_0 (w_sub03_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub03_u_r_w),
			.o_run_busy (w_sub03_run_busy),
			.i_run_req (r_sub03_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub02
		sub02_inst(
			.i_fld_result_1_addr_0 (w_sub02_result_addr),
			.i_fld_result_1_datain_0 (w_sub02_result_datain),
			.o_fld_result_1_dataout_0 (w_sub02_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub02_result_r_w),
			.i_fld_u_0_addr_0 (w_sub02_u_addr),
			.i_fld_u_0_datain_0 (w_sub02_u_datain),
			.o_fld_u_0_dataout_0 (w_sub02_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub02_u_r_w),
			.o_run_busy (w_sub02_run_busy),
			.i_run_req (r_sub02_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub11
		sub11_inst(
			.i_fld_result_1_addr_0 (w_sub11_result_addr),
			.i_fld_result_1_datain_0 (w_sub11_result_datain),
			.o_fld_result_1_dataout_0 (w_sub11_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub11_result_r_w),
			.i_fld_u_0_addr_0 (w_sub11_u_addr),
			.i_fld_u_0_datain_0 (w_sub11_u_datain),
			.o_fld_u_0_dataout_0 (w_sub11_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub11_u_r_w),
			.o_run_busy (w_sub11_run_busy),
			.i_run_req (r_sub11_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub14
		sub14_inst(
			.i_fld_result_1_addr_0 (w_sub14_result_addr),
			.i_fld_result_1_datain_0 (w_sub14_result_datain),
			.o_fld_result_1_dataout_0 (w_sub14_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub14_result_r_w),
			.i_fld_u_0_addr_0 (w_sub14_u_addr),
			.i_fld_u_0_datain_0 (w_sub14_u_datain),
			.o_fld_u_0_dataout_0 (w_sub14_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub14_u_r_w),
			.o_run_busy (w_sub14_run_busy),
			.i_run_req (r_sub14_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub01
		sub01_inst(
			.i_fld_result_1_addr_0 (w_sub01_result_addr),
			.i_fld_result_1_datain_0 (w_sub01_result_datain),
			.o_fld_result_1_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub01_result_r_w),
			.i_fld_u_0_addr_0 (w_sub01_u_addr),
			.i_fld_u_0_datain_0 (w_sub01_u_datain),
			.o_fld_u_0_dataout_0 (w_sub01_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub01_u_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub00
		sub00_inst(
			.i_fld_result_1_addr_0 (w_sub00_result_addr),
			.i_fld_result_1_datain_0 (w_sub00_result_datain),
			.o_fld_result_1_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub00_result_r_w),
			.i_fld_u_0_addr_0 (w_sub00_u_addr),
			.i_fld_u_0_datain_0 (w_sub00_u_datain),
			.o_fld_u_0_dataout_0 (w_sub00_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub00_u_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub13
		sub13_inst(
			.i_fld_result_1_addr_0 (w_sub13_result_addr),
			.i_fld_result_1_datain_0 (w_sub13_result_datain),
			.o_fld_result_1_dataout_0 (w_sub13_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub13_result_r_w),
			.i_fld_u_0_addr_0 (w_sub13_u_addr),
			.i_fld_u_0_datain_0 (w_sub13_u_datain),
			.o_fld_u_0_dataout_0 (w_sub13_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub13_u_r_w),
			.o_run_busy (w_sub13_run_busy),
			.i_run_req (r_sub13_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub07
		sub07_inst(
			.i_fld_result_1_addr_0 (w_sub07_result_addr),
			.i_fld_result_1_datain_0 (w_sub07_result_datain),
			.o_fld_result_1_dataout_0 (w_sub07_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub07_result_r_w),
			.i_fld_u_0_addr_0 (w_sub07_u_addr),
			.i_fld_u_0_datain_0 (w_sub07_u_datain),
			.o_fld_u_0_dataout_0 (w_sub07_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub07_u_r_w),
			.o_run_busy (w_sub07_run_busy),
			.i_run_req (r_sub07_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub16
		sub16_inst(
			.i_fld_result_1_addr_0 (w_sub16_result_addr),
			.i_fld_result_1_datain_0 (w_sub16_result_datain),
			.o_fld_result_1_dataout_0 (w_sub16_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub16_result_r_w),
			.i_fld_u_0_addr_0 (w_sub16_u_addr),
			.i_fld_u_0_datain_0 (w_sub16_u_datain),
			.o_fld_u_0_dataout_0 (w_sub16_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub16_u_r_w),
			.o_run_busy (w_sub16_run_busy),
			.i_run_req (r_sub16_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub06
		sub06_inst(
			.i_fld_result_1_addr_0 (w_sub06_result_addr),
			.i_fld_result_1_datain_0 (w_sub06_result_datain),
			.o_fld_result_1_dataout_0 (w_sub06_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub06_result_r_w),
			.i_fld_u_0_addr_0 (w_sub06_u_addr),
			.i_fld_u_0_datain_0 (w_sub06_u_datain),
			.o_fld_u_0_dataout_0 (w_sub06_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub06_u_r_w),
			.o_run_busy (w_sub06_run_busy),
			.i_run_req (r_sub06_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub15
		sub15_inst(
			.i_fld_result_1_addr_0 (w_sub15_result_addr),
			.i_fld_result_1_datain_0 (w_sub15_result_datain),
			.o_fld_result_1_dataout_0 (w_sub15_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub15_result_r_w),
			.i_fld_u_0_addr_0 (w_sub15_u_addr),
			.i_fld_u_0_datain_0 (w_sub15_u_datain),
			.o_fld_u_0_dataout_0 (w_sub15_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub15_u_r_w),
			.o_run_busy (w_sub15_run_busy),
			.i_run_req (r_sub15_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub05
		sub05_inst(
			.i_fld_q_1_addr_0 (w_sub05_q_addr),
			.i_fld_q_1_datain_0 (w_sub05_q_datain),
			.o_fld_q_1_dataout_0 (w_sub05_q_dataout),
			.i_fld_q_1_r_w_0 (w_sub05_q_r_w),
			.i_fld_result_2_addr_0 (w_sub05_result_addr),
			.i_fld_result_2_datain_0 (w_sub05_result_datain),
			.o_fld_result_2_dataout_0 (w_sub05_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub05_result_r_w),
			.i_fld_u_0_addr_0 (w_sub05_u_addr),
			.i_fld_u_0_datain_0 (w_sub05_u_datain),
			.o_fld_u_0_dataout_0 (w_sub05_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub05_u_r_w),
			.o_run_busy (w_sub05_run_busy),
			.i_run_req (r_sub05_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub18
		sub18_inst(
			.i_fld_result_1_addr_0 (w_sub18_result_addr),
			.i_fld_result_1_datain_0 (w_sub18_result_datain),
			.o_fld_result_1_dataout_0 (w_sub18_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub18_result_r_w),
			.i_fld_u_0_addr_0 (w_sub18_u_addr),
			.i_fld_u_0_datain_0 (w_sub18_u_datain),
			.o_fld_u_0_dataout_0 (w_sub18_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub18_u_r_w),
			.o_run_busy (w_sub18_run_busy),
			.i_run_req (r_sub18_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub04
		sub04_inst(
			.i_fld_result_1_addr_0 (w_sub04_result_addr),
			.i_fld_result_1_datain_0 (w_sub04_result_datain),
			.o_fld_result_1_dataout_0 (w_sub04_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub04_result_r_w),
			.i_fld_u_0_addr_0 (w_sub04_u_addr),
			.i_fld_u_0_datain_0 (w_sub04_u_datain),
			.o_fld_u_0_dataout_0 (w_sub04_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub04_u_r_w),
			.o_run_busy (w_sub04_run_busy),
			.i_run_req (r_sub04_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub17
		sub17_inst(
			.i_fld_result_1_addr_0 (w_sub17_result_addr),
			.i_fld_result_1_datain_0 (w_sub17_result_datain),
			.o_fld_result_1_dataout_0 (w_sub17_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub17_result_r_w),
			.i_fld_u_0_addr_0 (w_sub17_u_addr),
			.i_fld_u_0_datain_0 (w_sub17_u_datain),
			.o_fld_u_0_dataout_0 (w_sub17_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub17_u_r_w),
			.o_run_busy (w_sub17_run_busy),
			.i_run_req (r_sub17_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub10
		sub10_inst(
			.i_fld_result_1_addr_0 (w_sub10_result_addr),
			.i_fld_result_1_datain_0 (w_sub10_result_datain),
			.o_fld_result_1_dataout_0 (w_sub10_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub10_result_r_w),
			.i_fld_u_0_addr_0 (w_sub10_u_addr),
			.i_fld_u_0_datain_0 (w_sub10_u_datain),
			.o_fld_u_0_dataout_0 (w_sub10_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub10_u_r_w),
			.o_run_busy (w_sub10_run_busy),
			.i_run_req (r_sub10_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub20
		sub20_inst(
			.i_fld_result_1_addr_0 (w_sub20_result_addr),
			.i_fld_result_1_datain_0 (w_sub20_result_datain),
			.o_fld_result_1_dataout_0 (w_sub20_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub20_result_r_w),
			.i_fld_u_0_addr_0 (w_sub20_u_addr),
			.i_fld_u_0_datain_0 (w_sub20_u_datain),
			.o_fld_u_0_dataout_0 (w_sub20_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub20_u_r_w),
			.o_run_busy (w_sub20_run_busy),
			.i_run_req (r_sub20_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub21
		sub21_inst(
			.i_fld_q_1_addr_0 (w_sub21_q_addr),
			.i_fld_q_1_datain_0 (w_sub21_q_datain),
			.o_fld_q_1_dataout_0 (w_sub21_q_dataout),
			.i_fld_q_1_r_w_0 (w_sub21_q_r_w),
			.i_fld_result_2_addr_0 (w_sub21_result_addr),
			.i_fld_result_2_datain_0 (w_sub21_result_datain),
			.o_fld_result_2_dataout_0 (w_sub21_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub21_result_r_w),
			.i_fld_u_0_addr_0 (w_sub21_u_addr),
			.i_fld_u_0_datain_0 (w_sub21_u_datain),
			.o_fld_u_0_dataout_0 (w_sub21_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub21_u_r_w),
			.o_run_busy (w_sub21_run_busy),
			.i_run_req (r_sub21_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(9), .WORDS(484) )
		dpram_u_0(
			.clk (clock),
			.ce_0 (w_fld_u_0_ce_0),
			.addr_0 (w_fld_u_0_addr_0),
			.datain_0 (w_fld_u_0_datain_0),
			.dataout_0 (w_fld_u_0_dataout_0),
			.r_w_0 (w_fld_u_0_r_w_0),
			.ce_1 (w_fld_u_0_ce_1),
			.addr_1 (r_fld_u_0_addr_1),
			.datain_1 (r_fld_u_0_datain_1),
			.dataout_1 (w_fld_u_0_dataout_1),
			.r_w_1 (r_fld_u_0_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(9), .WORDS(484) )
		dpram_uu_1(
			.clk (clock),
			.ce_0 (w_fld_uu_1_ce_0),
			.addr_0 (w_fld_uu_1_addr_0),
			.datain_0 (w_fld_uu_1_datain_0),
			.dataout_0 (w_fld_uu_1_dataout_0),
			.r_w_0 (w_fld_uu_1_r_w_0),
			.ce_1 (w_fld_uu_1_ce_1),
			.addr_1 (r_fld_uu_1_addr_1),
			.datain_1 (r_fld_uu_1_datain_1),
			.dataout_1 (w_fld_uu_1_dataout_1),
			.r_w_1 (r_fld_uu_1_r_w_1)
		);

	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h3b: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 6'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_phase <= 6'h2;
						end

						6'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h4;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6) ? 6'h9 : 6'hf);

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'ha;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp9) ? 6'hd : 6'h6);

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_run_phase <= 6'ha;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h10;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp96) ? 6'h14 : 6'h3b);

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h10;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h15;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp99) ? 6'h18 : 6'h1a);

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1b)) begin
										r_sys_run_phase <= 6'h15;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h1b;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp263) ? 6'h1e : 6'h20);

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1e)) begin
										r_sys_run_phase <= 6'h1b;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h21;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp443) ? 6'h24 : 6'h25);

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h75)) begin
										r_sys_run_phase <= 6'h21;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h18: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_phase <= 6'h27;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h18: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_phase <= 6'h29;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h2a;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1145) ? 6'h2d : 6'h2f);

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h14)) begin
										r_sys_run_phase <= 6'h2a;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h30;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1249) ? 6'h33 : 6'h35);

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h14)) begin
										r_sys_run_phase <= 6'h30;

									end
								end

							endcase
						end

						6'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h36;

									end
								end

							endcase
						end

						6'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1353) ? 6'h39 : 6'h11);

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3a)) begin
										r_sys_run_phase <= 6'h36;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sys_run_phase <= 6'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 5'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1b)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1e)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h75)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h14)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h14)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3a)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 7'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h5)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1b)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h1a)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1e)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h1d)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h75)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h74)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h14)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h14)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3a)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h39)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						6'h3b: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_addr_1 <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp13[8:0] );

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp117[8:0] );

									end
									else
									if((r_sys_run_step==7'h1) || (r_sys_run_step==7'h5) || (r_sys_run_step==7'h9) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp107[8:0] );

									end
									else
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp112[8:0] );

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h4) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp103[8:0] );

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp280[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp274[8:0] );

									end
									else
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp286[8:0] );

									end
									else
									if((r_sys_run_step==7'h10) || (r_sys_run_step==7'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp364[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp424[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp310[8:0] );

									end
									else
									if((r_sys_run_step==7'h15) || (r_sys_run_step==7'h17)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp394[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp316[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp388[8:0] );

									end
									else
									if((r_sys_run_step==7'h16) || (r_sys_run_step==7'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp400[8:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp346[8:0] );

									end
									else
									if((r_sys_run_step==7'hf) || (r_sys_run_step==7'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp358[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp382[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp352[8:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp436[8:0] );

									end
									else
									if((r_sys_run_step==7'h4) || (r_sys_run_step==7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp292[8:0] );

									end
									else
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp322[8:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp418[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp268[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp430[8:0] );

									end
									else
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp328[8:0] );

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h61) || (r_sys_run_step==7'h63)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1030[8:0] );

									end
									else
									if((r_sys_run_step==7'h50) || (r_sys_run_step==7'h52)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp928[8:0] );

									end
									else
									if((r_sys_run_step==7'h16) || (r_sys_run_step==7'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp580[8:0] );

									end
									else
									if((r_sys_run_step==7'h3d) || (r_sys_run_step==7'h3f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp814[8:0] );

									end
									else
									if((r_sys_run_step==7'h55)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp958[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp448[8:0] );

									end
									else
									if((r_sys_run_step==7'h6d) || (r_sys_run_step==7'h6f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1102[8:0] );

									end
									else
									if((r_sys_run_step==7'h48)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp880[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp454[8:0] );

									end
									else
									if((r_sys_run_step==7'h66) || (r_sys_run_step==7'h68)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1060[8:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp616[8:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp598[8:0] );

									end
									else
									if((r_sys_run_step==7'h71)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1126[8:0] );

									end
									else
									if((r_sys_run_step==7'h65)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1054[8:0] );

									end
									else
									if((r_sys_run_step==7'h4d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp910[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp568[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp610[8:0] );

									end
									else
									if((r_sys_run_step==7'h70)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1120[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp604[8:0] );

									end
									else
									if((r_sys_run_step==7'h4) || (r_sys_run_step==7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp472[8:0] );

									end
									else
									if((r_sys_run_step==7'h39)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp790[8:0] );

									end
									else
									if((r_sys_run_step==7'h73)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1138[8:0] );

									end
									else
									if((r_sys_run_step==7'h2b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp706[8:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp634[8:0] );

									end
									else
									if((r_sys_run_step==7'h37)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp778[8:0] );

									end
									else
									if((r_sys_run_step==7'h24)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp664[8:0] );

									end
									else
									if((r_sys_run_step==7'hf) || (r_sys_run_step==7'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp538[8:0] );

									end
									else
									if((r_sys_run_step==7'h26) || (r_sys_run_step==7'h28)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp676[8:0] );

									end
									else
									if((r_sys_run_step==7'h49) || (r_sys_run_step==7'h4b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp886[8:0] );

									end
									else
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp466[8:0] );

									end
									else
									if((r_sys_run_step==7'h57)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp970[8:0] );

									end
									else
									if((r_sys_run_step==7'h3b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp802[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp496[8:0] );

									end
									else
									if((r_sys_run_step==7'h6c) || (r_sys_run_step==7'h6e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1096[8:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp622[8:0] );

									end
									else
									if((r_sys_run_step==7'h58)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp976[8:0] );

									end
									else
									if((r_sys_run_step==7'h27) || (r_sys_run_step==7'h29)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp682[8:0] );

									end
									else
									if((r_sys_run_step==7'h56)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp964[8:0] );

									end
									else
									if((r_sys_run_step==7'h3a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp796[8:0] );

									end
									else
									if((r_sys_run_step==7'h6a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1084[8:0] );

									end
									else
									if((r_sys_run_step==7'h53)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp946[8:0] );

									end
									else
									if((r_sys_run_step==7'h3c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp808[8:0] );

									end
									else
									if((r_sys_run_step==7'h36)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp772[8:0] );

									end
									else
									if((r_sys_run_step==7'h60) || (r_sys_run_step==7'h62)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1024[8:0] );

									end
									else
									if((r_sys_run_step==7'h4a) || (r_sys_run_step==7'h4c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp892[8:0] );

									end
									else
									if((r_sys_run_step==7'h15) || (r_sys_run_step==7'h17)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp574[8:0] );

									end
									else
									if((r_sys_run_step==7'h42)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp844[8:0] );

									end
									else
									if((r_sys_run_step==7'h10) || (r_sys_run_step==7'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp544[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp490[8:0] );

									end
									else
									if((r_sys_run_step==7'h31)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp742[8:0] );

									end
									else
									if((r_sys_run_step==7'h20) || (r_sys_run_step==7'h22)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp640[8:0] );

									end
									else
									if((r_sys_run_step==7'h2a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp700[8:0] );

									end
									else
									if((r_sys_run_step==7'h4e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp916[8:0] );

									end
									else
									if((r_sys_run_step==7'h43) || (r_sys_run_step==7'h45)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp850[8:0] );

									end
									else
									if((r_sys_run_step==7'h21) || (r_sys_run_step==7'h23)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp646[8:0] );

									end
									else
									if((r_sys_run_step==7'h2d) || (r_sys_run_step==7'h2f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp718[8:0] );

									end
									else
									if((r_sys_run_step==7'h32) || (r_sys_run_step==7'h34)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp748[8:0] );

									end
									else
									if((r_sys_run_step==7'h44) || (r_sys_run_step==7'h46)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp856[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp460[8:0] );

									end
									else
									if((r_sys_run_step==7'h33) || (r_sys_run_step==7'h35)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp754[8:0] );

									end
									else
									if((r_sys_run_step==7'h6b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1090[8:0] );

									end
									else
									if((r_sys_run_step==7'h72)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1132[8:0] );

									end
									else
									if((r_sys_run_step==7'h30)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp736[8:0] );

									end
									else
									if((r_sys_run_step==7'h38)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp784[8:0] );

									end
									else
									if((r_sys_run_step==7'h54)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp952[8:0] );

									end
									else
									if((r_sys_run_step==7'h25)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp670[8:0] );

									end
									else
									if((r_sys_run_step==7'h3e) || (r_sys_run_step==7'h40)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp820[8:0] );

									end
									else
									if((r_sys_run_step==7'h5a) || (r_sys_run_step==7'h5c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp988[8:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp628[8:0] );

									end
									else
									if((r_sys_run_step==7'h41)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp838[8:0] );

									end
									else
									if((r_sys_run_step==7'h47)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp874[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp562[8:0] );

									end
									else
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp502[8:0] );

									end
									else
									if((r_sys_run_step==7'h4f) || (r_sys_run_step==7'h51)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp922[8:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp526[8:0] );

									end
									else
									if((r_sys_run_step==7'h5e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1012[8:0] );

									end
									else
									if((r_sys_run_step==7'h5b) || (r_sys_run_step==7'h5d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp994[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp532[8:0] );

									end
									else
									if((r_sys_run_step==7'h59)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp982[8:0] );

									end
									else
									if((r_sys_run_step==7'h2c) || (r_sys_run_step==7'h2e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp712[8:0] );

									end
									else
									if((r_sys_run_step==7'h64)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1048[8:0] );

									end
									else
									if((r_sys_run_step==7'h67) || (r_sys_run_step==7'h69)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1066[8:0] );

									end
									else
									if((r_sys_run_step==7'h5f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1018[8:0] );

									end
									else
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp508[8:0] );

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1218[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1168[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1228[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1223[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1178[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1173[8:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1198[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1183[8:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1193[8:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1208[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1243[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1238[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1233[8:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1203[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1188[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1213[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1150[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1156[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1162[8:0] );

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1312[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1277[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1317[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1254[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1347[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1327[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1337[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1322[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1282[8:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1302[8:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1307[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1292[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1342[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1272[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1287[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1260[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1266[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1332[8:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1297[8:0] );

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1376[8:0] );

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1516[8:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1411[8:0] );

									end
									else
									if((r_sys_run_step==7'h3a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1641[8:0] );

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1461[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1358[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1396[8:0] );

									end
									else
									if((r_sys_run_step==7'h27)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1546[8:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1496[8:0] );

									end
									else
									if((r_sys_run_step==7'h28)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1551[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1451[8:0] );

									end
									else
									if((r_sys_run_step==7'h39)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1636[8:0] );

									end
									else
									if((r_sys_run_step==7'h32)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1601[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1364[8:0] );

									end
									else
									if((r_sys_run_step==7'h2c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1571[8:0] );

									end
									else
									if((r_sys_run_step==7'h2b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1566[8:0] );

									end
									else
									if((r_sys_run_step==7'h22)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1521[8:0] );

									end
									else
									if((r_sys_run_step==7'h31)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1596[8:0] );

									end
									else
									if((r_sys_run_step==7'h30)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1591[8:0] );

									end
									else
									if((r_sys_run_step==7'h38)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1631[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1436[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1381[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1481[8:0] );

									end
									else
									if((r_sys_run_step==7'h34)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1611[8:0] );

									end
									else
									if((r_sys_run_step==7'h23)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1526[8:0] );

									end
									else
									if((r_sys_run_step==7'h25)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1536[8:0] );

									end
									else
									if((r_sys_run_step==7'h37)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1626[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1426[8:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1471[8:0] );

									end
									else
									if((r_sys_run_step==7'h2f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1586[8:0] );

									end
									else
									if((r_sys_run_step==7'h2d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1576[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1441[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1431[8:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1406[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1370[8:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1501[8:0] );

									end
									else
									if((r_sys_run_step==7'h2a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1561[8:0] );

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1466[8:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1456[8:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1506[8:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1511[8:0] );

									end
									else
									if((r_sys_run_step==7'h29)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1556[8:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1401[8:0] );

									end
									else
									if((r_sys_run_step==7'h26)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1541[8:0] );

									end
									else
									if((r_sys_run_step==7'h24)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1531[8:0] );

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1616[8:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1416[8:0] );

									end
									else
									if((r_sys_run_step==7'h2e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1581[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1421[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1446[8:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1491[8:0] );

									end
									else
									if((r_sys_run_step==7'h36)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1621[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1391[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1386[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1486[8:0] );

									end
									else
									if((r_sys_run_step==7'h33)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1606[8:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1476[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp16;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h4) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h18)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp105;

									end
									else
									if((r_sys_run_step==7'h1) || (r_sys_run_step==7'h3) || (r_sys_run_step==7'h5) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'h9) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h1b)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp110;

									end
									else
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1a)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp115;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h3) || (r_sys_run_step==7'h4)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp1152;

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h8)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp14_float;

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp11_float;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h12)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h3) || (r_sys_run_step==7'h4)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp1256;

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h8)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp14_float;

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp11_float;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp21_float;

									end
									else
									if((r_sys_run_step==7'h24)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp44_float;

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h8)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp52_float;

									end
									else
									if((r_sys_run_step==7'h37)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp40_float;

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp48_float;

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp22_float;

									end
									else
									if((r_sys_run_step==7'h23)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==7'h2f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp42_float;

									end
									else
									if((r_sys_run_step==7'h39)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp14_float;

									end
									else
									if((r_sys_run_step==7'h22)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp19_float;

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==7'h29)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp31_float;

									end
									else
									if((r_sys_run_step==7'h33)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp41_float;

									end
									else
									if((r_sys_run_step==7'h25)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp32_float;

									end
									else
									if((r_sys_run_step==7'h2c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp30_float;

									end
									else
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h3) || (r_sys_run_step==7'h4)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp1360;

									end
									else
									if((r_sys_run_step==7'h2e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==7'h36)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==7'h2a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==7'h30)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp29_float;

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==7'h32)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==7'h27)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==7'h34)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp28_float;

									end
									else
									if((r_sys_run_step==7'h2d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp36_float;

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp25_float;

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp34_float;

									end
									else
									if((r_sys_run_step==7'h3a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp33_float;

									end
									else
									if((r_sys_run_step==7'h28)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp39_float;

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp26_float;

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp38_float;

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp37_float;

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp50_float;

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp51_float;

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp45_float;

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp23_float;

									end
									else
									if((r_sys_run_step==7'h38)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp27_float;

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp47_float;

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp46_float;

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp35_float;

									end
									else
									if((r_sys_run_step==7'h31)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp20_float;

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==7'h26)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp18_float;

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp24_float;

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp49_float;

									end
									else
									if((r_sys_run_step==7'h2b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp43_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h1b)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h1c)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h73)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h14)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h14)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h3a)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h3b: begin
							r_fld_u_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_uu_1_addr_1 <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_uu_1_addr_1 <= $signed( w_sys_tmp18[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_uu_1_datain_1 <= w_sys_tmp16;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_uu_1_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_uu_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h3b: begin
							r_fld_uu_1_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_27 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_27 <= w_sys_tmp8;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_27 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1e)) begin
										r_run_k_27 <= w_sys_tmp441;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_27 <= w_sys_tmp442;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h75)) begin
										r_run_k_27 <= w_sys_tmp1143;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_27 <= w_sys_tmp1144;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h14)) begin
										r_run_k_27 <= w_sys_tmp1247;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_27 <= w_sys_tmp1248;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h14)) begin
										r_run_k_27 <= w_sys_tmp1351;

									end
								end

							endcase
						end

						6'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_27 <= w_sys_tmp1352;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3a)) begin
										r_run_k_27 <= w_sys_tmp1645;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_28 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_28 <= w_sys_tmp23;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_28 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h4) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h18)) begin
										r_run_j_28 <= w_sys_tmp124;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_n_29 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_n_29 <= w_sys_tmp98;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_mx_30 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_my_31 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_nlast_32 <= w_sys_tmp5;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_dx_33 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_dy_34 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_35 <= r_run_j_28;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_35 <= w_sys_tmp22;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_36 <= r_run_j_28;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h1b)) begin
										r_run_copy0_j_36 <= w_sys_tmp121;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_37 <= r_run_j_28;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1a)) begin
										r_run_copy1_j_37 <= w_sys_tmp122;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy2_j_38 <= r_run_j_28;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1) || (r_sys_run_step==7'h5) || (r_sys_run_step==7'h9) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h19)) begin
										r_run_copy2_j_38 <= w_sys_tmp123;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub19_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub19_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h56)) begin
										r_sub19_u_addr <= $signed( w_sys_tmp952[8:0] );

									end
									else
									if((r_sys_run_step==7'h54)) begin
										r_sub19_u_addr <= $signed( w_sys_tmp928[8:0] );

									end
									else
									if((r_sys_run_step==7'h58)) begin
										r_sub19_u_addr <= $signed( w_sys_tmp964[8:0] );

									end
									else
									if((r_sys_run_step==7'h57)) begin
										r_sub19_u_addr <= $signed( w_sys_tmp958[8:0] );

									end
									else
									if((r_sys_run_step==7'h53)) begin
										r_sub19_u_addr <= $signed( w_sys_tmp922[8:0] );

									end
									else
									if((r_sys_run_step==7'h55)) begin
										r_sub19_u_addr <= $signed( w_sys_tmp946[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h53<=r_sys_run_step && r_sys_run_step<=7'h58)) begin
										r_sub19_u_datain <= w_sys_tmp450;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h53<=r_sys_run_step && r_sys_run_step<=7'h58)) begin
										r_sub19_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub19_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp1541[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp1536[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp1531[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp1546[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub19_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub09_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub09_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1e)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp616[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp598[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp580[8:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp574[8:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp610[8:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp604[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h19<=r_sys_run_step && r_sys_run_step<=7'h1e)) begin
										r_sub09_u_datain <= w_sys_tmp450;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h19<=r_sys_run_step && r_sys_run_step<=7'h1e)) begin
										r_sub09_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub09_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp1342[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp1347[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp1337[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp1332[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub09_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub08_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub08_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h18)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp580[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp538[8:0] );

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp574[8:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp562[8:0] );

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp568[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp544[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h13<=r_sys_run_step && r_sys_run_step<=7'h18)) begin
										r_sub08_u_datain <= w_sys_tmp450;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h13<=r_sys_run_step && r_sys_run_step<=7'h18)) begin
										r_sub08_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub08_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1312[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1317[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1327[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp1322[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub08_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub24_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub24_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h75)) begin
										r_sub24_u_addr <= $signed( w_sys_tmp1138[8:0] );

									end
									else
									if((r_sys_run_step==7'h70)) begin
										r_sub24_u_addr <= $signed( w_sys_tmp1096[8:0] );

									end
									else
									if((r_sys_run_step==7'h73)) begin
										r_sub24_u_addr <= $signed( w_sys_tmp1126[8:0] );

									end
									else
									if((r_sys_run_step==7'h72)) begin
										r_sub24_u_addr <= $signed( w_sys_tmp1120[8:0] );

									end
									else
									if((r_sys_run_step==7'h74)) begin
										r_sub24_u_addr <= $signed( w_sys_tmp1132[8:0] );

									end
									else
									if((r_sys_run_step==7'h71)) begin
										r_sub24_u_addr <= $signed( w_sys_tmp1102[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h70<=r_sys_run_step && r_sys_run_step<=7'h75)) begin
										r_sub24_u_datain <= w_sys_tmp450;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h70<=r_sys_run_step && r_sys_run_step<=7'h75)) begin
										r_sub24_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub24_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp1631[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp1636[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp1641[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp1626[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub24_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub22_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub22_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h68)) begin
										r_sub22_u_addr <= $signed( w_sys_tmp1060[8:0] );

									end
									else
									if((r_sys_run_step==7'h64)) begin
										r_sub22_u_addr <= $signed( w_sys_tmp1024[8:0] );

									end
									else
									if((r_sys_run_step==7'h65)) begin
										r_sub22_u_addr <= $signed( w_sys_tmp1030[8:0] );

									end
									else
									if((r_sys_run_step==7'h66)) begin
										r_sub22_u_addr <= $signed( w_sys_tmp1048[8:0] );

									end
									else
									if((r_sys_run_step==7'h67)) begin
										r_sub22_u_addr <= $signed( w_sys_tmp1054[8:0] );

									end
									else
									if((r_sys_run_step==7'h69)) begin
										r_sub22_u_addr <= $signed( w_sys_tmp1066[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h64<=r_sys_run_step && r_sys_run_step<=7'h69)) begin
										r_sub22_u_datain <= w_sys_tmp450;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h64<=r_sys_run_step && r_sys_run_step<=7'h69)) begin
										r_sub22_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub22_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp1586[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp1591[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp1601[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp1596[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub22_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub23_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub23_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6a)) begin
										r_sub23_u_addr <= $signed( w_sys_tmp1060[8:0] );

									end
									else
									if((r_sys_run_step==7'h6e)) begin
										r_sub23_u_addr <= $signed( w_sys_tmp1096[8:0] );

									end
									else
									if((r_sys_run_step==7'h6c)) begin
										r_sub23_u_addr <= $signed( w_sys_tmp1084[8:0] );

									end
									else
									if((r_sys_run_step==7'h6d)) begin
										r_sub23_u_addr <= $signed( w_sys_tmp1090[8:0] );

									end
									else
									if((r_sys_run_step==7'h6b)) begin
										r_sub23_u_addr <= $signed( w_sys_tmp1066[8:0] );

									end
									else
									if((r_sys_run_step==7'h6f)) begin
										r_sub23_u_addr <= $signed( w_sys_tmp1102[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h6a<=r_sys_run_step && r_sys_run_step<=7'h6f)) begin
										r_sub23_u_datain <= w_sys_tmp450;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h6a<=r_sys_run_step && r_sys_run_step<=7'h6f)) begin
										r_sub23_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub23_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp1611[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp1621[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp1616[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp1606[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub23_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub12_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub12_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2d)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp706[8:0] );

									end
									else
									if((r_sys_run_step==7'h2c)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp700[8:0] );

									end
									else
									if((r_sys_run_step==7'h2f)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp718[8:0] );

									end
									else
									if((r_sys_run_step==7'h2e)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp712[8:0] );

									end
									else
									if((r_sys_run_step==7'h2b)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp682[8:0] );

									end
									else
									if((r_sys_run_step==7'h2a)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp676[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2a<=r_sys_run_step && r_sys_run_step<=7'h2f)) begin
										r_sub12_u_datain <= w_sys_tmp450;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2a<=r_sys_run_step && r_sys_run_step<=7'h2f)) begin
										r_sub12_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub12_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp1401[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp1411[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp1406[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp1396[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub12_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h14)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp364[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp358[8:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp382[8:0] );

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp394[8:0] );

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp388[8:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp400[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h13<=r_sys_run_step && r_sys_run_step<=7'h18)) begin
										r_sub03_u_datain <= w_sys_tmp270;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h13<=r_sys_run_step && r_sys_run_step<=7'h18)) begin
										r_sub03_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub03_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1218[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1208[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1223[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1213[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub03_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hf)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp346[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp364[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp358[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp352[8:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp322[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp328[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'hd<=r_sys_run_step && r_sys_run_step<=7'h12)) begin
										r_sub02_u_datain <= w_sys_tmp270;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'hd<=r_sys_run_step && r_sys_run_step<=7'h12)) begin
										r_sub02_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub02_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1198[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1193[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1203[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1188[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub02_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub11_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub11_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h27)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp670[8:0] );

									end
									else
									if((r_sys_run_step==7'h24)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp640[8:0] );

									end
									else
									if((r_sys_run_step==7'h25)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp646[8:0] );

									end
									else
									if((r_sys_run_step==7'h26)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp664[8:0] );

									end
									else
									if((r_sys_run_step==7'h29)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp682[8:0] );

									end
									else
									if((r_sys_run_step==7'h28)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp676[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h24<=r_sys_run_step && r_sys_run_step<=7'h29)) begin
										r_sub11_u_datain <= w_sys_tmp450;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h24<=r_sys_run_step && r_sys_run_step<=7'h29)) begin
										r_sub11_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub11_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp1381[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp1376[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp1391[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp1386[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub11_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub14_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub14_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h39)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp778[8:0] );

									end
									else
									if((r_sys_run_step==7'h36)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp748[8:0] );

									end
									else
									if((r_sys_run_step==7'h37)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp754[8:0] );

									end
									else
									if((r_sys_run_step==7'h3b)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp790[8:0] );

									end
									else
									if((r_sys_run_step==7'h3a)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp784[8:0] );

									end
									else
									if((r_sys_run_step==7'h38)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp772[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h36<=r_sys_run_step && r_sys_run_step<=7'h3b)) begin
										r_sub14_u_datain <= w_sys_tmp450;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h36<=r_sys_run_step && r_sys_run_step<=7'h3b)) begin
										r_sub14_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub14_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp1446[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp1436[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp1451[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp1441[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub14_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp286[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp310[8:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp316[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp292[8:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp322[8:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp328[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h7<=r_sys_run_step && r_sys_run_step<=7'hc)) begin
										r_sub01_u_datain <= w_sys_tmp270;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h7<=r_sys_run_step && r_sys_run_step<=7'hc)) begin
										r_sub01_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub01_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1168[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1183[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1178[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1173[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp280[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp286[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp274[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp292[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp268[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub00_u_datain <= w_sys_tmp270;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub00_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub00_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1156[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1150[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1162[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h1) || (r_sys_run_step==7'h2)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub13_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub13_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h34)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp748[8:0] );

									end
									else
									if((r_sys_run_step==7'h31)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp718[8:0] );

									end
									else
									if((r_sys_run_step==7'h30)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp712[8:0] );

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp754[8:0] );

									end
									else
									if((r_sys_run_step==7'h32)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp736[8:0] );

									end
									else
									if((r_sys_run_step==7'h33)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp742[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h30<=r_sys_run_step && r_sys_run_step<=7'h35)) begin
										r_sub13_u_datain <= w_sys_tmp450;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h30<=r_sys_run_step && r_sys_run_step<=7'h35)) begin
										r_sub13_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub13_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp1421[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp1431[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp1426[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp1416[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub13_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub07_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub07_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h10)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp532[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp538[8:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp502[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp544[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp526[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp508[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'hd<=r_sys_run_step && r_sys_run_step<=7'h12)) begin
										r_sub07_u_datain <= w_sys_tmp450;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'hd<=r_sys_run_step && r_sys_run_step<=7'h12)) begin
										r_sub07_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub07_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1292[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1297[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1307[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp1302[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub07_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub16_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub16_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h42)) begin
										r_sub16_u_addr <= $signed( w_sys_tmp820[8:0] );

									end
									else
									if((r_sys_run_step==7'h45)) begin
										r_sub16_u_addr <= $signed( w_sys_tmp850[8:0] );

									end
									else
									if((r_sys_run_step==7'h43)) begin
										r_sub16_u_addr <= $signed( w_sys_tmp838[8:0] );

									end
									else
									if((r_sys_run_step==7'h46)) begin
										r_sub16_u_addr <= $signed( w_sys_tmp856[8:0] );

									end
									else
									if((r_sys_run_step==7'h41)) begin
										r_sub16_u_addr <= $signed( w_sys_tmp814[8:0] );

									end
									else
									if((r_sys_run_step==7'h44)) begin
										r_sub16_u_addr <= $signed( w_sys_tmp844[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h41<=r_sys_run_step && r_sys_run_step<=7'h46)) begin
										r_sub16_u_datain <= w_sys_tmp450;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h41<=r_sys_run_step && r_sys_run_step<=7'h46)) begin
										r_sub16_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub16_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp1471[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp1481[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp1486[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp1476[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub16_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub06_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub06_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp496[8:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp502[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp466[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp472[8:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp508[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp490[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h7<=r_sys_run_step && r_sys_run_step<=7'hc)) begin
										r_sub06_u_datain <= w_sys_tmp450;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h7<=r_sys_run_step && r_sys_run_step<=7'hc)) begin
										r_sub06_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub06_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1277[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1272[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1287[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp1282[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub06_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub15_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub15_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h40)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp820[8:0] );

									end
									else
									if((r_sys_run_step==7'h3f)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp814[8:0] );

									end
									else
									if((r_sys_run_step==7'h3c)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp796[8:0] );

									end
									else
									if((r_sys_run_step==7'h3d)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp802[8:0] );

									end
									else
									if((r_sys_run_step==7'h3e)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp808[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h3c<=r_sys_run_step && r_sys_run_step<=7'h40)) begin
										r_sub15_u_datain <= w_sys_tmp450;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h3c<=r_sys_run_step && r_sys_run_step<=7'h40)) begin
										r_sub15_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub15_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp1466[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp1456[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp1461[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h1) || (r_sys_run_step==7'h2)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub15_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub05_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub05_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp460[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp466[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp472[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp448[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp454[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub05_u_datain <= w_sys_tmp450;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub05_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub05_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_q_addr <= 9'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_q_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_q_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub05_q_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1254[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1266[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp1260[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h1) || (r_sys_run_step==7'h2)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub05_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub18_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub18_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h52)) begin
										r_sub18_u_addr <= $signed( w_sys_tmp928[8:0] );

									end
									else
									if((r_sys_run_step==7'h50)) begin
										r_sub18_u_addr <= $signed( w_sys_tmp916[8:0] );

									end
									else
									if((r_sys_run_step==7'h4e)) begin
										r_sub18_u_addr <= $signed( w_sys_tmp892[8:0] );

									end
									else
									if((r_sys_run_step==7'h4d)) begin
										r_sub18_u_addr <= $signed( w_sys_tmp886[8:0] );

									end
									else
									if((r_sys_run_step==7'h4f)) begin
										r_sub18_u_addr <= $signed( w_sys_tmp910[8:0] );

									end
									else
									if((r_sys_run_step==7'h51)) begin
										r_sub18_u_addr <= $signed( w_sys_tmp922[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h4d<=r_sys_run_step && r_sys_run_step<=7'h52)) begin
										r_sub18_u_datain <= w_sys_tmp450;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h4d<=r_sys_run_step && r_sys_run_step<=7'h52)) begin
										r_sub18_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub18_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp1511[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp1526[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp1516[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp1521[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub18_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub04_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub04_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1c)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp424[8:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp436[8:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp394[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp418[8:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp430[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp400[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h19<=r_sys_run_step && r_sys_run_step<=7'h1e)) begin
										r_sub04_u_datain <= w_sys_tmp270;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h19<=r_sys_run_step && r_sys_run_step<=7'h1e)) begin
										r_sub04_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub04_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1243[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1228[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1238[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1233[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub04_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub17_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub17_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4c)) begin
										r_sub17_u_addr <= $signed( w_sys_tmp892[8:0] );

									end
									else
									if((r_sys_run_step==7'h47)) begin
										r_sub17_u_addr <= $signed( w_sys_tmp850[8:0] );

									end
									else
									if((r_sys_run_step==7'h48)) begin
										r_sub17_u_addr <= $signed( w_sys_tmp856[8:0] );

									end
									else
									if((r_sys_run_step==7'h49)) begin
										r_sub17_u_addr <= $signed( w_sys_tmp874[8:0] );

									end
									else
									if((r_sys_run_step==7'h4b)) begin
										r_sub17_u_addr <= $signed( w_sys_tmp886[8:0] );

									end
									else
									if((r_sys_run_step==7'h4a)) begin
										r_sub17_u_addr <= $signed( w_sys_tmp880[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h47<=r_sys_run_step && r_sys_run_step<=7'h4c)) begin
										r_sub17_u_datain <= w_sys_tmp450;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h47<=r_sys_run_step && r_sys_run_step<=7'h4c)) begin
										r_sub17_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub17_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp1496[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp1506[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp1491[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp1501[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub17_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub10_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub10_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h22)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp640[8:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp628[8:0] );

									end
									else
									if((r_sys_run_step==7'h23)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp646[8:0] );

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp634[8:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp622[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h1f<=r_sys_run_step && r_sys_run_step<=7'h23)) begin
										r_sub10_u_datain <= w_sys_tmp450;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h1f<=r_sys_run_step && r_sys_run_step<=7'h23)) begin
										r_sub10_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub10_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp1364[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp1370[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp1358[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h1) || (r_sys_run_step==7'h2)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub10_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub20_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub20_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5c)) begin
										r_sub20_u_addr <= $signed( w_sys_tmp988[8:0] );

									end
									else
									if((r_sys_run_step==7'h5a)) begin
										r_sub20_u_addr <= $signed( w_sys_tmp976[8:0] );

									end
									else
									if((r_sys_run_step==7'h5b)) begin
										r_sub20_u_addr <= $signed( w_sys_tmp982[8:0] );

									end
									else
									if((r_sys_run_step==7'h59)) begin
										r_sub20_u_addr <= $signed( w_sys_tmp970[8:0] );

									end
									else
									if((r_sys_run_step==7'h5d)) begin
										r_sub20_u_addr <= $signed( w_sys_tmp994[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h59<=r_sys_run_step && r_sys_run_step<=7'h5d)) begin
										r_sub20_u_datain <= w_sys_tmp450;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h59<=r_sys_run_step && r_sys_run_step<=7'h5d)) begin
										r_sub20_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub20_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp1561[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp1551[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp1556[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h1) || (r_sys_run_step==7'h2)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub20_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub21_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub21_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h62)) begin
										r_sub21_u_addr <= $signed( w_sys_tmp1024[8:0] );

									end
									else
									if((r_sys_run_step==7'h5e)) begin
										r_sub21_u_addr <= $signed( w_sys_tmp988[8:0] );

									end
									else
									if((r_sys_run_step==7'h63)) begin
										r_sub21_u_addr <= $signed( w_sys_tmp1030[8:0] );

									end
									else
									if((r_sys_run_step==7'h61)) begin
										r_sub21_u_addr <= $signed( w_sys_tmp1018[8:0] );

									end
									else
									if((r_sys_run_step==7'h60)) begin
										r_sub21_u_addr <= $signed( w_sys_tmp1012[8:0] );

									end
									else
									if((r_sys_run_step==7'h5f)) begin
										r_sub21_u_addr <= $signed( w_sys_tmp994[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h5e<=r_sys_run_step && r_sys_run_step<=7'h63)) begin
										r_sub21_u_datain <= w_sys_tmp450;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h5e<=r_sys_run_step && r_sys_run_step<=7'h63)) begin
										r_sub21_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub21_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_q_addr <= 9'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_q_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_q_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub21_q_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp1576[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp1581[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp1571[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp1566[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h3b: begin
							r_sub21_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp0_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp0_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp0_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp1_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp1_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp1_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp2_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp2_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp2_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp3_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp3_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp3_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp4_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp4_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp4_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp5_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp5_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp5_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp6_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp6_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp6_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp7_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp7_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp7_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp8_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp8_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp8_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp9_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp9_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp9_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp10_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp10_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp10_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp11_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp11_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp11_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp12_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp12_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp12_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp13_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp13_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp13_float <= w_sub20_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h5)) begin
										r_sys_tmp14_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h5)) begin
										r_sys_tmp14_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp14_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp15_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp16_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp17_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp18_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp19_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp20_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp21_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp22_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp23_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp24_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp25_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp26_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp27_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp28_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp29_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp30_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp31_float <= w_sub20_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp32_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp33_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp34_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp35_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp36_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp37_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp38_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp39_float <= w_sub20_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp40_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp41_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp42_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp43_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp44_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp45_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp46_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp47_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp48_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp49_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp50_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp51_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h5)) begin
										r_sys_tmp52_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
