/*
TimeStamp:	2016/9/27		15:22
*/


module c1(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy	
);

	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 8:0] r_sys_run_phase;
	reg         [ 4:0] r_sys_run_stage;
	reg         [ 4:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 4:0] w_sys_run_stage_p1;
	wire        [ 4:0] w_sys_run_step_p1;
	wire signed [14:0] w_fld_u_0_addr_0;
	wire        [31:0] w_fld_u_0_datain_0;
	wire        [31:0] w_fld_u_0_dataout_0;
	wire               w_fld_u_0_r_w_0;
	wire               w_fld_u_0_ce_0;
	reg  signed [14:0] r_fld_u_0_addr_1;
	reg         [31:0] r_fld_u_0_datain_1;
	wire        [31:0] w_fld_u_0_dataout_1;
	reg                r_fld_u_0_r_w_1;
	wire               w_fld_u_0_ce_1;
	reg  signed [31:0] r_run_k_17;
	reg  signed [31:0] r_run_j_18;
	reg  signed [31:0] r_run_n_19;
	reg  signed [31:0] r_run_mx_20;
	reg  signed [31:0] r_run_my_21;
	reg  signed [31:0] r_run_nlast_22;
	reg  signed [31:0] r_run_copy0_j_23;
	reg  signed [31:0] r_run_copy1_j_24;
	reg  signed [31:0] r_run_copy2_j_25;
	reg  signed [31:0] r_run_copy0_j_26;
	reg  signed [31:0] r_run_copy0_j_27;
	reg  signed [31:0] r_run_copy0_j_28;
	reg  signed [31:0] r_run_copy0_j_29;
	reg  signed [31:0] r_run_copy0_j_30;
	reg  signed [31:0] r_run_copy0_j_31;
	reg  signed [31:0] r_run_copy0_j_32;
	reg  signed [31:0] r_run_copy0_j_33;
	reg  signed [31:0] r_run_copy0_j_34;
	reg  signed [31:0] r_run_copy0_j_35;
	reg  signed [31:0] r_run_copy0_j_36;
	reg  signed [31:0] r_run_copy0_j_37;
	reg  signed [31:0] r_run_copy0_j_38;
	reg  signed [31:0] r_run_copy0_j_39;
	reg  signed [31:0] r_run_copy0_j_40;
	reg  signed [31:0] r_run_copy0_j_41;
	reg  signed [31:0] r_run_copy0_j_42;
	reg  signed [31:0] r_run_copy0_j_43;
	reg  signed [31:0] r_run_copy0_j_44;
	reg  signed [31:0] r_run_copy0_j_45;
	reg  signed [31:0] r_run_copy0_j_46;
	reg  signed [31:0] r_run_copy0_j_47;
	reg  signed [31:0] r_run_copy0_j_48;
	reg  signed [31:0] r_run_copy0_j_49;
	reg  signed [31:0] r_run_copy0_j_50;
	reg  signed [31:0] r_run_copy0_j_51;
	reg  signed [31:0] r_run_copy0_j_52;
	reg  signed [31:0] r_run_copy0_j_53;
	reg  signed [31:0] r_run_copy0_j_54;
	reg  signed [31:0] r_run_copy0_j_55;
	reg  signed [31:0] r_run_copy0_j_56;
	reg  signed [31:0] r_run_copy0_j_57;
	reg                r_sub09_run_req;
	wire               w_sub09_run_busy;
	wire signed [12:0] w_sub09_u_addr;
	reg  signed [12:0] r_sub09_u_addr;
	wire        [31:0] w_sub09_u_datain;
	reg         [31:0] r_sub09_u_datain;
	wire        [31:0] w_sub09_u_dataout;
	wire               w_sub09_u_r_w;
	reg                r_sub09_u_r_w;
	wire signed [12:0] w_sub09_result_addr;
	reg  signed [12:0] r_sub09_result_addr;
	wire        [31:0] w_sub09_result_datain;
	reg         [31:0] r_sub09_result_datain;
	wire        [31:0] w_sub09_result_dataout;
	wire               w_sub09_result_r_w;
	reg                r_sub09_result_r_w;
	reg                r_sub08_run_req;
	wire               w_sub08_run_busy;
	wire signed [12:0] w_sub08_u_addr;
	reg  signed [12:0] r_sub08_u_addr;
	wire        [31:0] w_sub08_u_datain;
	reg         [31:0] r_sub08_u_datain;
	wire        [31:0] w_sub08_u_dataout;
	wire               w_sub08_u_r_w;
	reg                r_sub08_u_r_w;
	wire signed [12:0] w_sub08_result_addr;
	reg  signed [12:0] r_sub08_result_addr;
	wire        [31:0] w_sub08_result_datain;
	reg         [31:0] r_sub08_result_datain;
	wire        [31:0] w_sub08_result_dataout;
	wire               w_sub08_result_r_w;
	reg                r_sub08_result_r_w;
	reg                r_sub12_run_req;
	wire               w_sub12_run_busy;
	wire signed [12:0] w_sub12_u_addr;
	reg  signed [12:0] r_sub12_u_addr;
	wire        [31:0] w_sub12_u_datain;
	reg         [31:0] r_sub12_u_datain;
	wire        [31:0] w_sub12_u_dataout;
	wire               w_sub12_u_r_w;
	reg                r_sub12_u_r_w;
	wire signed [12:0] w_sub12_result_addr;
	reg  signed [12:0] r_sub12_result_addr;
	wire        [31:0] w_sub12_result_datain;
	reg         [31:0] r_sub12_result_datain;
	wire        [31:0] w_sub12_result_dataout;
	wire               w_sub12_result_r_w;
	reg                r_sub12_result_r_w;
	reg                r_sub03_run_req;
	wire               w_sub03_run_busy;
	wire signed [12:0] w_sub03_u_addr;
	reg  signed [12:0] r_sub03_u_addr;
	wire        [31:0] w_sub03_u_datain;
	reg         [31:0] r_sub03_u_datain;
	wire        [31:0] w_sub03_u_dataout;
	wire               w_sub03_u_r_w;
	reg                r_sub03_u_r_w;
	wire signed [12:0] w_sub03_result_addr;
	reg  signed [12:0] r_sub03_result_addr;
	wire        [31:0] w_sub03_result_datain;
	reg         [31:0] r_sub03_result_datain;
	wire        [31:0] w_sub03_result_dataout;
	wire               w_sub03_result_r_w;
	reg                r_sub03_result_r_w;
	reg                r_sub02_run_req;
	wire               w_sub02_run_busy;
	wire signed [12:0] w_sub02_u_addr;
	reg  signed [12:0] r_sub02_u_addr;
	wire        [31:0] w_sub02_u_datain;
	reg         [31:0] r_sub02_u_datain;
	wire        [31:0] w_sub02_u_dataout;
	wire               w_sub02_u_r_w;
	reg                r_sub02_u_r_w;
	wire signed [12:0] w_sub02_result_addr;
	reg  signed [12:0] r_sub02_result_addr;
	wire        [31:0] w_sub02_result_datain;
	reg         [31:0] r_sub02_result_datain;
	wire        [31:0] w_sub02_result_dataout;
	wire               w_sub02_result_r_w;
	reg                r_sub02_result_r_w;
	reg                r_sub11_run_req;
	wire               w_sub11_run_busy;
	wire signed [12:0] w_sub11_u_addr;
	reg  signed [12:0] r_sub11_u_addr;
	wire        [31:0] w_sub11_u_datain;
	reg         [31:0] r_sub11_u_datain;
	wire        [31:0] w_sub11_u_dataout;
	wire               w_sub11_u_r_w;
	reg                r_sub11_u_r_w;
	wire signed [12:0] w_sub11_result_addr;
	reg  signed [12:0] r_sub11_result_addr;
	wire        [31:0] w_sub11_result_datain;
	reg         [31:0] r_sub11_result_datain;
	wire        [31:0] w_sub11_result_dataout;
	wire               w_sub11_result_r_w;
	reg                r_sub11_result_r_w;
	reg                r_sub14_run_req;
	wire               w_sub14_run_busy;
	wire signed [12:0] w_sub14_u_addr;
	reg  signed [12:0] r_sub14_u_addr;
	wire        [31:0] w_sub14_u_datain;
	reg         [31:0] r_sub14_u_datain;
	wire        [31:0] w_sub14_u_dataout;
	wire               w_sub14_u_r_w;
	reg                r_sub14_u_r_w;
	wire signed [12:0] w_sub14_result_addr;
	reg  signed [12:0] r_sub14_result_addr;
	wire        [31:0] w_sub14_result_datain;
	reg         [31:0] r_sub14_result_datain;
	wire        [31:0] w_sub14_result_dataout;
	wire               w_sub14_result_r_w;
	reg                r_sub14_result_r_w;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [12:0] w_sub01_u_addr;
	reg  signed [12:0] r_sub01_u_addr;
	wire        [31:0] w_sub01_u_datain;
	reg         [31:0] r_sub01_u_datain;
	wire        [31:0] w_sub01_u_dataout;
	wire               w_sub01_u_r_w;
	reg                r_sub01_u_r_w;
	wire signed [12:0] w_sub01_result_addr;
	reg  signed [12:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub13_run_req;
	wire               w_sub13_run_busy;
	wire signed [12:0] w_sub13_u_addr;
	reg  signed [12:0] r_sub13_u_addr;
	wire        [31:0] w_sub13_u_datain;
	reg         [31:0] r_sub13_u_datain;
	wire        [31:0] w_sub13_u_dataout;
	wire               w_sub13_u_r_w;
	reg                r_sub13_u_r_w;
	wire signed [12:0] w_sub13_result_addr;
	reg  signed [12:0] r_sub13_result_addr;
	wire        [31:0] w_sub13_result_datain;
	reg         [31:0] r_sub13_result_datain;
	wire        [31:0] w_sub13_result_dataout;
	wire               w_sub13_result_r_w;
	reg                r_sub13_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [12:0] w_sub00_u_addr;
	reg  signed [12:0] r_sub00_u_addr;
	wire        [31:0] w_sub00_u_datain;
	reg         [31:0] r_sub00_u_datain;
	wire        [31:0] w_sub00_u_dataout;
	wire               w_sub00_u_r_w;
	reg                r_sub00_u_r_w;
	wire signed [12:0] w_sub00_result_addr;
	reg  signed [12:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	reg                r_sub07_run_req;
	wire               w_sub07_run_busy;
	wire signed [12:0] w_sub07_u_addr;
	reg  signed [12:0] r_sub07_u_addr;
	wire        [31:0] w_sub07_u_datain;
	reg         [31:0] r_sub07_u_datain;
	wire        [31:0] w_sub07_u_dataout;
	wire               w_sub07_u_r_w;
	reg                r_sub07_u_r_w;
	wire signed [12:0] w_sub07_result_addr;
	reg  signed [12:0] r_sub07_result_addr;
	wire        [31:0] w_sub07_result_datain;
	reg         [31:0] r_sub07_result_datain;
	wire        [31:0] w_sub07_result_dataout;
	wire               w_sub07_result_r_w;
	reg                r_sub07_result_r_w;
	reg                r_sub06_run_req;
	wire               w_sub06_run_busy;
	wire signed [12:0] w_sub06_u_addr;
	reg  signed [12:0] r_sub06_u_addr;
	wire        [31:0] w_sub06_u_datain;
	reg         [31:0] r_sub06_u_datain;
	wire        [31:0] w_sub06_u_dataout;
	wire               w_sub06_u_r_w;
	reg                r_sub06_u_r_w;
	wire signed [12:0] w_sub06_result_addr;
	reg  signed [12:0] r_sub06_result_addr;
	wire        [31:0] w_sub06_result_datain;
	reg         [31:0] r_sub06_result_datain;
	wire        [31:0] w_sub06_result_dataout;
	wire               w_sub06_result_r_w;
	reg                r_sub06_result_r_w;
	reg                r_sub15_run_req;
	wire               w_sub15_run_busy;
	wire signed [12:0] w_sub15_u_addr;
	reg  signed [12:0] r_sub15_u_addr;
	wire        [31:0] w_sub15_u_datain;
	reg         [31:0] r_sub15_u_datain;
	wire        [31:0] w_sub15_u_dataout;
	wire               w_sub15_u_r_w;
	reg                r_sub15_u_r_w;
	wire signed [12:0] w_sub15_result_addr;
	reg  signed [12:0] r_sub15_result_addr;
	wire        [31:0] w_sub15_result_datain;
	reg         [31:0] r_sub15_result_datain;
	wire        [31:0] w_sub15_result_dataout;
	wire               w_sub15_result_r_w;
	reg                r_sub15_result_r_w;
	reg                r_sub05_run_req;
	wire               w_sub05_run_busy;
	wire signed [12:0] w_sub05_u_addr;
	reg  signed [12:0] r_sub05_u_addr;
	wire        [31:0] w_sub05_u_datain;
	reg         [31:0] r_sub05_u_datain;
	wire        [31:0] w_sub05_u_dataout;
	wire               w_sub05_u_r_w;
	reg                r_sub05_u_r_w;
	wire signed [12:0] w_sub05_result_addr;
	reg  signed [12:0] r_sub05_result_addr;
	wire        [31:0] w_sub05_result_datain;
	reg         [31:0] r_sub05_result_datain;
	wire        [31:0] w_sub05_result_dataout;
	wire               w_sub05_result_r_w;
	reg                r_sub05_result_r_w;
	reg                r_sub04_run_req;
	wire               w_sub04_run_busy;
	wire signed [12:0] w_sub04_u_addr;
	reg  signed [12:0] r_sub04_u_addr;
	wire        [31:0] w_sub04_u_datain;
	reg         [31:0] r_sub04_u_datain;
	wire        [31:0] w_sub04_u_dataout;
	wire               w_sub04_u_r_w;
	reg                r_sub04_u_r_w;
	wire signed [12:0] w_sub04_result_addr;
	reg  signed [12:0] r_sub04_result_addr;
	wire        [31:0] w_sub04_result_datain;
	reg         [31:0] r_sub04_result_datain;
	wire        [31:0] w_sub04_result_dataout;
	wire               w_sub04_result_r_w;
	reg                r_sub04_result_r_w;
	reg                r_sub10_run_req;
	wire               w_sub10_run_busy;
	wire signed [12:0] w_sub10_u_addr;
	reg  signed [12:0] r_sub10_u_addr;
	wire        [31:0] w_sub10_u_datain;
	reg         [31:0] r_sub10_u_datain;
	wire        [31:0] w_sub10_u_dataout;
	wire               w_sub10_u_r_w;
	reg                r_sub10_u_r_w;
	wire signed [12:0] w_sub10_result_addr;
	reg  signed [12:0] r_sub10_result_addr;
	wire        [31:0] w_sub10_result_datain;
	reg         [31:0] r_sub10_result_datain;
	wire        [31:0] w_sub10_result_dataout;
	wire               w_sub10_result_r_w;
	reg                r_sub10_result_r_w;
	wire signed [31:0] w_sys_tmp1;
	wire               w_sys_tmp3;
	wire               w_sys_tmp4;
	wire signed [31:0] w_sys_tmp5;
	wire               w_sys_tmp6;
	wire               w_sys_tmp7;
	wire signed [31:0] w_sys_tmp10;
	wire signed [31:0] w_sys_tmp11;
	wire signed [31:0] w_sys_tmp12;
	wire        [31:0] w_sys_tmp13;
	wire signed [31:0] w_sys_tmp14;
	wire               w_sys_tmp51;
	wire               w_sys_tmp52;
	wire signed [31:0] w_sys_tmp53;
	wire               w_sys_tmp54;
	wire               w_sys_tmp55;
	wire signed [31:0] w_sys_tmp58;
	wire signed [31:0] w_sys_tmp59;
	wire        [31:0] w_sys_tmp60;
	wire signed [31:0] w_sys_tmp62;
	wire signed [31:0] w_sys_tmp63;
	wire        [31:0] w_sys_tmp64;
	wire signed [31:0] w_sys_tmp66;
	wire signed [31:0] w_sys_tmp67;
	wire        [31:0] w_sys_tmp69;
	wire signed [31:0] w_sys_tmp71;
	wire signed [31:0] w_sys_tmp72;
	wire signed [31:0] w_sys_tmp75;
	wire signed [31:0] w_sys_tmp76;
	wire signed [31:0] w_sys_tmp77;
	wire signed [31:0] w_sys_tmp78;
	wire               w_sys_tmp211;
	wire               w_sys_tmp212;
	wire signed [31:0] w_sys_tmp213;
	wire signed [31:0] w_sys_tmp214;
	wire               w_sys_tmp215;
	wire               w_sys_tmp216;
	wire signed [31:0] w_sys_tmp217;
	wire signed [31:0] w_sys_tmp220;
	wire signed [31:0] w_sys_tmp221;
	wire signed [31:0] w_sys_tmp222;
	wire        [31:0] w_sys_tmp223;
	wire signed [31:0] w_sys_tmp224;
	wire signed [31:0] w_sys_tmp225;
	wire signed [31:0] w_sys_tmp227;
	wire signed [31:0] w_sys_tmp228;
	wire signed [31:0] w_sys_tmp289;
	wire               w_sys_tmp290;
	wire               w_sys_tmp291;
	wire signed [31:0] w_sys_tmp292;
	wire signed [31:0] w_sys_tmp295;
	wire signed [31:0] w_sys_tmp296;
	wire signed [31:0] w_sys_tmp297;
	wire signed [31:0] w_sys_tmp298;
	wire signed [31:0] w_sys_tmp299;
	wire        [31:0] w_sys_tmp300;
	wire signed [31:0] w_sys_tmp301;
	wire signed [31:0] w_sys_tmp302;
	wire signed [31:0] w_sys_tmp303;
	wire signed [31:0] w_sys_tmp304;
	wire signed [31:0] w_sys_tmp305;
	wire signed [31:0] w_sys_tmp378;
	wire               w_sys_tmp379;
	wire               w_sys_tmp380;
	wire signed [31:0] w_sys_tmp381;
	wire signed [31:0] w_sys_tmp384;
	wire signed [31:0] w_sys_tmp385;
	wire signed [31:0] w_sys_tmp386;
	wire signed [31:0] w_sys_tmp387;
	wire signed [31:0] w_sys_tmp388;
	wire        [31:0] w_sys_tmp389;
	wire signed [31:0] w_sys_tmp390;
	wire signed [31:0] w_sys_tmp391;
	wire signed [31:0] w_sys_tmp393;
	wire signed [31:0] w_sys_tmp394;
	wire signed [31:0] w_sys_tmp467;
	wire               w_sys_tmp468;
	wire               w_sys_tmp469;
	wire signed [31:0] w_sys_tmp470;
	wire signed [31:0] w_sys_tmp473;
	wire signed [31:0] w_sys_tmp474;
	wire signed [31:0] w_sys_tmp475;
	wire signed [31:0] w_sys_tmp476;
	wire signed [31:0] w_sys_tmp477;
	wire        [31:0] w_sys_tmp478;
	wire signed [31:0] w_sys_tmp479;
	wire signed [31:0] w_sys_tmp480;
	wire signed [31:0] w_sys_tmp482;
	wire signed [31:0] w_sys_tmp483;
	wire signed [31:0] w_sys_tmp556;
	wire               w_sys_tmp557;
	wire               w_sys_tmp558;
	wire signed [31:0] w_sys_tmp559;
	wire signed [31:0] w_sys_tmp560;
	wire               w_sys_tmp561;
	wire               w_sys_tmp562;
	wire signed [31:0] w_sys_tmp563;
	wire signed [31:0] w_sys_tmp566;
	wire signed [31:0] w_sys_tmp567;
	wire signed [31:0] w_sys_tmp568;
	wire        [31:0] w_sys_tmp569;
	wire signed [31:0] w_sys_tmp570;
	wire signed [31:0] w_sys_tmp571;
	wire signed [31:0] w_sys_tmp573;
	wire signed [31:0] w_sys_tmp574;
	wire signed [31:0] w_sys_tmp635;
	wire               w_sys_tmp636;
	wire               w_sys_tmp637;
	wire signed [31:0] w_sys_tmp638;
	wire signed [31:0] w_sys_tmp641;
	wire signed [31:0] w_sys_tmp642;
	wire signed [31:0] w_sys_tmp643;
	wire signed [31:0] w_sys_tmp644;
	wire signed [31:0] w_sys_tmp645;
	wire        [31:0] w_sys_tmp646;
	wire signed [31:0] w_sys_tmp647;
	wire signed [31:0] w_sys_tmp648;
	wire signed [31:0] w_sys_tmp650;
	wire signed [31:0] w_sys_tmp651;
	wire signed [31:0] w_sys_tmp724;
	wire               w_sys_tmp725;
	wire               w_sys_tmp726;
	wire signed [31:0] w_sys_tmp727;
	wire signed [31:0] w_sys_tmp730;
	wire signed [31:0] w_sys_tmp731;
	wire signed [31:0] w_sys_tmp732;
	wire signed [31:0] w_sys_tmp733;
	wire signed [31:0] w_sys_tmp734;
	wire        [31:0] w_sys_tmp735;
	wire signed [31:0] w_sys_tmp736;
	wire signed [31:0] w_sys_tmp737;
	wire signed [31:0] w_sys_tmp739;
	wire signed [31:0] w_sys_tmp740;
	wire signed [31:0] w_sys_tmp813;
	wire               w_sys_tmp814;
	wire               w_sys_tmp815;
	wire signed [31:0] w_sys_tmp816;
	wire signed [31:0] w_sys_tmp819;
	wire signed [31:0] w_sys_tmp820;
	wire signed [31:0] w_sys_tmp821;
	wire signed [31:0] w_sys_tmp822;
	wire signed [31:0] w_sys_tmp823;
	wire        [31:0] w_sys_tmp824;
	wire signed [31:0] w_sys_tmp825;
	wire signed [31:0] w_sys_tmp826;
	wire signed [31:0] w_sys_tmp828;
	wire signed [31:0] w_sys_tmp829;
	wire signed [31:0] w_sys_tmp902;
	wire               w_sys_tmp903;
	wire               w_sys_tmp904;
	wire signed [31:0] w_sys_tmp905;
	wire signed [31:0] w_sys_tmp906;
	wire               w_sys_tmp907;
	wire               w_sys_tmp908;
	wire signed [31:0] w_sys_tmp909;
	wire signed [31:0] w_sys_tmp912;
	wire signed [31:0] w_sys_tmp913;
	wire signed [31:0] w_sys_tmp914;
	wire        [31:0] w_sys_tmp915;
	wire signed [31:0] w_sys_tmp916;
	wire signed [31:0] w_sys_tmp917;
	wire signed [31:0] w_sys_tmp919;
	wire signed [31:0] w_sys_tmp920;
	wire signed [31:0] w_sys_tmp981;
	wire               w_sys_tmp982;
	wire               w_sys_tmp983;
	wire signed [31:0] w_sys_tmp984;
	wire signed [31:0] w_sys_tmp987;
	wire signed [31:0] w_sys_tmp988;
	wire signed [31:0] w_sys_tmp989;
	wire signed [31:0] w_sys_tmp990;
	wire signed [31:0] w_sys_tmp991;
	wire        [31:0] w_sys_tmp992;
	wire signed [31:0] w_sys_tmp993;
	wire signed [31:0] w_sys_tmp994;
	wire signed [31:0] w_sys_tmp996;
	wire signed [31:0] w_sys_tmp997;
	wire signed [31:0] w_sys_tmp1070;
	wire               w_sys_tmp1071;
	wire               w_sys_tmp1072;
	wire signed [31:0] w_sys_tmp1073;
	wire signed [31:0] w_sys_tmp1076;
	wire signed [31:0] w_sys_tmp1077;
	wire signed [31:0] w_sys_tmp1078;
	wire signed [31:0] w_sys_tmp1079;
	wire signed [31:0] w_sys_tmp1080;
	wire        [31:0] w_sys_tmp1081;
	wire signed [31:0] w_sys_tmp1082;
	wire signed [31:0] w_sys_tmp1083;
	wire signed [31:0] w_sys_tmp1085;
	wire signed [31:0] w_sys_tmp1086;
	wire signed [31:0] w_sys_tmp1159;
	wire               w_sys_tmp1160;
	wire               w_sys_tmp1161;
	wire signed [31:0] w_sys_tmp1162;
	wire signed [31:0] w_sys_tmp1165;
	wire signed [31:0] w_sys_tmp1166;
	wire signed [31:0] w_sys_tmp1167;
	wire signed [31:0] w_sys_tmp1168;
	wire signed [31:0] w_sys_tmp1169;
	wire        [31:0] w_sys_tmp1170;
	wire signed [31:0] w_sys_tmp1171;
	wire signed [31:0] w_sys_tmp1172;
	wire signed [31:0] w_sys_tmp1174;
	wire signed [31:0] w_sys_tmp1175;
	wire signed [31:0] w_sys_tmp1248;
	wire               w_sys_tmp1249;
	wire               w_sys_tmp1250;
	wire signed [31:0] w_sys_tmp1251;
	wire signed [31:0] w_sys_tmp1252;
	wire               w_sys_tmp1253;
	wire               w_sys_tmp1254;
	wire signed [31:0] w_sys_tmp1255;
	wire signed [31:0] w_sys_tmp1258;
	wire signed [31:0] w_sys_tmp1259;
	wire signed [31:0] w_sys_tmp1260;
	wire        [31:0] w_sys_tmp1261;
	wire signed [31:0] w_sys_tmp1262;
	wire signed [31:0] w_sys_tmp1263;
	wire signed [31:0] w_sys_tmp1265;
	wire signed [31:0] w_sys_tmp1266;
	wire signed [31:0] w_sys_tmp1327;
	wire               w_sys_tmp1328;
	wire               w_sys_tmp1329;
	wire signed [31:0] w_sys_tmp1330;
	wire signed [31:0] w_sys_tmp1333;
	wire signed [31:0] w_sys_tmp1334;
	wire signed [31:0] w_sys_tmp1335;
	wire signed [31:0] w_sys_tmp1336;
	wire signed [31:0] w_sys_tmp1337;
	wire        [31:0] w_sys_tmp1338;
	wire signed [31:0] w_sys_tmp1339;
	wire signed [31:0] w_sys_tmp1340;
	wire signed [31:0] w_sys_tmp1342;
	wire signed [31:0] w_sys_tmp1343;
	wire signed [31:0] w_sys_tmp1416;
	wire               w_sys_tmp1417;
	wire               w_sys_tmp1418;
	wire signed [31:0] w_sys_tmp1419;
	wire signed [31:0] w_sys_tmp1422;
	wire signed [31:0] w_sys_tmp1423;
	wire signed [31:0] w_sys_tmp1424;
	wire signed [31:0] w_sys_tmp1425;
	wire signed [31:0] w_sys_tmp1426;
	wire        [31:0] w_sys_tmp1427;
	wire signed [31:0] w_sys_tmp1428;
	wire signed [31:0] w_sys_tmp1429;
	wire signed [31:0] w_sys_tmp1431;
	wire signed [31:0] w_sys_tmp1432;
	wire signed [31:0] w_sys_tmp1505;
	wire               w_sys_tmp1506;
	wire               w_sys_tmp1507;
	wire signed [31:0] w_sys_tmp1508;
	wire signed [31:0] w_sys_tmp1511;
	wire signed [31:0] w_sys_tmp1512;
	wire signed [31:0] w_sys_tmp1513;
	wire signed [31:0] w_sys_tmp1514;
	wire signed [31:0] w_sys_tmp1515;
	wire        [31:0] w_sys_tmp1516;
	wire signed [31:0] w_sys_tmp1517;
	wire signed [31:0] w_sys_tmp1518;
	wire signed [31:0] w_sys_tmp1520;
	wire signed [31:0] w_sys_tmp1521;
	wire signed [31:0] w_sys_tmp1594;
	wire               w_sys_tmp1595;
	wire               w_sys_tmp1596;
	wire signed [31:0] w_sys_tmp1597;
	wire signed [31:0] w_sys_tmp1598;
	wire signed [31:0] w_sys_tmp1599;
	wire               w_sys_tmp1600;
	wire               w_sys_tmp1601;
	wire signed [31:0] w_sys_tmp1602;
	wire signed [31:0] w_sys_tmp1605;
	wire signed [31:0] w_sys_tmp1606;
	wire signed [31:0] w_sys_tmp1607;
	wire        [31:0] w_sys_tmp1608;
	wire signed [31:0] w_sys_tmp1609;
	wire signed [31:0] w_sys_tmp1610;
	wire signed [31:0] w_sys_tmp1612;
	wire signed [31:0] w_sys_tmp1613;
	wire signed [31:0] w_sys_tmp1674;
	wire               w_sys_tmp1675;
	wire               w_sys_tmp1676;
	wire signed [31:0] w_sys_tmp1677;
	wire signed [31:0] w_sys_tmp1680;
	wire signed [31:0] w_sys_tmp1681;
	wire signed [31:0] w_sys_tmp1682;
	wire        [31:0] w_sys_tmp1683;
	wire signed [31:0] w_sys_tmp1684;
	wire signed [31:0] w_sys_tmp1685;
	wire signed [31:0] w_sys_tmp1686;
	wire signed [31:0] w_sys_tmp1687;
	wire signed [31:0] w_sys_tmp1689;
	wire signed [31:0] w_sys_tmp1690;
	wire signed [31:0] w_sys_tmp1763;
	wire               w_sys_tmp1764;
	wire               w_sys_tmp1765;
	wire signed [31:0] w_sys_tmp1766;
	wire signed [31:0] w_sys_tmp1769;
	wire signed [31:0] w_sys_tmp1770;
	wire signed [31:0] w_sys_tmp1771;
	wire        [31:0] w_sys_tmp1772;
	wire signed [31:0] w_sys_tmp1773;
	wire signed [31:0] w_sys_tmp1774;
	wire signed [31:0] w_sys_tmp1775;
	wire signed [31:0] w_sys_tmp1776;
	wire signed [31:0] w_sys_tmp1778;
	wire signed [31:0] w_sys_tmp1779;
	wire signed [31:0] w_sys_tmp1852;
	wire               w_sys_tmp1853;
	wire               w_sys_tmp1854;
	wire signed [31:0] w_sys_tmp1855;
	wire signed [31:0] w_sys_tmp1858;
	wire signed [31:0] w_sys_tmp1859;
	wire signed [31:0] w_sys_tmp1860;
	wire        [31:0] w_sys_tmp1861;
	wire signed [31:0] w_sys_tmp1862;
	wire signed [31:0] w_sys_tmp1863;
	wire signed [31:0] w_sys_tmp1864;
	wire signed [31:0] w_sys_tmp1865;
	wire signed [31:0] w_sys_tmp1867;
	wire signed [31:0] w_sys_tmp1868;
	wire signed [31:0] w_sys_tmp1941;
	wire               w_sys_tmp1942;
	wire               w_sys_tmp1943;
	wire signed [31:0] w_sys_tmp1944;
	wire signed [31:0] w_sys_tmp1945;
	wire signed [31:0] w_sys_tmp1946;
	wire               w_sys_tmp1947;
	wire               w_sys_tmp1948;
	wire signed [31:0] w_sys_tmp1949;
	wire signed [31:0] w_sys_tmp1952;
	wire signed [31:0] w_sys_tmp1953;
	wire signed [31:0] w_sys_tmp1954;
	wire        [31:0] w_sys_tmp1955;
	wire signed [31:0] w_sys_tmp1956;
	wire signed [31:0] w_sys_tmp1957;
	wire signed [31:0] w_sys_tmp1959;
	wire signed [31:0] w_sys_tmp1960;
	wire signed [31:0] w_sys_tmp2021;
	wire               w_sys_tmp2022;
	wire               w_sys_tmp2023;
	wire signed [31:0] w_sys_tmp2024;
	wire signed [31:0] w_sys_tmp2027;
	wire signed [31:0] w_sys_tmp2028;
	wire signed [31:0] w_sys_tmp2029;
	wire        [31:0] w_sys_tmp2030;
	wire signed [31:0] w_sys_tmp2031;
	wire signed [31:0] w_sys_tmp2032;
	wire signed [31:0] w_sys_tmp2033;
	wire signed [31:0] w_sys_tmp2034;
	wire signed [31:0] w_sys_tmp2036;
	wire signed [31:0] w_sys_tmp2037;
	wire signed [31:0] w_sys_tmp2110;
	wire               w_sys_tmp2111;
	wire               w_sys_tmp2112;
	wire signed [31:0] w_sys_tmp2113;
	wire signed [31:0] w_sys_tmp2116;
	wire signed [31:0] w_sys_tmp2117;
	wire signed [31:0] w_sys_tmp2118;
	wire        [31:0] w_sys_tmp2119;
	wire signed [31:0] w_sys_tmp2120;
	wire signed [31:0] w_sys_tmp2121;
	wire signed [31:0] w_sys_tmp2122;
	wire signed [31:0] w_sys_tmp2123;
	wire signed [31:0] w_sys_tmp2125;
	wire signed [31:0] w_sys_tmp2126;
	wire signed [31:0] w_sys_tmp2199;
	wire               w_sys_tmp2200;
	wire               w_sys_tmp2201;
	wire signed [31:0] w_sys_tmp2202;
	wire signed [31:0] w_sys_tmp2205;
	wire signed [31:0] w_sys_tmp2206;
	wire signed [31:0] w_sys_tmp2207;
	wire        [31:0] w_sys_tmp2208;
	wire signed [31:0] w_sys_tmp2209;
	wire signed [31:0] w_sys_tmp2210;
	wire signed [31:0] w_sys_tmp2211;
	wire signed [31:0] w_sys_tmp2212;
	wire signed [31:0] w_sys_tmp2214;
	wire signed [31:0] w_sys_tmp2215;
	wire signed [31:0] w_sys_tmp2288;
	wire               w_sys_tmp2289;
	wire               w_sys_tmp2290;
	wire signed [31:0] w_sys_tmp2291;
	wire signed [31:0] w_sys_tmp2292;
	wire signed [31:0] w_sys_tmp2293;
	wire               w_sys_tmp2294;
	wire               w_sys_tmp2295;
	wire signed [31:0] w_sys_tmp2296;
	wire signed [31:0] w_sys_tmp2299;
	wire signed [31:0] w_sys_tmp2300;
	wire signed [31:0] w_sys_tmp2301;
	wire        [31:0] w_sys_tmp2302;
	wire signed [31:0] w_sys_tmp2303;
	wire signed [31:0] w_sys_tmp2304;
	wire signed [31:0] w_sys_tmp2306;
	wire signed [31:0] w_sys_tmp2307;
	wire signed [31:0] w_sys_tmp2368;
	wire               w_sys_tmp2369;
	wire               w_sys_tmp2370;
	wire signed [31:0] w_sys_tmp2371;
	wire signed [31:0] w_sys_tmp2374;
	wire signed [31:0] w_sys_tmp2375;
	wire signed [31:0] w_sys_tmp2376;
	wire        [31:0] w_sys_tmp2377;
	wire signed [31:0] w_sys_tmp2378;
	wire signed [31:0] w_sys_tmp2379;
	wire signed [31:0] w_sys_tmp2380;
	wire signed [31:0] w_sys_tmp2381;
	wire signed [31:0] w_sys_tmp2383;
	wire signed [31:0] w_sys_tmp2384;
	wire signed [31:0] w_sys_tmp2457;
	wire               w_sys_tmp2458;
	wire               w_sys_tmp2459;
	wire signed [31:0] w_sys_tmp2460;
	wire signed [31:0] w_sys_tmp2463;
	wire signed [31:0] w_sys_tmp2464;
	wire signed [31:0] w_sys_tmp2465;
	wire        [31:0] w_sys_tmp2466;
	wire signed [31:0] w_sys_tmp2467;
	wire signed [31:0] w_sys_tmp2468;
	wire signed [31:0] w_sys_tmp2469;
	wire signed [31:0] w_sys_tmp2470;
	wire signed [31:0] w_sys_tmp2472;
	wire signed [31:0] w_sys_tmp2473;
	wire signed [31:0] w_sys_tmp2546;
	wire               w_sys_tmp2547;
	wire               w_sys_tmp2548;
	wire signed [31:0] w_sys_tmp2549;
	wire signed [31:0] w_sys_tmp2552;
	wire signed [31:0] w_sys_tmp2553;
	wire signed [31:0] w_sys_tmp2554;
	wire        [31:0] w_sys_tmp2555;
	wire signed [31:0] w_sys_tmp2556;
	wire signed [31:0] w_sys_tmp2557;
	wire signed [31:0] w_sys_tmp2558;
	wire signed [31:0] w_sys_tmp2559;
	wire signed [31:0] w_sys_tmp2561;
	wire signed [31:0] w_sys_tmp2562;
	wire signed [31:0] w_sys_tmp2635;
	wire               w_sys_tmp2636;
	wire               w_sys_tmp2637;
	wire signed [31:0] w_sys_tmp2638;
	wire signed [31:0] w_sys_tmp2639;
	wire signed [31:0] w_sys_tmp2640;
	wire               w_sys_tmp2641;
	wire               w_sys_tmp2642;
	wire signed [31:0] w_sys_tmp2643;
	wire signed [31:0] w_sys_tmp2646;
	wire signed [31:0] w_sys_tmp2647;
	wire signed [31:0] w_sys_tmp2648;
	wire        [31:0] w_sys_tmp2649;
	wire signed [31:0] w_sys_tmp2650;
	wire signed [31:0] w_sys_tmp2651;
	wire signed [31:0] w_sys_tmp2653;
	wire signed [31:0] w_sys_tmp2654;
	wire signed [31:0] w_sys_tmp2715;
	wire               w_sys_tmp2716;
	wire               w_sys_tmp2717;
	wire signed [31:0] w_sys_tmp2718;
	wire signed [31:0] w_sys_tmp2721;
	wire signed [31:0] w_sys_tmp2722;
	wire signed [31:0] w_sys_tmp2723;
	wire        [31:0] w_sys_tmp2724;
	wire signed [31:0] w_sys_tmp2725;
	wire signed [31:0] w_sys_tmp2726;
	wire signed [31:0] w_sys_tmp2727;
	wire signed [31:0] w_sys_tmp2728;
	wire signed [31:0] w_sys_tmp2730;
	wire signed [31:0] w_sys_tmp2731;
	wire signed [31:0] w_sys_tmp2804;
	wire               w_sys_tmp2805;
	wire               w_sys_tmp2806;
	wire signed [31:0] w_sys_tmp2807;
	wire signed [31:0] w_sys_tmp2810;
	wire signed [31:0] w_sys_tmp2811;
	wire signed [31:0] w_sys_tmp2812;
	wire        [31:0] w_sys_tmp2813;
	wire signed [31:0] w_sys_tmp2814;
	wire signed [31:0] w_sys_tmp2815;
	wire signed [31:0] w_sys_tmp2816;
	wire signed [31:0] w_sys_tmp2817;
	wire signed [31:0] w_sys_tmp2819;
	wire signed [31:0] w_sys_tmp2820;
	wire signed [31:0] w_sys_tmp2893;
	wire               w_sys_tmp2894;
	wire               w_sys_tmp2895;
	wire signed [31:0] w_sys_tmp2896;
	wire signed [31:0] w_sys_tmp2899;
	wire signed [31:0] w_sys_tmp2900;
	wire signed [31:0] w_sys_tmp2901;
	wire        [31:0] w_sys_tmp2902;
	wire signed [31:0] w_sys_tmp2903;
	wire signed [31:0] w_sys_tmp2904;
	wire signed [31:0] w_sys_tmp2905;
	wire signed [31:0] w_sys_tmp2906;
	wire signed [31:0] w_sys_tmp2908;
	wire signed [31:0] w_sys_tmp2909;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 5'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 5'h1);
	assign w_fld_u_0_addr_0 = 15'sh0;
	assign w_fld_u_0_datain_0 = 32'h0;
	assign w_fld_u_0_r_w_0 = 1'h0;
	assign w_fld_u_0_ce_0 = w_sys_ce;
	assign w_fld_u_0_ce_1 = w_sys_ce;
	assign w_sub09_u_addr = ( (|r_sys_processing_methodID) ? r_sub09_u_addr : 13'sh0 ) ;
	assign w_sub09_u_datain = ( (|r_sys_processing_methodID) ? r_sub09_u_datain : 32'h0 ) ;
	assign w_sub09_u_r_w = ( (|r_sys_processing_methodID) ? r_sub09_u_r_w : 1'h0 ) ;
	assign w_sub09_result_addr = ( (|r_sys_processing_methodID) ? r_sub09_result_addr : 13'sh0 ) ;
	assign w_sub09_result_datain = ( (|r_sys_processing_methodID) ? r_sub09_result_datain : 32'h0 ) ;
	assign w_sub09_result_r_w = ( (|r_sys_processing_methodID) ? r_sub09_result_r_w : 1'h0 ) ;
	assign w_sub08_u_addr = ( (|r_sys_processing_methodID) ? r_sub08_u_addr : 13'sh0 ) ;
	assign w_sub08_u_datain = ( (|r_sys_processing_methodID) ? r_sub08_u_datain : 32'h0 ) ;
	assign w_sub08_u_r_w = ( (|r_sys_processing_methodID) ? r_sub08_u_r_w : 1'h0 ) ;
	assign w_sub08_result_addr = ( (|r_sys_processing_methodID) ? r_sub08_result_addr : 13'sh0 ) ;
	assign w_sub08_result_datain = ( (|r_sys_processing_methodID) ? r_sub08_result_datain : 32'h0 ) ;
	assign w_sub08_result_r_w = ( (|r_sys_processing_methodID) ? r_sub08_result_r_w : 1'h0 ) ;
	assign w_sub12_u_addr = ( (|r_sys_processing_methodID) ? r_sub12_u_addr : 13'sh0 ) ;
	assign w_sub12_u_datain = ( (|r_sys_processing_methodID) ? r_sub12_u_datain : 32'h0 ) ;
	assign w_sub12_u_r_w = ( (|r_sys_processing_methodID) ? r_sub12_u_r_w : 1'h0 ) ;
	assign w_sub12_result_addr = ( (|r_sys_processing_methodID) ? r_sub12_result_addr : 13'sh0 ) ;
	assign w_sub12_result_datain = ( (|r_sys_processing_methodID) ? r_sub12_result_datain : 32'h0 ) ;
	assign w_sub12_result_r_w = ( (|r_sys_processing_methodID) ? r_sub12_result_r_w : 1'h0 ) ;
	assign w_sub03_u_addr = ( (|r_sys_processing_methodID) ? r_sub03_u_addr : 13'sh0 ) ;
	assign w_sub03_u_datain = ( (|r_sys_processing_methodID) ? r_sub03_u_datain : 32'h0 ) ;
	assign w_sub03_u_r_w = ( (|r_sys_processing_methodID) ? r_sub03_u_r_w : 1'h0 ) ;
	assign w_sub03_result_addr = ( (|r_sys_processing_methodID) ? r_sub03_result_addr : 13'sh0 ) ;
	assign w_sub03_result_datain = ( (|r_sys_processing_methodID) ? r_sub03_result_datain : 32'h0 ) ;
	assign w_sub03_result_r_w = ( (|r_sys_processing_methodID) ? r_sub03_result_r_w : 1'h0 ) ;
	assign w_sub02_u_addr = ( (|r_sys_processing_methodID) ? r_sub02_u_addr : 13'sh0 ) ;
	assign w_sub02_u_datain = ( (|r_sys_processing_methodID) ? r_sub02_u_datain : 32'h0 ) ;
	assign w_sub02_u_r_w = ( (|r_sys_processing_methodID) ? r_sub02_u_r_w : 1'h0 ) ;
	assign w_sub02_result_addr = ( (|r_sys_processing_methodID) ? r_sub02_result_addr : 13'sh0 ) ;
	assign w_sub02_result_datain = ( (|r_sys_processing_methodID) ? r_sub02_result_datain : 32'h0 ) ;
	assign w_sub02_result_r_w = ( (|r_sys_processing_methodID) ? r_sub02_result_r_w : 1'h0 ) ;
	assign w_sub11_u_addr = ( (|r_sys_processing_methodID) ? r_sub11_u_addr : 13'sh0 ) ;
	assign w_sub11_u_datain = ( (|r_sys_processing_methodID) ? r_sub11_u_datain : 32'h0 ) ;
	assign w_sub11_u_r_w = ( (|r_sys_processing_methodID) ? r_sub11_u_r_w : 1'h0 ) ;
	assign w_sub11_result_addr = ( (|r_sys_processing_methodID) ? r_sub11_result_addr : 13'sh0 ) ;
	assign w_sub11_result_datain = ( (|r_sys_processing_methodID) ? r_sub11_result_datain : 32'h0 ) ;
	assign w_sub11_result_r_w = ( (|r_sys_processing_methodID) ? r_sub11_result_r_w : 1'h0 ) ;
	assign w_sub14_u_addr = ( (|r_sys_processing_methodID) ? r_sub14_u_addr : 13'sh0 ) ;
	assign w_sub14_u_datain = ( (|r_sys_processing_methodID) ? r_sub14_u_datain : 32'h0 ) ;
	assign w_sub14_u_r_w = ( (|r_sys_processing_methodID) ? r_sub14_u_r_w : 1'h0 ) ;
	assign w_sub14_result_addr = ( (|r_sys_processing_methodID) ? r_sub14_result_addr : 13'sh0 ) ;
	assign w_sub14_result_datain = ( (|r_sys_processing_methodID) ? r_sub14_result_datain : 32'h0 ) ;
	assign w_sub14_result_r_w = ( (|r_sys_processing_methodID) ? r_sub14_result_r_w : 1'h0 ) ;
	assign w_sub01_u_addr = ( (|r_sys_processing_methodID) ? r_sub01_u_addr : 13'sh0 ) ;
	assign w_sub01_u_datain = ( (|r_sys_processing_methodID) ? r_sub01_u_datain : 32'h0 ) ;
	assign w_sub01_u_r_w = ( (|r_sys_processing_methodID) ? r_sub01_u_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 13'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub13_u_addr = ( (|r_sys_processing_methodID) ? r_sub13_u_addr : 13'sh0 ) ;
	assign w_sub13_u_datain = ( (|r_sys_processing_methodID) ? r_sub13_u_datain : 32'h0 ) ;
	assign w_sub13_u_r_w = ( (|r_sys_processing_methodID) ? r_sub13_u_r_w : 1'h0 ) ;
	assign w_sub13_result_addr = ( (|r_sys_processing_methodID) ? r_sub13_result_addr : 13'sh0 ) ;
	assign w_sub13_result_datain = ( (|r_sys_processing_methodID) ? r_sub13_result_datain : 32'h0 ) ;
	assign w_sub13_result_r_w = ( (|r_sys_processing_methodID) ? r_sub13_result_r_w : 1'h0 ) ;
	assign w_sub00_u_addr = ( (|r_sys_processing_methodID) ? r_sub00_u_addr : 13'sh0 ) ;
	assign w_sub00_u_datain = ( (|r_sys_processing_methodID) ? r_sub00_u_datain : 32'h0 ) ;
	assign w_sub00_u_r_w = ( (|r_sys_processing_methodID) ? r_sub00_u_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 13'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sub07_u_addr = ( (|r_sys_processing_methodID) ? r_sub07_u_addr : 13'sh0 ) ;
	assign w_sub07_u_datain = ( (|r_sys_processing_methodID) ? r_sub07_u_datain : 32'h0 ) ;
	assign w_sub07_u_r_w = ( (|r_sys_processing_methodID) ? r_sub07_u_r_w : 1'h0 ) ;
	assign w_sub07_result_addr = ( (|r_sys_processing_methodID) ? r_sub07_result_addr : 13'sh0 ) ;
	assign w_sub07_result_datain = ( (|r_sys_processing_methodID) ? r_sub07_result_datain : 32'h0 ) ;
	assign w_sub07_result_r_w = ( (|r_sys_processing_methodID) ? r_sub07_result_r_w : 1'h0 ) ;
	assign w_sub06_u_addr = ( (|r_sys_processing_methodID) ? r_sub06_u_addr : 13'sh0 ) ;
	assign w_sub06_u_datain = ( (|r_sys_processing_methodID) ? r_sub06_u_datain : 32'h0 ) ;
	assign w_sub06_u_r_w = ( (|r_sys_processing_methodID) ? r_sub06_u_r_w : 1'h0 ) ;
	assign w_sub06_result_addr = ( (|r_sys_processing_methodID) ? r_sub06_result_addr : 13'sh0 ) ;
	assign w_sub06_result_datain = ( (|r_sys_processing_methodID) ? r_sub06_result_datain : 32'h0 ) ;
	assign w_sub06_result_r_w = ( (|r_sys_processing_methodID) ? r_sub06_result_r_w : 1'h0 ) ;
	assign w_sub15_u_addr = ( (|r_sys_processing_methodID) ? r_sub15_u_addr : 13'sh0 ) ;
	assign w_sub15_u_datain = ( (|r_sys_processing_methodID) ? r_sub15_u_datain : 32'h0 ) ;
	assign w_sub15_u_r_w = ( (|r_sys_processing_methodID) ? r_sub15_u_r_w : 1'h0 ) ;
	assign w_sub15_result_addr = ( (|r_sys_processing_methodID) ? r_sub15_result_addr : 13'sh0 ) ;
	assign w_sub15_result_datain = ( (|r_sys_processing_methodID) ? r_sub15_result_datain : 32'h0 ) ;
	assign w_sub15_result_r_w = ( (|r_sys_processing_methodID) ? r_sub15_result_r_w : 1'h0 ) ;
	assign w_sub05_u_addr = ( (|r_sys_processing_methodID) ? r_sub05_u_addr : 13'sh0 ) ;
	assign w_sub05_u_datain = ( (|r_sys_processing_methodID) ? r_sub05_u_datain : 32'h0 ) ;
	assign w_sub05_u_r_w = ( (|r_sys_processing_methodID) ? r_sub05_u_r_w : 1'h0 ) ;
	assign w_sub05_result_addr = ( (|r_sys_processing_methodID) ? r_sub05_result_addr : 13'sh0 ) ;
	assign w_sub05_result_datain = ( (|r_sys_processing_methodID) ? r_sub05_result_datain : 32'h0 ) ;
	assign w_sub05_result_r_w = ( (|r_sys_processing_methodID) ? r_sub05_result_r_w : 1'h0 ) ;
	assign w_sub04_u_addr = ( (|r_sys_processing_methodID) ? r_sub04_u_addr : 13'sh0 ) ;
	assign w_sub04_u_datain = ( (|r_sys_processing_methodID) ? r_sub04_u_datain : 32'h0 ) ;
	assign w_sub04_u_r_w = ( (|r_sys_processing_methodID) ? r_sub04_u_r_w : 1'h0 ) ;
	assign w_sub04_result_addr = ( (|r_sys_processing_methodID) ? r_sub04_result_addr : 13'sh0 ) ;
	assign w_sub04_result_datain = ( (|r_sys_processing_methodID) ? r_sub04_result_datain : 32'h0 ) ;
	assign w_sub04_result_r_w = ( (|r_sys_processing_methodID) ? r_sub04_result_r_w : 1'h0 ) ;
	assign w_sub10_u_addr = ( (|r_sys_processing_methodID) ? r_sub10_u_addr : 13'sh0 ) ;
	assign w_sub10_u_datain = ( (|r_sys_processing_methodID) ? r_sub10_u_datain : 32'h0 ) ;
	assign w_sub10_u_r_w = ( (|r_sys_processing_methodID) ? r_sub10_u_r_w : 1'h0 ) ;
	assign w_sub10_result_addr = ( (|r_sys_processing_methodID) ? r_sub10_result_addr : 13'sh0 ) ;
	assign w_sub10_result_datain = ( (|r_sys_processing_methodID) ? r_sub10_result_datain : 32'h0 ) ;
	assign w_sub10_result_r_w = ( (|r_sys_processing_methodID) ? r_sub10_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh00000081;
	assign w_sys_tmp3 = ( !w_sys_tmp4 );
	assign w_sys_tmp4 = (r_run_my_21 < r_run_k_17);
	assign w_sys_tmp5 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp6 = ( !w_sys_tmp7 );
	assign w_sys_tmp7 = (r_run_mx_20 < r_run_j_18);
	assign w_sys_tmp10 = (w_sys_tmp11 + r_run_k_17);
	assign w_sys_tmp11 = (r_run_j_18 * w_sys_tmp12);
	assign w_sys_tmp12 = 32'sh00000081;
	assign w_sys_tmp13 = 32'h0;
	assign w_sys_tmp14 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp51 = ( !w_sys_tmp52 );
	assign w_sys_tmp52 = (r_run_nlast_22 < r_run_n_19);
	assign w_sys_tmp53 = (r_run_n_19 + w_sys_intOne);
	assign w_sys_tmp54 = ( !w_sys_tmp55 );
	assign w_sys_tmp55 = (r_run_my_21 < r_run_j_18);
	assign w_sys_tmp58 = (w_sys_tmp59 + r_run_j_18);
	assign w_sys_tmp59 = 32'sh00000081;
	assign w_sys_tmp60 = 32'h3f000000;
	assign w_sys_tmp62 = (w_sys_tmp63 + r_run_copy2_j_25);
	assign w_sys_tmp63 = 32'sh00004101;
	assign w_sys_tmp64 = 32'h0;
	assign w_sys_tmp66 = (w_sys_tmp67 + w_sys_intOne);
	assign w_sys_tmp67 = (r_run_copy1_j_24 * w_sys_tmp59);
	assign w_sys_tmp69 = 32'h3f800000;
	assign w_sys_tmp71 = (w_sys_tmp72 + r_run_my_21);
	assign w_sys_tmp72 = (r_run_copy0_j_23 * w_sys_tmp59);
	assign w_sys_tmp75 = (r_run_copy0_j_23 + w_sys_intOne);
	assign w_sys_tmp76 = (r_run_copy1_j_24 + w_sys_intOne);
	assign w_sys_tmp77 = (r_run_copy2_j_25 + w_sys_intOne);
	assign w_sys_tmp78 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp211 = ( !w_sys_tmp212 );
	assign w_sys_tmp212 = (w_sys_tmp213 < r_run_k_17);
	assign w_sys_tmp213 = 32'sh00000021;
	assign w_sys_tmp214 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp215 = ( !w_sys_tmp216 );
	assign w_sys_tmp216 = (w_sys_tmp217 < r_run_j_18);
	assign w_sys_tmp217 = 32'sh00000021;
	assign w_sys_tmp220 = (w_sys_tmp221 + r_run_k_17);
	assign w_sys_tmp221 = (r_run_j_18 * w_sys_tmp222);
	assign w_sys_tmp222 = 32'sh00000081;
	assign w_sys_tmp223 = w_fld_u_0_dataout_1;
	assign w_sys_tmp224 = (w_sys_tmp225 + r_run_k_17);
	assign w_sys_tmp225 = (r_run_copy0_j_26 * w_sys_tmp222);
	assign w_sys_tmp227 = (r_run_copy0_j_26 + w_sys_intOne);
	assign w_sys_tmp228 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp289 = 32'sh00000020;
	assign w_sys_tmp290 = ( !w_sys_tmp291 );
	assign w_sys_tmp291 = (w_sys_tmp292 < r_run_j_18);
	assign w_sys_tmp292 = 32'sh00000041;
	assign w_sys_tmp295 = (w_sys_tmp296 + r_run_k_17);
	assign w_sys_tmp296 = (w_sys_tmp297 * w_sys_tmp299);
	assign w_sys_tmp297 = (r_run_j_18 - w_sys_tmp298);
	assign w_sys_tmp298 = 32'sh0000001f;
	assign w_sys_tmp299 = 32'sh00000081;
	assign w_sys_tmp300 = w_fld_u_0_dataout_1;
	assign w_sys_tmp301 = (w_sys_tmp302 + r_run_k_17);
	assign w_sys_tmp302 = (r_run_copy0_j_27 - w_sys_tmp303);
	assign w_sys_tmp303 = 32'sh00000f9f;
	assign w_sys_tmp304 = (r_run_copy0_j_27 + w_sys_intOne);
	assign w_sys_tmp305 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp378 = 32'sh00000040;
	assign w_sys_tmp379 = ( !w_sys_tmp380 );
	assign w_sys_tmp380 = (w_sys_tmp381 < r_run_j_18);
	assign w_sys_tmp381 = 32'sh00000061;
	assign w_sys_tmp384 = (w_sys_tmp385 + r_run_k_17);
	assign w_sys_tmp385 = (w_sys_tmp386 * w_sys_tmp388);
	assign w_sys_tmp386 = (r_run_j_18 - w_sys_tmp387);
	assign w_sys_tmp387 = 32'sh0000003f;
	assign w_sys_tmp388 = 32'sh00000081;
	assign w_sys_tmp389 = w_fld_u_0_dataout_1;
	assign w_sys_tmp390 = (w_sys_tmp391 + r_run_k_17);
	assign w_sys_tmp391 = (r_run_copy0_j_28 * w_sys_tmp388);
	assign w_sys_tmp393 = (r_run_copy0_j_28 + w_sys_intOne);
	assign w_sys_tmp394 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp467 = 32'sh00000060;
	assign w_sys_tmp468 = ( !w_sys_tmp469 );
	assign w_sys_tmp469 = (w_sys_tmp470 < r_run_j_18);
	assign w_sys_tmp470 = 32'sh00000081;
	assign w_sys_tmp473 = (w_sys_tmp474 + r_run_k_17);
	assign w_sys_tmp474 = (w_sys_tmp475 * w_sys_tmp477);
	assign w_sys_tmp475 = (r_run_j_18 - w_sys_tmp476);
	assign w_sys_tmp476 = 32'sh0000005f;
	assign w_sys_tmp477 = 32'sh00000081;
	assign w_sys_tmp478 = w_fld_u_0_dataout_1;
	assign w_sys_tmp479 = (w_sys_tmp480 + r_run_k_17);
	assign w_sys_tmp480 = (r_run_copy0_j_29 * w_sys_tmp477);
	assign w_sys_tmp482 = (r_run_copy0_j_29 + w_sys_intOne);
	assign w_sys_tmp483 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp556 = 32'sh00000020;
	assign w_sys_tmp557 = ( !w_sys_tmp558 );
	assign w_sys_tmp558 = (w_sys_tmp559 < r_run_k_17);
	assign w_sys_tmp559 = 32'sh00000041;
	assign w_sys_tmp560 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp561 = ( !w_sys_tmp562 );
	assign w_sys_tmp562 = (w_sys_tmp563 < r_run_j_18);
	assign w_sys_tmp563 = 32'sh00000021;
	assign w_sys_tmp566 = (w_sys_tmp567 + r_run_k_17);
	assign w_sys_tmp567 = (r_run_j_18 * w_sys_tmp568);
	assign w_sys_tmp568 = 32'sh00000081;
	assign w_sys_tmp569 = w_fld_u_0_dataout_1;
	assign w_sys_tmp570 = (w_sys_tmp571 + r_run_k_17);
	assign w_sys_tmp571 = (r_run_copy0_j_30 * w_sys_tmp568);
	assign w_sys_tmp573 = (r_run_copy0_j_30 + w_sys_intOne);
	assign w_sys_tmp574 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp635 = 32'sh00000020;
	assign w_sys_tmp636 = ( !w_sys_tmp637 );
	assign w_sys_tmp637 = (w_sys_tmp638 < r_run_j_18);
	assign w_sys_tmp638 = 32'sh00000041;
	assign w_sys_tmp641 = (w_sys_tmp642 + r_run_k_17);
	assign w_sys_tmp642 = (w_sys_tmp643 * w_sys_tmp645);
	assign w_sys_tmp643 = (r_run_j_18 - w_sys_tmp644);
	assign w_sys_tmp644 = 32'sh0000001f;
	assign w_sys_tmp645 = 32'sh00000081;
	assign w_sys_tmp646 = w_fld_u_0_dataout_1;
	assign w_sys_tmp647 = (w_sys_tmp648 + r_run_k_17);
	assign w_sys_tmp648 = (r_run_copy0_j_31 * w_sys_tmp645);
	assign w_sys_tmp650 = (r_run_copy0_j_31 + w_sys_intOne);
	assign w_sys_tmp651 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp724 = 32'sh00000040;
	assign w_sys_tmp725 = ( !w_sys_tmp726 );
	assign w_sys_tmp726 = (w_sys_tmp727 < r_run_j_18);
	assign w_sys_tmp727 = 32'sh00000061;
	assign w_sys_tmp730 = (w_sys_tmp731 + r_run_k_17);
	assign w_sys_tmp731 = (w_sys_tmp732 * w_sys_tmp734);
	assign w_sys_tmp732 = (r_run_j_18 - w_sys_tmp733);
	assign w_sys_tmp733 = 32'sh0000003f;
	assign w_sys_tmp734 = 32'sh00000081;
	assign w_sys_tmp735 = w_fld_u_0_dataout_1;
	assign w_sys_tmp736 = (w_sys_tmp737 + r_run_k_17);
	assign w_sys_tmp737 = (r_run_copy0_j_32 * w_sys_tmp734);
	assign w_sys_tmp739 = (r_run_copy0_j_32 + w_sys_intOne);
	assign w_sys_tmp740 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp813 = 32'sh00000060;
	assign w_sys_tmp814 = ( !w_sys_tmp815 );
	assign w_sys_tmp815 = (w_sys_tmp816 < r_run_j_18);
	assign w_sys_tmp816 = 32'sh00000081;
	assign w_sys_tmp819 = (w_sys_tmp820 + r_run_k_17);
	assign w_sys_tmp820 = (w_sys_tmp821 * w_sys_tmp823);
	assign w_sys_tmp821 = (r_run_j_18 - w_sys_tmp822);
	assign w_sys_tmp822 = 32'sh0000005f;
	assign w_sys_tmp823 = 32'sh00000081;
	assign w_sys_tmp824 = w_fld_u_0_dataout_1;
	assign w_sys_tmp825 = (w_sys_tmp826 + r_run_k_17);
	assign w_sys_tmp826 = (r_run_copy0_j_33 * w_sys_tmp823);
	assign w_sys_tmp828 = (r_run_copy0_j_33 + w_sys_intOne);
	assign w_sys_tmp829 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp902 = 32'sh00000040;
	assign w_sys_tmp903 = ( !w_sys_tmp904 );
	assign w_sys_tmp904 = (w_sys_tmp905 < r_run_k_17);
	assign w_sys_tmp905 = 32'sh00000061;
	assign w_sys_tmp906 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp907 = ( !w_sys_tmp908 );
	assign w_sys_tmp908 = (w_sys_tmp909 < r_run_j_18);
	assign w_sys_tmp909 = 32'sh00000021;
	assign w_sys_tmp912 = (w_sys_tmp913 + r_run_k_17);
	assign w_sys_tmp913 = (r_run_j_18 * w_sys_tmp914);
	assign w_sys_tmp914 = 32'sh00000081;
	assign w_sys_tmp915 = w_fld_u_0_dataout_1;
	assign w_sys_tmp916 = (w_sys_tmp917 + r_run_k_17);
	assign w_sys_tmp917 = (r_run_copy0_j_34 * w_sys_tmp914);
	assign w_sys_tmp919 = (r_run_copy0_j_34 + w_sys_intOne);
	assign w_sys_tmp920 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp981 = 32'sh00000020;
	assign w_sys_tmp982 = ( !w_sys_tmp983 );
	assign w_sys_tmp983 = (w_sys_tmp984 < r_run_j_18);
	assign w_sys_tmp984 = 32'sh00000041;
	assign w_sys_tmp987 = (w_sys_tmp988 + r_run_k_17);
	assign w_sys_tmp988 = (w_sys_tmp989 * w_sys_tmp991);
	assign w_sys_tmp989 = (r_run_j_18 - w_sys_tmp990);
	assign w_sys_tmp990 = 32'sh0000001f;
	assign w_sys_tmp991 = 32'sh00000081;
	assign w_sys_tmp992 = w_fld_u_0_dataout_1;
	assign w_sys_tmp993 = (w_sys_tmp994 + r_run_k_17);
	assign w_sys_tmp994 = (r_run_copy0_j_35 * w_sys_tmp991);
	assign w_sys_tmp996 = (r_run_copy0_j_35 + w_sys_intOne);
	assign w_sys_tmp997 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp1070 = 32'sh00000040;
	assign w_sys_tmp1071 = ( !w_sys_tmp1072 );
	assign w_sys_tmp1072 = (w_sys_tmp1073 < r_run_j_18);
	assign w_sys_tmp1073 = 32'sh00000061;
	assign w_sys_tmp1076 = (w_sys_tmp1077 + r_run_k_17);
	assign w_sys_tmp1077 = (w_sys_tmp1078 * w_sys_tmp1080);
	assign w_sys_tmp1078 = (r_run_j_18 - w_sys_tmp1079);
	assign w_sys_tmp1079 = 32'sh0000003f;
	assign w_sys_tmp1080 = 32'sh00000081;
	assign w_sys_tmp1081 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1082 = (w_sys_tmp1083 + r_run_k_17);
	assign w_sys_tmp1083 = (r_run_copy0_j_36 * w_sys_tmp1080);
	assign w_sys_tmp1085 = (r_run_copy0_j_36 + w_sys_intOne);
	assign w_sys_tmp1086 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp1159 = 32'sh00000060;
	assign w_sys_tmp1160 = ( !w_sys_tmp1161 );
	assign w_sys_tmp1161 = (w_sys_tmp1162 < r_run_j_18);
	assign w_sys_tmp1162 = 32'sh00000081;
	assign w_sys_tmp1165 = (w_sys_tmp1166 + r_run_k_17);
	assign w_sys_tmp1166 = (w_sys_tmp1167 * w_sys_tmp1169);
	assign w_sys_tmp1167 = (r_run_j_18 - w_sys_tmp1168);
	assign w_sys_tmp1168 = 32'sh0000005f;
	assign w_sys_tmp1169 = 32'sh00000081;
	assign w_sys_tmp1170 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1171 = (w_sys_tmp1172 + r_run_k_17);
	assign w_sys_tmp1172 = (r_run_copy0_j_37 * w_sys_tmp1169);
	assign w_sys_tmp1174 = (r_run_copy0_j_37 + w_sys_intOne);
	assign w_sys_tmp1175 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp1248 = 32'sh00000060;
	assign w_sys_tmp1249 = ( !w_sys_tmp1250 );
	assign w_sys_tmp1250 = (w_sys_tmp1251 < r_run_k_17);
	assign w_sys_tmp1251 = 32'sh00000081;
	assign w_sys_tmp1252 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp1253 = ( !w_sys_tmp1254 );
	assign w_sys_tmp1254 = (w_sys_tmp1255 < r_run_j_18);
	assign w_sys_tmp1255 = 32'sh00000021;
	assign w_sys_tmp1258 = (w_sys_tmp1259 + r_run_k_17);
	assign w_sys_tmp1259 = (r_run_j_18 * w_sys_tmp1260);
	assign w_sys_tmp1260 = 32'sh00000081;
	assign w_sys_tmp1261 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1262 = (w_sys_tmp1263 + r_run_k_17);
	assign w_sys_tmp1263 = (r_run_copy0_j_38 * w_sys_tmp1260);
	assign w_sys_tmp1265 = (r_run_copy0_j_38 + w_sys_intOne);
	assign w_sys_tmp1266 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp1327 = 32'sh00000020;
	assign w_sys_tmp1328 = ( !w_sys_tmp1329 );
	assign w_sys_tmp1329 = (w_sys_tmp1330 < r_run_j_18);
	assign w_sys_tmp1330 = 32'sh00000041;
	assign w_sys_tmp1333 = (w_sys_tmp1334 + r_run_k_17);
	assign w_sys_tmp1334 = (w_sys_tmp1335 * w_sys_tmp1337);
	assign w_sys_tmp1335 = (r_run_j_18 - w_sys_tmp1336);
	assign w_sys_tmp1336 = 32'sh0000001f;
	assign w_sys_tmp1337 = 32'sh00000081;
	assign w_sys_tmp1338 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1339 = (w_sys_tmp1340 + r_run_k_17);
	assign w_sys_tmp1340 = (r_run_copy0_j_39 * w_sys_tmp1337);
	assign w_sys_tmp1342 = (r_run_copy0_j_39 + w_sys_intOne);
	assign w_sys_tmp1343 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp1416 = 32'sh00000040;
	assign w_sys_tmp1417 = ( !w_sys_tmp1418 );
	assign w_sys_tmp1418 = (w_sys_tmp1419 < r_run_j_18);
	assign w_sys_tmp1419 = 32'sh00000061;
	assign w_sys_tmp1422 = (w_sys_tmp1423 + r_run_k_17);
	assign w_sys_tmp1423 = (w_sys_tmp1424 * w_sys_tmp1426);
	assign w_sys_tmp1424 = (r_run_j_18 - w_sys_tmp1425);
	assign w_sys_tmp1425 = 32'sh0000003f;
	assign w_sys_tmp1426 = 32'sh00000081;
	assign w_sys_tmp1427 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1428 = (w_sys_tmp1429 + r_run_k_17);
	assign w_sys_tmp1429 = (r_run_copy0_j_40 * w_sys_tmp1426);
	assign w_sys_tmp1431 = (r_run_copy0_j_40 + w_sys_intOne);
	assign w_sys_tmp1432 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp1505 = 32'sh00000060;
	assign w_sys_tmp1506 = ( !w_sys_tmp1507 );
	assign w_sys_tmp1507 = (w_sys_tmp1508 < r_run_j_18);
	assign w_sys_tmp1508 = 32'sh00000081;
	assign w_sys_tmp1511 = (w_sys_tmp1512 + r_run_k_17);
	assign w_sys_tmp1512 = (w_sys_tmp1513 * w_sys_tmp1515);
	assign w_sys_tmp1513 = (r_run_j_18 - w_sys_tmp1514);
	assign w_sys_tmp1514 = 32'sh0000005f;
	assign w_sys_tmp1515 = 32'sh00000081;
	assign w_sys_tmp1516 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1517 = (w_sys_tmp1518 + r_run_k_17);
	assign w_sys_tmp1518 = (r_run_copy0_j_41 * w_sys_tmp1515);
	assign w_sys_tmp1520 = (r_run_copy0_j_41 + w_sys_intOne);
	assign w_sys_tmp1521 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp1594 = 32'sh00000002;
	assign w_sys_tmp1595 = ( !w_sys_tmp1596 );
	assign w_sys_tmp1596 = (w_sys_tmp1597 < r_run_k_17);
	assign w_sys_tmp1597 = 32'sh00000020;
	assign w_sys_tmp1598 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp1599 = 32'sh00000002;
	assign w_sys_tmp1600 = ( !w_sys_tmp1601 );
	assign w_sys_tmp1601 = (w_sys_tmp1602 < r_run_j_18);
	assign w_sys_tmp1602 = 32'sh00000020;
	assign w_sys_tmp1605 = (w_sys_tmp1606 + r_run_k_17);
	assign w_sys_tmp1606 = (r_run_j_18 * w_sys_tmp1607);
	assign w_sys_tmp1607 = 32'sh00000081;
	assign w_sys_tmp1608 = w_sub00_result_dataout;
	assign w_sys_tmp1609 = (w_sys_tmp1610 + r_run_k_17);
	assign w_sys_tmp1610 = (r_run_copy0_j_42 * w_sys_tmp1607);
	assign w_sys_tmp1612 = (r_run_copy0_j_42 + w_sys_intOne);
	assign w_sys_tmp1613 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp1674 = 32'sh00000021;
	assign w_sys_tmp1675 = ( !w_sys_tmp1676 );
	assign w_sys_tmp1676 = (w_sys_tmp1677 < r_run_j_18);
	assign w_sys_tmp1677 = 32'sh00000040;
	assign w_sys_tmp1680 = (w_sys_tmp1681 + r_run_k_17);
	assign w_sys_tmp1681 = (r_run_j_18 * w_sys_tmp1682);
	assign w_sys_tmp1682 = 32'sh00000081;
	assign w_sys_tmp1683 = w_sub01_result_dataout;
	assign w_sys_tmp1684 = (w_sys_tmp1685 + r_run_k_17);
	assign w_sys_tmp1685 = (w_sys_tmp1686 * w_sys_tmp1682);
	assign w_sys_tmp1686 = (r_run_copy0_j_43 - w_sys_tmp1687);
	assign w_sys_tmp1687 = 32'sh0000001f;
	assign w_sys_tmp1689 = (r_run_copy0_j_43 + w_sys_intOne);
	assign w_sys_tmp1690 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp1763 = 32'sh00000041;
	assign w_sys_tmp1764 = ( !w_sys_tmp1765 );
	assign w_sys_tmp1765 = (w_sys_tmp1766 < r_run_j_18);
	assign w_sys_tmp1766 = 32'sh00000060;
	assign w_sys_tmp1769 = (w_sys_tmp1770 + r_run_k_17);
	assign w_sys_tmp1770 = (r_run_j_18 * w_sys_tmp1771);
	assign w_sys_tmp1771 = 32'sh00000081;
	assign w_sys_tmp1772 = w_sub02_result_dataout;
	assign w_sys_tmp1773 = (w_sys_tmp1774 + r_run_k_17);
	assign w_sys_tmp1774 = (w_sys_tmp1775 * w_sys_tmp1771);
	assign w_sys_tmp1775 = (r_run_copy0_j_44 - w_sys_tmp1776);
	assign w_sys_tmp1776 = 32'sh0000003f;
	assign w_sys_tmp1778 = (r_run_copy0_j_44 + w_sys_intOne);
	assign w_sys_tmp1779 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp1852 = 32'sh00000061;
	assign w_sys_tmp1853 = ( !w_sys_tmp1854 );
	assign w_sys_tmp1854 = (w_sys_tmp1855 < r_run_j_18);
	assign w_sys_tmp1855 = 32'sh00000080;
	assign w_sys_tmp1858 = (w_sys_tmp1859 + r_run_k_17);
	assign w_sys_tmp1859 = (r_run_j_18 * w_sys_tmp1860);
	assign w_sys_tmp1860 = 32'sh00000081;
	assign w_sys_tmp1861 = w_sub03_result_dataout;
	assign w_sys_tmp1862 = (w_sys_tmp1863 + r_run_k_17);
	assign w_sys_tmp1863 = (w_sys_tmp1864 * w_sys_tmp1860);
	assign w_sys_tmp1864 = (r_run_copy0_j_45 - w_sys_tmp1865);
	assign w_sys_tmp1865 = 32'sh0000005f;
	assign w_sys_tmp1867 = (r_run_copy0_j_45 + w_sys_intOne);
	assign w_sys_tmp1868 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp1941 = 32'sh00000021;
	assign w_sys_tmp1942 = ( !w_sys_tmp1943 );
	assign w_sys_tmp1943 = (w_sys_tmp1944 < r_run_k_17);
	assign w_sys_tmp1944 = 32'sh00000040;
	assign w_sys_tmp1945 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp1946 = 32'sh00000002;
	assign w_sys_tmp1947 = ( !w_sys_tmp1948 );
	assign w_sys_tmp1948 = (w_sys_tmp1949 < r_run_j_18);
	assign w_sys_tmp1949 = 32'sh00000020;
	assign w_sys_tmp1952 = (w_sys_tmp1953 + r_run_k_17);
	assign w_sys_tmp1953 = (r_run_j_18 * w_sys_tmp1954);
	assign w_sys_tmp1954 = 32'sh00000081;
	assign w_sys_tmp1955 = w_sub04_result_dataout;
	assign w_sys_tmp1956 = (w_sys_tmp1957 + r_run_k_17);
	assign w_sys_tmp1957 = (r_run_copy0_j_46 * w_sys_tmp1954);
	assign w_sys_tmp1959 = (r_run_copy0_j_46 + w_sys_intOne);
	assign w_sys_tmp1960 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp2021 = 32'sh00000021;
	assign w_sys_tmp2022 = ( !w_sys_tmp2023 );
	assign w_sys_tmp2023 = (w_sys_tmp2024 < r_run_j_18);
	assign w_sys_tmp2024 = 32'sh00000040;
	assign w_sys_tmp2027 = (w_sys_tmp2028 + r_run_k_17);
	assign w_sys_tmp2028 = (r_run_j_18 * w_sys_tmp2029);
	assign w_sys_tmp2029 = 32'sh00000081;
	assign w_sys_tmp2030 = w_sub05_result_dataout;
	assign w_sys_tmp2031 = (w_sys_tmp2032 + r_run_k_17);
	assign w_sys_tmp2032 = (w_sys_tmp2033 * w_sys_tmp2029);
	assign w_sys_tmp2033 = (r_run_copy0_j_47 - w_sys_tmp2034);
	assign w_sys_tmp2034 = 32'sh0000001f;
	assign w_sys_tmp2036 = (r_run_copy0_j_47 + w_sys_intOne);
	assign w_sys_tmp2037 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp2110 = 32'sh00000041;
	assign w_sys_tmp2111 = ( !w_sys_tmp2112 );
	assign w_sys_tmp2112 = (w_sys_tmp2113 < r_run_j_18);
	assign w_sys_tmp2113 = 32'sh00000060;
	assign w_sys_tmp2116 = (w_sys_tmp2117 + r_run_k_17);
	assign w_sys_tmp2117 = (r_run_j_18 * w_sys_tmp2118);
	assign w_sys_tmp2118 = 32'sh00000081;
	assign w_sys_tmp2119 = w_sub06_result_dataout;
	assign w_sys_tmp2120 = (w_sys_tmp2121 + r_run_k_17);
	assign w_sys_tmp2121 = (w_sys_tmp2122 * w_sys_tmp2118);
	assign w_sys_tmp2122 = (r_run_copy0_j_48 - w_sys_tmp2123);
	assign w_sys_tmp2123 = 32'sh0000003f;
	assign w_sys_tmp2125 = (r_run_copy0_j_48 + w_sys_intOne);
	assign w_sys_tmp2126 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp2199 = 32'sh00000061;
	assign w_sys_tmp2200 = ( !w_sys_tmp2201 );
	assign w_sys_tmp2201 = (w_sys_tmp2202 < r_run_j_18);
	assign w_sys_tmp2202 = 32'sh00000080;
	assign w_sys_tmp2205 = (w_sys_tmp2206 + r_run_k_17);
	assign w_sys_tmp2206 = (r_run_j_18 * w_sys_tmp2207);
	assign w_sys_tmp2207 = 32'sh00000081;
	assign w_sys_tmp2208 = w_sub07_result_dataout;
	assign w_sys_tmp2209 = (w_sys_tmp2210 + r_run_k_17);
	assign w_sys_tmp2210 = (w_sys_tmp2211 * w_sys_tmp2207);
	assign w_sys_tmp2211 = (r_run_copy0_j_49 - w_sys_tmp2212);
	assign w_sys_tmp2212 = 32'sh0000005f;
	assign w_sys_tmp2214 = (r_run_copy0_j_49 + w_sys_intOne);
	assign w_sys_tmp2215 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp2288 = 32'sh00000041;
	assign w_sys_tmp2289 = ( !w_sys_tmp2290 );
	assign w_sys_tmp2290 = (w_sys_tmp2291 < r_run_k_17);
	assign w_sys_tmp2291 = 32'sh00000060;
	assign w_sys_tmp2292 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp2293 = 32'sh00000002;
	assign w_sys_tmp2294 = ( !w_sys_tmp2295 );
	assign w_sys_tmp2295 = (w_sys_tmp2296 < r_run_j_18);
	assign w_sys_tmp2296 = 32'sh00000020;
	assign w_sys_tmp2299 = (w_sys_tmp2300 + r_run_k_17);
	assign w_sys_tmp2300 = (r_run_j_18 * w_sys_tmp2301);
	assign w_sys_tmp2301 = 32'sh00000081;
	assign w_sys_tmp2302 = w_sub08_result_dataout;
	assign w_sys_tmp2303 = (w_sys_tmp2304 + r_run_k_17);
	assign w_sys_tmp2304 = (r_run_copy0_j_50 * w_sys_tmp2301);
	assign w_sys_tmp2306 = (r_run_copy0_j_50 + w_sys_intOne);
	assign w_sys_tmp2307 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp2368 = 32'sh00000021;
	assign w_sys_tmp2369 = ( !w_sys_tmp2370 );
	assign w_sys_tmp2370 = (w_sys_tmp2371 < r_run_j_18);
	assign w_sys_tmp2371 = 32'sh00000040;
	assign w_sys_tmp2374 = (w_sys_tmp2375 + r_run_k_17);
	assign w_sys_tmp2375 = (r_run_j_18 * w_sys_tmp2376);
	assign w_sys_tmp2376 = 32'sh00000081;
	assign w_sys_tmp2377 = w_sub09_result_dataout;
	assign w_sys_tmp2378 = (w_sys_tmp2379 + r_run_k_17);
	assign w_sys_tmp2379 = (w_sys_tmp2380 * w_sys_tmp2376);
	assign w_sys_tmp2380 = (r_run_copy0_j_51 - w_sys_tmp2381);
	assign w_sys_tmp2381 = 32'sh0000001f;
	assign w_sys_tmp2383 = (r_run_copy0_j_51 + w_sys_intOne);
	assign w_sys_tmp2384 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp2457 = 32'sh00000041;
	assign w_sys_tmp2458 = ( !w_sys_tmp2459 );
	assign w_sys_tmp2459 = (w_sys_tmp2460 < r_run_j_18);
	assign w_sys_tmp2460 = 32'sh00000060;
	assign w_sys_tmp2463 = (w_sys_tmp2464 + r_run_k_17);
	assign w_sys_tmp2464 = (r_run_j_18 * w_sys_tmp2465);
	assign w_sys_tmp2465 = 32'sh00000081;
	assign w_sys_tmp2466 = w_sub10_result_dataout;
	assign w_sys_tmp2467 = (w_sys_tmp2468 + r_run_k_17);
	assign w_sys_tmp2468 = (w_sys_tmp2469 * w_sys_tmp2465);
	assign w_sys_tmp2469 = (r_run_copy0_j_52 - w_sys_tmp2470);
	assign w_sys_tmp2470 = 32'sh0000003f;
	assign w_sys_tmp2472 = (r_run_copy0_j_52 + w_sys_intOne);
	assign w_sys_tmp2473 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp2546 = 32'sh00000061;
	assign w_sys_tmp2547 = ( !w_sys_tmp2548 );
	assign w_sys_tmp2548 = (w_sys_tmp2549 < r_run_j_18);
	assign w_sys_tmp2549 = 32'sh00000080;
	assign w_sys_tmp2552 = (w_sys_tmp2553 + r_run_k_17);
	assign w_sys_tmp2553 = (r_run_j_18 * w_sys_tmp2554);
	assign w_sys_tmp2554 = 32'sh00000081;
	assign w_sys_tmp2555 = w_sub11_result_dataout;
	assign w_sys_tmp2556 = (w_sys_tmp2557 + r_run_k_17);
	assign w_sys_tmp2557 = (w_sys_tmp2558 * w_sys_tmp2554);
	assign w_sys_tmp2558 = (r_run_copy0_j_53 - w_sys_tmp2559);
	assign w_sys_tmp2559 = 32'sh0000005f;
	assign w_sys_tmp2561 = (r_run_copy0_j_53 + w_sys_intOne);
	assign w_sys_tmp2562 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp2635 = 32'sh00000061;
	assign w_sys_tmp2636 = ( !w_sys_tmp2637 );
	assign w_sys_tmp2637 = (w_sys_tmp2638 < r_run_k_17);
	assign w_sys_tmp2638 = 32'sh00000080;
	assign w_sys_tmp2639 = (r_run_k_17 + w_sys_intOne);
	assign w_sys_tmp2640 = 32'sh00000002;
	assign w_sys_tmp2641 = ( !w_sys_tmp2642 );
	assign w_sys_tmp2642 = (w_sys_tmp2643 < r_run_j_18);
	assign w_sys_tmp2643 = 32'sh00000020;
	assign w_sys_tmp2646 = (w_sys_tmp2647 + r_run_k_17);
	assign w_sys_tmp2647 = (r_run_j_18 * w_sys_tmp2648);
	assign w_sys_tmp2648 = 32'sh00000081;
	assign w_sys_tmp2649 = w_sub12_result_dataout;
	assign w_sys_tmp2650 = (w_sys_tmp2651 + r_run_k_17);
	assign w_sys_tmp2651 = (r_run_copy0_j_54 * w_sys_tmp2648);
	assign w_sys_tmp2653 = (r_run_copy0_j_54 + w_sys_intOne);
	assign w_sys_tmp2654 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp2715 = 32'sh00000021;
	assign w_sys_tmp2716 = ( !w_sys_tmp2717 );
	assign w_sys_tmp2717 = (w_sys_tmp2718 < r_run_j_18);
	assign w_sys_tmp2718 = 32'sh00000040;
	assign w_sys_tmp2721 = (w_sys_tmp2722 + r_run_k_17);
	assign w_sys_tmp2722 = (r_run_j_18 * w_sys_tmp2723);
	assign w_sys_tmp2723 = 32'sh00000081;
	assign w_sys_tmp2724 = w_sub13_result_dataout;
	assign w_sys_tmp2725 = (w_sys_tmp2726 + r_run_k_17);
	assign w_sys_tmp2726 = (w_sys_tmp2727 * w_sys_tmp2723);
	assign w_sys_tmp2727 = (r_run_copy0_j_55 - w_sys_tmp2728);
	assign w_sys_tmp2728 = 32'sh0000001f;
	assign w_sys_tmp2730 = (r_run_copy0_j_55 + w_sys_intOne);
	assign w_sys_tmp2731 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp2804 = 32'sh00000041;
	assign w_sys_tmp2805 = ( !w_sys_tmp2806 );
	assign w_sys_tmp2806 = (w_sys_tmp2807 < r_run_j_18);
	assign w_sys_tmp2807 = 32'sh00000060;
	assign w_sys_tmp2810 = (w_sys_tmp2811 + r_run_k_17);
	assign w_sys_tmp2811 = (r_run_j_18 * w_sys_tmp2812);
	assign w_sys_tmp2812 = 32'sh00000081;
	assign w_sys_tmp2813 = w_sub14_result_dataout;
	assign w_sys_tmp2814 = (w_sys_tmp2815 + r_run_k_17);
	assign w_sys_tmp2815 = (w_sys_tmp2816 * w_sys_tmp2812);
	assign w_sys_tmp2816 = (r_run_copy0_j_56 - w_sys_tmp2817);
	assign w_sys_tmp2817 = 32'sh0000003f;
	assign w_sys_tmp2819 = (r_run_copy0_j_56 + w_sys_intOne);
	assign w_sys_tmp2820 = (r_run_j_18 + w_sys_intOne);
	assign w_sys_tmp2893 = 32'sh00000061;
	assign w_sys_tmp2894 = ( !w_sys_tmp2895 );
	assign w_sys_tmp2895 = (w_sys_tmp2896 < r_run_j_18);
	assign w_sys_tmp2896 = 32'sh00000080;
	assign w_sys_tmp2899 = (w_sys_tmp2900 + r_run_k_17);
	assign w_sys_tmp2900 = (r_run_j_18 * w_sys_tmp2901);
	assign w_sys_tmp2901 = 32'sh00000081;
	assign w_sys_tmp2902 = w_sub15_result_dataout;
	assign w_sys_tmp2903 = (w_sys_tmp2904 + r_run_k_17);
	assign w_sys_tmp2904 = (w_sys_tmp2905 * w_sys_tmp2901);
	assign w_sys_tmp2905 = (r_run_copy0_j_57 - w_sys_tmp2906);
	assign w_sys_tmp2906 = 32'sh0000005f;
	assign w_sys_tmp2908 = (r_run_copy0_j_57 + w_sys_intOne);
	assign w_sys_tmp2909 = (r_run_j_18 + w_sys_intOne);


	sub09
		sub09_inst(
			.i_fld_result_1_addr_0 (w_sub09_result_addr),
			.i_fld_result_1_datain_0 (w_sub09_result_datain),
			.o_fld_result_1_dataout_0 (w_sub09_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub09_result_r_w),
			.i_fld_u_0_addr_0 (w_sub09_u_addr),
			.i_fld_u_0_datain_0 (w_sub09_u_datain),
			.o_fld_u_0_dataout_0 (w_sub09_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub09_u_r_w),
			.o_run_busy (w_sub09_run_busy),
			.i_run_req (r_sub09_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub08
		sub08_inst(
			.i_fld_result_1_addr_0 (w_sub08_result_addr),
			.i_fld_result_1_datain_0 (w_sub08_result_datain),
			.o_fld_result_1_dataout_0 (w_sub08_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub08_result_r_w),
			.i_fld_u_0_addr_0 (w_sub08_u_addr),
			.i_fld_u_0_datain_0 (w_sub08_u_datain),
			.o_fld_u_0_dataout_0 (w_sub08_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub08_u_r_w),
			.o_run_busy (w_sub08_run_busy),
			.i_run_req (r_sub08_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub12
		sub12_inst(
			.i_fld_result_1_addr_0 (w_sub12_result_addr),
			.i_fld_result_1_datain_0 (w_sub12_result_datain),
			.o_fld_result_1_dataout_0 (w_sub12_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub12_result_r_w),
			.i_fld_u_0_addr_0 (w_sub12_u_addr),
			.i_fld_u_0_datain_0 (w_sub12_u_datain),
			.o_fld_u_0_dataout_0 (w_sub12_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub12_u_r_w),
			.o_run_busy (w_sub12_run_busy),
			.i_run_req (r_sub12_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub03
		sub03_inst(
			.i_fld_result_1_addr_0 (w_sub03_result_addr),
			.i_fld_result_1_datain_0 (w_sub03_result_datain),
			.o_fld_result_1_dataout_0 (w_sub03_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub03_result_r_w),
			.i_fld_u_0_addr_0 (w_sub03_u_addr),
			.i_fld_u_0_datain_0 (w_sub03_u_datain),
			.o_fld_u_0_dataout_0 (w_sub03_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub03_u_r_w),
			.o_run_busy (w_sub03_run_busy),
			.i_run_req (r_sub03_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub02
		sub02_inst(
			.i_fld_result_1_addr_0 (w_sub02_result_addr),
			.i_fld_result_1_datain_0 (w_sub02_result_datain),
			.o_fld_result_1_dataout_0 (w_sub02_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub02_result_r_w),
			.i_fld_u_0_addr_0 (w_sub02_u_addr),
			.i_fld_u_0_datain_0 (w_sub02_u_datain),
			.o_fld_u_0_dataout_0 (w_sub02_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub02_u_r_w),
			.o_run_busy (w_sub02_run_busy),
			.i_run_req (r_sub02_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub11
		sub11_inst(
			.i_fld_result_1_addr_0 (w_sub11_result_addr),
			.i_fld_result_1_datain_0 (w_sub11_result_datain),
			.o_fld_result_1_dataout_0 (w_sub11_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub11_result_r_w),
			.i_fld_u_0_addr_0 (w_sub11_u_addr),
			.i_fld_u_0_datain_0 (w_sub11_u_datain),
			.o_fld_u_0_dataout_0 (w_sub11_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub11_u_r_w),
			.o_run_busy (w_sub11_run_busy),
			.i_run_req (r_sub11_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub14
		sub14_inst(
			.i_fld_result_1_addr_0 (w_sub14_result_addr),
			.i_fld_result_1_datain_0 (w_sub14_result_datain),
			.o_fld_result_1_dataout_0 (w_sub14_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub14_result_r_w),
			.i_fld_u_0_addr_0 (w_sub14_u_addr),
			.i_fld_u_0_datain_0 (w_sub14_u_datain),
			.o_fld_u_0_dataout_0 (w_sub14_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub14_u_r_w),
			.o_run_busy (w_sub14_run_busy),
			.i_run_req (r_sub14_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub01
		sub01_inst(
			.i_fld_result_1_addr_0 (w_sub01_result_addr),
			.i_fld_result_1_datain_0 (w_sub01_result_datain),
			.o_fld_result_1_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub01_result_r_w),
			.i_fld_u_0_addr_0 (w_sub01_u_addr),
			.i_fld_u_0_datain_0 (w_sub01_u_datain),
			.o_fld_u_0_dataout_0 (w_sub01_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub01_u_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub13
		sub13_inst(
			.i_fld_result_1_addr_0 (w_sub13_result_addr),
			.i_fld_result_1_datain_0 (w_sub13_result_datain),
			.o_fld_result_1_dataout_0 (w_sub13_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub13_result_r_w),
			.i_fld_u_0_addr_0 (w_sub13_u_addr),
			.i_fld_u_0_datain_0 (w_sub13_u_datain),
			.o_fld_u_0_dataout_0 (w_sub13_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub13_u_r_w),
			.o_run_busy (w_sub13_run_busy),
			.i_run_req (r_sub13_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub00
		sub00_inst(
			.i_fld_result_1_addr_0 (w_sub00_result_addr),
			.i_fld_result_1_datain_0 (w_sub00_result_datain),
			.o_fld_result_1_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub00_result_r_w),
			.i_fld_u_0_addr_0 (w_sub00_u_addr),
			.i_fld_u_0_datain_0 (w_sub00_u_datain),
			.o_fld_u_0_dataout_0 (w_sub00_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub00_u_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub07
		sub07_inst(
			.i_fld_result_1_addr_0 (w_sub07_result_addr),
			.i_fld_result_1_datain_0 (w_sub07_result_datain),
			.o_fld_result_1_dataout_0 (w_sub07_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub07_result_r_w),
			.i_fld_u_0_addr_0 (w_sub07_u_addr),
			.i_fld_u_0_datain_0 (w_sub07_u_datain),
			.o_fld_u_0_dataout_0 (w_sub07_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub07_u_r_w),
			.o_run_busy (w_sub07_run_busy),
			.i_run_req (r_sub07_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub06
		sub06_inst(
			.i_fld_result_1_addr_0 (w_sub06_result_addr),
			.i_fld_result_1_datain_0 (w_sub06_result_datain),
			.o_fld_result_1_dataout_0 (w_sub06_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub06_result_r_w),
			.i_fld_u_0_addr_0 (w_sub06_u_addr),
			.i_fld_u_0_datain_0 (w_sub06_u_datain),
			.o_fld_u_0_dataout_0 (w_sub06_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub06_u_r_w),
			.o_run_busy (w_sub06_run_busy),
			.i_run_req (r_sub06_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub15
		sub15_inst(
			.i_fld_result_1_addr_0 (w_sub15_result_addr),
			.i_fld_result_1_datain_0 (w_sub15_result_datain),
			.o_fld_result_1_dataout_0 (w_sub15_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub15_result_r_w),
			.i_fld_u_0_addr_0 (w_sub15_u_addr),
			.i_fld_u_0_datain_0 (w_sub15_u_datain),
			.o_fld_u_0_dataout_0 (w_sub15_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub15_u_r_w),
			.o_run_busy (w_sub15_run_busy),
			.i_run_req (r_sub15_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub05
		sub05_inst(
			.i_fld_result_1_addr_0 (w_sub05_result_addr),
			.i_fld_result_1_datain_0 (w_sub05_result_datain),
			.o_fld_result_1_dataout_0 (w_sub05_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub05_result_r_w),
			.i_fld_u_0_addr_0 (w_sub05_u_addr),
			.i_fld_u_0_datain_0 (w_sub05_u_datain),
			.o_fld_u_0_dataout_0 (w_sub05_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub05_u_r_w),
			.o_run_busy (w_sub05_run_busy),
			.i_run_req (r_sub05_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub04
		sub04_inst(
			.i_fld_result_1_addr_0 (w_sub04_result_addr),
			.i_fld_result_1_datain_0 (w_sub04_result_datain),
			.o_fld_result_1_dataout_0 (w_sub04_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub04_result_r_w),
			.i_fld_u_0_addr_0 (w_sub04_u_addr),
			.i_fld_u_0_datain_0 (w_sub04_u_datain),
			.o_fld_u_0_dataout_0 (w_sub04_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub04_u_r_w),
			.o_run_busy (w_sub04_run_busy),
			.i_run_req (r_sub04_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub10
		sub10_inst(
			.i_fld_result_1_addr_0 (w_sub10_result_addr),
			.i_fld_result_1_datain_0 (w_sub10_result_datain),
			.o_fld_result_1_dataout_0 (w_sub10_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub10_result_r_w),
			.i_fld_u_0_addr_0 (w_sub10_u_addr),
			.i_fld_u_0_datain_0 (w_sub10_u_datain),
			.o_fld_u_0_dataout_0 (w_sub10_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub10_u_r_w),
			.o_run_busy (w_sub10_run_busy),
			.i_run_req (r_sub10_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_u_0(
			.clk (clock),
			.ce_0 (w_fld_u_0_ce_0),
			.addr_0 (w_fld_u_0_addr_0),
			.datain_0 (w_fld_u_0_datain_0),
			.dataout_0 (w_fld_u_0_dataout_0),
			.r_w_0 (w_fld_u_0_r_w_0),
			.ce_1 (w_fld_u_0_ce_1),
			.addr_1 (r_fld_u_0_addr_1),
			.datain_1 (r_fld_u_0_datain_1),
			.dataout_1 (w_fld_u_0_dataout_1),
			.r_w_1 (r_fld_u_0_r_w_1)
		);

	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						9'h105: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 9'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h0: begin
							r_sys_run_phase <= 9'h2;
						end

						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h4;

									end
								end

							endcase
						end

						9'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h5;

									end
								end

							endcase
						end

						9'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3) ? 9'h9 : 9'hf);

									end
								end

							endcase
						end

						9'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h5;

									end
								end

							endcase
						end

						9'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'ha;

									end
								end

							endcase
						end

						9'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6) ? 9'hd : 9'h6);

									end
								end

							endcase
						end

						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h6)) begin
										r_sys_run_phase <= 9'ha;

									end
								end

							endcase
						end

						9'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h10;

									end
								end

							endcase
						end

						9'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp51) ? 9'h14 : 9'h105);

									end
								end

							endcase
						end

						9'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h10;

									end
								end

							endcase
						end

						9'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h15;

									end
								end

							endcase
						end

						9'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp54) ? 9'h18 : 9'h1a);

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h1b)) begin
										r_sys_run_phase <= 9'h15;

									end
								end

							endcase
						end

						9'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h1b;

									end
								end

							endcase
						end

						9'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp211) ? 9'h1f : 9'h37);

									end
								end

							endcase
						end

						9'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h1b;

									end
								end

							endcase
						end

						9'h1f: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h20;

									end
								end

							endcase
						end

						9'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp215) ? 9'h23 : 9'h25);

									end
								end

							endcase
						end

						9'h23: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'h20;

									end
								end

							endcase
						end

						9'h25: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h26;

									end
								end

							endcase
						end

						9'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp290) ? 9'h29 : 9'h2b);

									end
								end

							endcase
						end

						9'h29: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'h26;

									end
								end

							endcase
						end

						9'h2b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h2c;

									end
								end

							endcase
						end

						9'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp379) ? 9'h2f : 9'h31);

									end
								end

							endcase
						end

						9'h2f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'h2c;

									end
								end

							endcase
						end

						9'h31: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h32;

									end
								end

							endcase
						end

						9'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp468) ? 9'h35 : 9'h1c);

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'h32;

									end
								end

							endcase
						end

						9'h37: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h38;

									end
								end

							endcase
						end

						9'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp557) ? 9'h3c : 9'h54);

									end
								end

							endcase
						end

						9'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h38;

									end
								end

							endcase
						end

						9'h3c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h3d;

									end
								end

							endcase
						end

						9'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp561) ? 9'h40 : 9'h42);

									end
								end

							endcase
						end

						9'h40: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'h3d;

									end
								end

							endcase
						end

						9'h42: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h43;

									end
								end

							endcase
						end

						9'h43: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp636) ? 9'h46 : 9'h48);

									end
								end

							endcase
						end

						9'h46: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'h43;

									end
								end

							endcase
						end

						9'h48: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h49;

									end
								end

							endcase
						end

						9'h49: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp725) ? 9'h4c : 9'h4e);

									end
								end

							endcase
						end

						9'h4c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'h49;

									end
								end

							endcase
						end

						9'h4e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h4f;

									end
								end

							endcase
						end

						9'h4f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp814) ? 9'h52 : 9'h39);

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'h4f;

									end
								end

							endcase
						end

						9'h54: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h55;

									end
								end

							endcase
						end

						9'h55: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp903) ? 9'h59 : 9'h71);

									end
								end

							endcase
						end

						9'h56: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h55;

									end
								end

							endcase
						end

						9'h59: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h5a;

									end
								end

							endcase
						end

						9'h5a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp907) ? 9'h5d : 9'h5f);

									end
								end

							endcase
						end

						9'h5d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'h5a;

									end
								end

							endcase
						end

						9'h5f: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h60;

									end
								end

							endcase
						end

						9'h60: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp982) ? 9'h63 : 9'h65);

									end
								end

							endcase
						end

						9'h63: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'h60;

									end
								end

							endcase
						end

						9'h65: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h66;

									end
								end

							endcase
						end

						9'h66: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1071) ? 9'h69 : 9'h6b);

									end
								end

							endcase
						end

						9'h69: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'h66;

									end
								end

							endcase
						end

						9'h6b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h6c;

									end
								end

							endcase
						end

						9'h6c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1160) ? 9'h6f : 9'h56);

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'h6c;

									end
								end

							endcase
						end

						9'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h72;

									end
								end

							endcase
						end

						9'h72: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1249) ? 9'h76 : 9'h8d);

									end
								end

							endcase
						end

						9'h73: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h72;

									end
								end

							endcase
						end

						9'h76: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h77;

									end
								end

							endcase
						end

						9'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1253) ? 9'h7a : 9'h7c);

									end
								end

							endcase
						end

						9'h7a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'h77;

									end
								end

							endcase
						end

						9'h7c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h7d;

									end
								end

							endcase
						end

						9'h7d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1328) ? 9'h80 : 9'h82);

									end
								end

							endcase
						end

						9'h80: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'h7d;

									end
								end

							endcase
						end

						9'h82: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h83;

									end
								end

							endcase
						end

						9'h83: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1417) ? 9'h86 : 9'h88);

									end
								end

							endcase
						end

						9'h86: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'h83;

									end
								end

							endcase
						end

						9'h88: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h89;

									end
								end

							endcase
						end

						9'h89: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1506) ? 9'h8c : 9'h73);

									end
								end

							endcase
						end

						9'h8c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'h89;

									end
								end

							endcase
						end

						9'h8d: begin

							case(r_sys_run_stage) 
								5'h10: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_phase <= 9'h8f;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_phase <= 9'h91;

									end
								end

							endcase
						end

						9'h91: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h92;

									end
								end

							endcase
						end

						9'h92: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1595) ? 9'h96 : 9'hae);

									end
								end

							endcase
						end

						9'h93: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h92;

									end
								end

							endcase
						end

						9'h96: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h97;

									end
								end

							endcase
						end

						9'h97: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1600) ? 9'h9a : 9'h9c);

									end
								end

							endcase
						end

						9'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'h97;

									end
								end

							endcase
						end

						9'h9c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h9d;

									end
								end

							endcase
						end

						9'h9d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1675) ? 9'ha0 : 9'ha2);

									end
								end

							endcase
						end

						9'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'h9d;

									end
								end

							endcase
						end

						9'ha2: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'ha3;

									end
								end

							endcase
						end

						9'ha3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1764) ? 9'ha6 : 9'ha8);

									end
								end

							endcase
						end

						9'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'ha3;

									end
								end

							endcase
						end

						9'ha8: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'ha9;

									end
								end

							endcase
						end

						9'ha9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1853) ? 9'hac : 9'h93);

									end
								end

							endcase
						end

						9'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'ha9;

									end
								end

							endcase
						end

						9'hae: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'haf;

									end
								end

							endcase
						end

						9'haf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1942) ? 9'hb3 : 9'hcb);

									end
								end

							endcase
						end

						9'hb0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'haf;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'hb4;

									end
								end

							endcase
						end

						9'hb4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1947) ? 9'hb7 : 9'hb9);

									end
								end

							endcase
						end

						9'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'hb4;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'hba;

									end
								end

							endcase
						end

						9'hba: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2022) ? 9'hbd : 9'hbf);

									end
								end

							endcase
						end

						9'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'hba;

									end
								end

							endcase
						end

						9'hbf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'hc0;

									end
								end

							endcase
						end

						9'hc0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2111) ? 9'hc3 : 9'hc5);

									end
								end

							endcase
						end

						9'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'hc0;

									end
								end

							endcase
						end

						9'hc5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'hc6;

									end
								end

							endcase
						end

						9'hc6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2200) ? 9'hc9 : 9'hb0);

									end
								end

							endcase
						end

						9'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'hc6;

									end
								end

							endcase
						end

						9'hcb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'hcc;

									end
								end

							endcase
						end

						9'hcc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2289) ? 9'hd0 : 9'he8);

									end
								end

							endcase
						end

						9'hcd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'hcc;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'hd1;

									end
								end

							endcase
						end

						9'hd1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2294) ? 9'hd4 : 9'hd6);

									end
								end

							endcase
						end

						9'hd4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'hd1;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'hd7;

									end
								end

							endcase
						end

						9'hd7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2369) ? 9'hda : 9'hdc);

									end
								end

							endcase
						end

						9'hda: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'hd7;

									end
								end

							endcase
						end

						9'hdc: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'hdd;

									end
								end

							endcase
						end

						9'hdd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2458) ? 9'he0 : 9'he2);

									end
								end

							endcase
						end

						9'he0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'hdd;

									end
								end

							endcase
						end

						9'he2: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'he3;

									end
								end

							endcase
						end

						9'he3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2547) ? 9'he6 : 9'hcd);

									end
								end

							endcase
						end

						9'he6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'he3;

									end
								end

							endcase
						end

						9'he8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'he9;

									end
								end

							endcase
						end

						9'he9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2636) ? 9'hed : 9'h11);

									end
								end

							endcase
						end

						9'hea: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'he9;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'hee;

									end
								end

							endcase
						end

						9'hee: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2641) ? 9'hf1 : 9'hf3);

									end
								end

							endcase
						end

						9'hf1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'hee;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'hf4;

									end
								end

							endcase
						end

						9'hf4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2716) ? 9'hf7 : 9'hf9);

									end
								end

							endcase
						end

						9'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'hf4;

									end
								end

							endcase
						end

						9'hf9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'hfa;

									end
								end

							endcase
						end

						9'hfa: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2805) ? 9'hfd : 9'hff);

									end
								end

							endcase
						end

						9'hfd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'hfa;

									end
								end

							endcase
						end

						9'hff: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 9'h100;

									end
								end

							endcase
						end

						9'h100: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2894) ? 9'h103 : 9'hea);

									end
								end

							endcase
						end

						9'h103: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 9'h100;

									end
								end

							endcase
						end

						9'h105: begin
							r_sys_run_phase <= 9'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 5'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h6)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h1b)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h1f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h23: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h29: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h2b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h2f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h31: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h37: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h40: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h43: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h46: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h48: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h49: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h4c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h4e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h4f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h54: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h55: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h56: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h59: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h5a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h5d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h5f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h60: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h63: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h66: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h69: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h6c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h72: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h73: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h76: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h7a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h7c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h7d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h80: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h83: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h86: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h88: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h89: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h8c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h91: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h92: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h93: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h96: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h97: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h9c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h9d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hae: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'haf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hb0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hb4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hba: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hbf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hc0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hc5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hc6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hcb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hcc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hcd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hda: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hdc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hdd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'he0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'he2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'he3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'he6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'he8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'he9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hea: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hee: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hfa: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hfd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hff: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h100: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h103: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 5'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h6)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h5)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h1b)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h1a)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h1f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h23: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h29: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h2b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h2f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h31: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h37: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h40: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h43: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h46: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h48: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h49: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h4c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h4e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h4f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h54: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h55: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h56: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h59: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h5a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h5d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h5f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h60: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h63: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h66: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h69: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h6c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h72: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h73: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h76: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h7a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h7c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h7d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h80: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h83: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h86: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h88: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h89: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h8c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub00_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub01_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub02_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub03_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub04_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub05_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub06_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub07_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub08_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub09_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub10_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub11_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub12_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub13_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub14_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub15_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

							endcase
						end

						9'h91: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h92: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h93: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h96: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h97: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h9c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h9d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'ha2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'ha3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'ha8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'ha9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hae: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'haf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hb0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hb4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hba: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hbf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hc0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hc5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hc6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hcb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hcc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hcd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hd1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hd4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hd7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hda: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hdc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hdd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'he0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'he2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'he3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'he6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'he8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'he9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hea: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hee: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hf1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hf4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hf9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hfa: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hfd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'hff: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h100: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						9'h103: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						9'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						9'h105: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp10[14:0] );

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0) || (r_sys_run_step==5'h4) || (r_sys_run_step==5'h8) || (r_sys_run_step==5'hc) || (r_sys_run_step==5'h10) || (r_sys_run_step==5'h14) || (r_sys_run_step==5'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp58[14:0] );

									end
									else
									if((r_sys_run_step==5'h1) || (r_sys_run_step==5'h5) || (r_sys_run_step==5'h9) || (r_sys_run_step==5'hd) || (r_sys_run_step==5'h11) || (r_sys_run_step==5'h15) || (r_sys_run_step==5'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp62[14:0] );

									end
									else
									if((r_sys_run_step==5'h3) || (r_sys_run_step==5'h7) || (r_sys_run_step==5'hb) || (r_sys_run_step==5'hf) || (r_sys_run_step==5'h13) || (r_sys_run_step==5'h17) || (r_sys_run_step==5'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp71[14:0] );

									end
									else
									if((r_sys_run_step==5'h2) || (r_sys_run_step==5'h6) || (r_sys_run_step==5'ha) || (r_sys_run_step==5'he) || (r_sys_run_step==5'h12) || (r_sys_run_step==5'h16) || (r_sys_run_step==5'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp66[14:0] );

									end
								end

							endcase
						end

						9'h23: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp224[14:0] );

									end
								end

							endcase
						end

						9'h29: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp301[14:0] );

									end
								end

							endcase
						end

						9'h2f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp390[14:0] );

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp479[14:0] );

									end
								end

							endcase
						end

						9'h40: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp570[14:0] );

									end
								end

							endcase
						end

						9'h46: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp647[14:0] );

									end
								end

							endcase
						end

						9'h4c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp736[14:0] );

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp825[14:0] );

									end
								end

							endcase
						end

						9'h5d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp916[14:0] );

									end
								end

							endcase
						end

						9'h63: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp993[14:0] );

									end
								end

							endcase
						end

						9'h69: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1082[14:0] );

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1171[14:0] );

									end
								end

							endcase
						end

						9'h7a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1262[14:0] );

									end
								end

							endcase
						end

						9'h80: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1339[14:0] );

									end
								end

							endcase
						end

						9'h86: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1428[14:0] );

									end
								end

							endcase
						end

						9'h8c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1517[14:0] );

									end
								end

							endcase
						end

						9'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1605[14:0] );

									end
								end

							endcase
						end

						9'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1680[14:0] );

									end
								end

							endcase
						end

						9'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1769[14:0] );

									end
								end

							endcase
						end

						9'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1858[14:0] );

									end
								end

							endcase
						end

						9'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1952[14:0] );

									end
								end

							endcase
						end

						9'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2027[14:0] );

									end
								end

							endcase
						end

						9'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2116[14:0] );

									end
								end

							endcase
						end

						9'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2205[14:0] );

									end
								end

							endcase
						end

						9'hd4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2299[14:0] );

									end
								end

							endcase
						end

						9'hda: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2374[14:0] );

									end
								end

							endcase
						end

						9'he0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2463[14:0] );

									end
								end

							endcase
						end

						9'he6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2552[14:0] );

									end
								end

							endcase
						end

						9'hf1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2646[14:0] );

									end
								end

							endcase
						end

						9'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2721[14:0] );

									end
								end

							endcase
						end

						9'hfd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2810[14:0] );

									end
								end

							endcase
						end

						9'h103: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2899[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp13;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h2) || (r_sys_run_step==5'h6) || (r_sys_run_step==5'ha) || (r_sys_run_step==5'he) || (r_sys_run_step==5'h12) || (r_sys_run_step==5'h16) || (r_sys_run_step==5'h1a)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp69;

									end
									else
									if((r_sys_run_step==5'h0) || (r_sys_run_step==5'h4) || (r_sys_run_step==5'h8) || (r_sys_run_step==5'hc) || (r_sys_run_step==5'h10) || (r_sys_run_step==5'h14) || (r_sys_run_step==5'h18)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp60;

									end
									else
									if((r_sys_run_step==5'h1) || (r_sys_run_step==5'h3) || (r_sys_run_step==5'h5) || (r_sys_run_step==5'h7) || (r_sys_run_step==5'h9) || (r_sys_run_step==5'hb) || (r_sys_run_step==5'hd) || (r_sys_run_step==5'hf) || (r_sys_run_step==5'h11) || (r_sys_run_step==5'h13) || (r_sys_run_step==5'h15) || (r_sys_run_step==5'h17) || (r_sys_run_step==5'h19) || (r_sys_run_step==5'h1b)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp64;

									end
								end

							endcase
						end

						9'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp1608;

									end
								end

							endcase
						end

						9'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp1683;

									end
								end

							endcase
						end

						9'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp1772;

									end
								end

							endcase
						end

						9'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp1861;

									end
								end

							endcase
						end

						9'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp1955;

									end
								end

							endcase
						end

						9'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp2030;

									end
								end

							endcase
						end

						9'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp2119;

									end
								end

							endcase
						end

						9'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp2208;

									end
								end

							endcase
						end

						9'hd4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp2302;

									end
								end

							endcase
						end

						9'hda: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp2377;

									end
								end

							endcase
						end

						9'he0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp2466;

									end
								end

							endcase
						end

						9'he6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp2555;

									end
								end

							endcase
						end

						9'hf1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp2649;

									end
								end

							endcase
						end

						9'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp2724;

									end
								end

							endcase
						end

						9'hfd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp2813;

									end
								end

							endcase
						end

						9'h103: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp2902;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h1b)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h23: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h29: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h2f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h40: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h46: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h4c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h5d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h63: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h69: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h7a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h80: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h86: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h8c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hd4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hda: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'he0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'he6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hf1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hfd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h103: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h105: begin
							r_fld_u_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_17 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_17 <= w_sys_tmp5;

									end
								end

							endcase
						end

						9'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_17 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_17 <= w_sys_tmp214;

									end
								end

							endcase
						end

						9'h37: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_17 <= w_sys_tmp556;

									end
								end

							endcase
						end

						9'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_17 <= w_sys_tmp560;

									end
								end

							endcase
						end

						9'h54: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_17 <= w_sys_tmp902;

									end
								end

							endcase
						end

						9'h56: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_17 <= w_sys_tmp906;

									end
								end

							endcase
						end

						9'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_17 <= w_sys_tmp1248;

									end
								end

							endcase
						end

						9'h73: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_17 <= w_sys_tmp1252;

									end
								end

							endcase
						end

						9'h91: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_17 <= w_sys_tmp1594;

									end
								end

							endcase
						end

						9'h93: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_17 <= w_sys_tmp1598;

									end
								end

							endcase
						end

						9'hae: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_17 <= w_sys_tmp1941;

									end
								end

							endcase
						end

						9'hb0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_17 <= w_sys_tmp1945;

									end
								end

							endcase
						end

						9'hcb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_17 <= w_sys_tmp2288;

									end
								end

							endcase
						end

						9'hcd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_17 <= w_sys_tmp2292;

									end
								end

							endcase
						end

						9'he8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_17 <= w_sys_tmp2635;

									end
								end

							endcase
						end

						9'hea: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_17 <= w_sys_tmp2639;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_j_18 <= w_sys_tmp14;

									end
								end

							endcase
						end

						9'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0) || (r_sys_run_step==5'h4) || (r_sys_run_step==5'h8) || (r_sys_run_step==5'hc) || (r_sys_run_step==5'h10) || (r_sys_run_step==5'h14) || (r_sys_run_step==5'h18)) begin
										r_run_j_18 <= w_sys_tmp78;

									end
								end

							endcase
						end

						9'h1f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h23: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp228;

									end
								end

							endcase
						end

						9'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_tmp289;

									end
								end

							endcase
						end

						9'h29: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp305;

									end
								end

							endcase
						end

						9'h2b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_tmp378;

									end
								end

							endcase
						end

						9'h2f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp394;

									end
								end

							endcase
						end

						9'h31: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_tmp467;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp483;

									end
								end

							endcase
						end

						9'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h40: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp574;

									end
								end

							endcase
						end

						9'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_tmp635;

									end
								end

							endcase
						end

						9'h46: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp651;

									end
								end

							endcase
						end

						9'h48: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_tmp724;

									end
								end

							endcase
						end

						9'h4c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp740;

									end
								end

							endcase
						end

						9'h4e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_tmp813;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp829;

									end
								end

							endcase
						end

						9'h59: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h5d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp920;

									end
								end

							endcase
						end

						9'h5f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_tmp981;

									end
								end

							endcase
						end

						9'h63: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp997;

									end
								end

							endcase
						end

						9'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_tmp1070;

									end
								end

							endcase
						end

						9'h69: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp1086;

									end
								end

							endcase
						end

						9'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_tmp1159;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp1175;

									end
								end

							endcase
						end

						9'h76: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h7a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp1266;

									end
								end

							endcase
						end

						9'h7c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_tmp1327;

									end
								end

							endcase
						end

						9'h80: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp1343;

									end
								end

							endcase
						end

						9'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_tmp1416;

									end
								end

							endcase
						end

						9'h86: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp1432;

									end
								end

							endcase
						end

						9'h88: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_tmp1505;

									end
								end

							endcase
						end

						9'h8c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp1521;

									end
								end

							endcase
						end

						9'h96: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_tmp1599;

									end
								end

							endcase
						end

						9'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp1613;

									end
								end

							endcase
						end

						9'h9c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_tmp1674;

									end
								end

							endcase
						end

						9'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp1690;

									end
								end

							endcase
						end

						9'ha2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_tmp1763;

									end
								end

							endcase
						end

						9'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp1779;

									end
								end

							endcase
						end

						9'ha8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_tmp1852;

									end
								end

							endcase
						end

						9'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp1868;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_tmp1946;

									end
								end

							endcase
						end

						9'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp1960;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_tmp2021;

									end
								end

							endcase
						end

						9'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp2037;

									end
								end

							endcase
						end

						9'hbf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_tmp2110;

									end
								end

							endcase
						end

						9'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp2126;

									end
								end

							endcase
						end

						9'hc5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_tmp2199;

									end
								end

							endcase
						end

						9'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp2215;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_tmp2293;

									end
								end

							endcase
						end

						9'hd4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp2307;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_tmp2368;

									end
								end

							endcase
						end

						9'hda: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp2384;

									end
								end

							endcase
						end

						9'hdc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_tmp2457;

									end
								end

							endcase
						end

						9'he0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp2473;

									end
								end

							endcase
						end

						9'he2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_tmp2546;

									end
								end

							endcase
						end

						9'he6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp2562;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_tmp2640;

									end
								end

							endcase
						end

						9'hf1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp2654;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_tmp2715;

									end
								end

							endcase
						end

						9'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp2731;

									end
								end

							endcase
						end

						9'hf9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_tmp2804;

									end
								end

							endcase
						end

						9'hfd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp2820;

									end
								end

							endcase
						end

						9'hff: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_18 <= w_sys_tmp2893;

									end
								end

							endcase
						end

						9'h103: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_18 <= w_sys_tmp2909;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_n_19 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_n_19 <= w_sys_tmp53;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_mx_20 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_my_21 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_nlast_22 <= w_sys_intOne;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_23 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h3) || (r_sys_run_step==5'h7) || (r_sys_run_step==5'hb) || (r_sys_run_step==5'hf) || (r_sys_run_step==5'h13) || (r_sys_run_step==5'h17) || (r_sys_run_step==5'h1b)) begin
										r_run_copy0_j_23 <= w_sys_tmp75;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy1_j_24 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h2) || (r_sys_run_step==5'h6) || (r_sys_run_step==5'ha) || (r_sys_run_step==5'he) || (r_sys_run_step==5'h12) || (r_sys_run_step==5'h16) || (r_sys_run_step==5'h1a)) begin
										r_run_copy1_j_24 <= w_sys_tmp76;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy2_j_25 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h1) || (r_sys_run_step==5'h5) || (r_sys_run_step==5'h9) || (r_sys_run_step==5'hd) || (r_sys_run_step==5'h11) || (r_sys_run_step==5'h15) || (r_sys_run_step==5'h19)) begin
										r_run_copy2_j_25 <= w_sys_tmp77;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1f: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_26 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h23: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_26 <= w_sys_tmp227;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h25: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_27 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h29: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_27 <= w_sys_tmp304;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_28 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h2f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_28 <= w_sys_tmp393;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h31: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_29 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_29 <= w_sys_tmp482;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_30 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h40: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_30 <= w_sys_tmp573;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h42: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_31 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h46: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_31 <= w_sys_tmp650;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h48: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_32 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h4c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_32 <= w_sys_tmp739;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h4e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_33 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_33 <= w_sys_tmp828;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h59: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_34 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h5d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_34 <= w_sys_tmp919;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5f: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_35 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h63: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_35 <= w_sys_tmp996;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h65: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_36 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h69: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_36 <= w_sys_tmp1085;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_37 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_37 <= w_sys_tmp1174;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h76: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_38 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h7a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_38 <= w_sys_tmp1265;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_39 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h80: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_39 <= w_sys_tmp1342;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h82: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_40 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h86: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_40 <= w_sys_tmp1431;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h88: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_41 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h8c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_41 <= w_sys_tmp1520;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h96: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_42 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_42 <= w_sys_tmp1612;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_43 <= r_run_j_18;

									end
								end

							endcase
						end

						9'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_43 <= w_sys_tmp1689;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha2: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_44 <= r_run_j_18;

									end
								end

							endcase
						end

						9'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_44 <= w_sys_tmp1778;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha8: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_45 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_45 <= w_sys_tmp1867;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hb3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_46 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_46 <= w_sys_tmp1959;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hb9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_47 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_47 <= w_sys_tmp2036;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hbf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_48 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_48 <= w_sys_tmp2125;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hc5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_49 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_49 <= w_sys_tmp2214;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd0: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_50 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hd4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_50 <= w_sys_tmp2306;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd6: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_51 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hda: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_51 <= w_sys_tmp2383;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hdc: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_52 <= r_run_j_18;

									end
								end

							endcase
						end

						9'he0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_52 <= w_sys_tmp2472;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'he2: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_53 <= r_run_j_18;

									end
								end

							endcase
						end

						9'he6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_53 <= w_sys_tmp2561;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hed: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_54 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hf1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_54 <= w_sys_tmp2653;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hf3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_55 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_55 <= w_sys_tmp2730;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hf9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_56 <= r_run_j_18;

									end
								end

							endcase
						end

						9'hfd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_56 <= w_sys_tmp2819;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hff: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_57 <= r_run_j_18;

									end
								end

							endcase
						end

						9'h103: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_57 <= w_sys_tmp2908;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'h7: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub09_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub09_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h63: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp987[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h63: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub09_u_datain <= w_sys_tmp992;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h63: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub09_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub09_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hda: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp2378[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hda: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub09_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub08_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub08_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp912[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub08_u_datain <= w_sys_tmp915;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub08_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub08_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp2303[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hd4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub08_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'h10: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub12_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub12_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp1258[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub12_u_datain <= w_sys_tmp1261;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub12_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub12_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hf1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp2650[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hf1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub12_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'h3: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp473[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub03_u_datain <= w_sys_tmp478;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub03_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub03_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1862[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub03_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'h2: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp384[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub02_u_datain <= w_sys_tmp389;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub02_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub02_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1773[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub02_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'h9: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub11_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub11_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1165[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub11_u_datain <= w_sys_tmp1170;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub11_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub11_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'he6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp2556[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'he6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub11_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'hb: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub14_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub14_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h86: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp1422[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h86: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub14_u_datain <= w_sys_tmp1427;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h86: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub14_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub14_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hfd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp2814[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hfd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub14_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h29: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp295[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h29: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub01_u_datain <= w_sys_tmp300;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h29: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub01_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub01_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1684[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'ha: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub13_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub13_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h80: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp1333[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h80: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub13_u_datain <= w_sys_tmp1338;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h80: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub13_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub13_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp2725[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub13_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h23: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp220[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h23: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub00_u_datain <= w_sys_tmp223;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h23: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub00_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub00_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1609[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'h6: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub07_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub07_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp819[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub07_u_datain <= w_sys_tmp824;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub07_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub07_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2209[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub07_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'h5: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub06_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub06_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h4c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp730[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h4c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub06_u_datain <= w_sys_tmp735;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h4c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub06_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub06_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2120[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub06_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'hc: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub15_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub15_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp1511[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub15_u_datain <= w_sys_tmp1516;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub15_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub15_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h103: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp2903[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h103: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub15_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'h4: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub05_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub05_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h46: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp641[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h46: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub05_u_datain <= w_sys_tmp646;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h46: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub05_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub05_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2031[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub05_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'he: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub04_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub04_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h40: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp566[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h40: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub04_u_datain <= w_sys_tmp569;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h40: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub04_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub04_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp1956[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub04_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'h8: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub10_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub10_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_u_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h69: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp1076[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h69: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub10_u_datain <= w_sys_tmp1081;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h69: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub10_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub10_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_addr <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'he0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp2467[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'he0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h105: begin
							r_sub10_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


endmodule
