/*
TimeStamp:	2016/12/2		14:42
*/


module Jacobi(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy,	
	output signed  [31:0] o_run_return	
);

	reg         [31:0] r_ip_AddFloat_portA_0;
	reg         [31:0] r_ip_AddFloat_portB_0;
	wire        [31:0] w_ip_AddFloat_result_0;
	reg         [31:0] r_ip_MultFloat_multiplicand_0;
	reg         [31:0] r_ip_MultFloat_multiplier_0;
	wire        [31:0] w_ip_MultFloat_product_0;
	reg         [31:0] r_ip_DivFloat_dividend_0;
	reg         [31:0] r_ip_DivFloat_divisor_0;
	wire        [31:0] w_ip_DivFloat_quotient_0;
	reg         [31:0] r_ip_CompareFloatLT_portA_0;
	reg         [31:0] r_ip_CompareFloatLT_portB_0;
	wire               w_ip_CompareFloatLT_result_0;
	reg  signed [31:0] r_ip_FixedToFloat_fixed_0;
	wire        [31:0] w_ip_FixedToFloat_floating_0;
	reg         [ 2:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [31:0] r_sys_max_return;
	reg         [ 2:0] r_sys_max_caller;
	reg                r_sys_max_req;
	reg         [ 3:0] r_sys_max_phase;
	reg         [ 1:0] r_sys_max_stage;
	reg         [ 2:0] r_sys_max_step;
	reg                r_sys_max_busy;
	wire        [ 1:0] w_sys_max_stage_p1;
	wire        [ 2:0] w_sys_max_step_p1;
	reg         [31:0] r_sys_sqrt_return;
	reg         [ 2:0] r_sys_sqrt_caller;
	reg                r_sys_sqrt_req;
	reg         [ 3:0] r_sys_sqrt_phase;
	reg         [ 1:0] r_sys_sqrt_stage;
	reg         [ 6:0] r_sys_sqrt_step;
	reg                r_sys_sqrt_busy;
	wire        [ 1:0] w_sys_sqrt_stage_p1;
	wire        [ 6:0] w_sys_sqrt_step_p1;
	reg         [31:0] r_sys_run_return;
	reg         [ 2:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 6:0] r_sys_run_phase;
	reg         [ 3:0] r_sys_run_stage;
	reg         [ 5:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 3:0] w_sys_run_stage_p1;
	wire        [ 5:0] w_sys_run_step_p1;
	wire signed [ 3:0] w_fld_a_0_addr_0;
	wire        [31:0] w_fld_a_0_datain_0;
	wire        [31:0] w_fld_a_0_dataout_0;
	wire               w_fld_a_0_r_w_0;
	wire               w_fld_a_0_ce_0;
	reg  signed [ 3:0] r_fld_a_0_addr_1;
	reg         [31:0] r_fld_a_0_datain_1;
	wire        [31:0] w_fld_a_0_dataout_1;
	reg                r_fld_a_0_r_w_1;
	wire               w_fld_a_0_ce_1;
	wire signed [ 3:0] w_fld_x_1_addr_0;
	wire        [31:0] w_fld_x_1_datain_0;
	wire        [31:0] w_fld_x_1_dataout_0;
	wire               w_fld_x_1_r_w_0;
	wire               w_fld_x_1_ce_0;
	reg  signed [ 3:0] r_fld_x_1_addr_1;
	reg         [31:0] r_fld_x_1_datain_1;
	wire        [31:0] w_fld_x_1_dataout_1;
	reg                r_fld_x_1_r_w_1;
	wire               w_fld_x_1_ce_1;
	reg         [31:0] r_max_a_2;
	reg         [31:0] r_max_b_3;
	reg         [31:0] r_sqrt_s_4;
	reg         [31:0] r_sqrt_x_5;
	reg         [31:0] r_sqrt_last_x_6;
	reg  signed [31:0] r_run_i_7;
	reg  signed [31:0] r_run_j_8;
	reg  signed [31:0] r_run_k_9;
	reg  signed [31:0] r_run_n_10;
	reg         [31:0] r_run_abserr_11;
	reg         [31:0] r_run_b2_12;
	reg         [31:0] r_run_bar_13;
	reg         [31:0] r_run_beta_14;
	reg         [31:0] r_run_coeff_15;
	reg         [31:0] r_run_c_16;
	reg         [31:0] r_run_s_17;
	reg         [31:0] r_run_cs_18;
	reg         [31:0] r_run_sc_19;
	reg         [31:0] r_run_tmp_20;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg         [31:0] r_sys_tmp4_float;
	wire               w_sys_tmp1;
	wire        [31:0] w_sys_tmp2;
	wire        [31:0] w_sys_tmp3;
	wire        [31:0] w_sys_tmp4;
	wire        [31:0] w_sys_tmp5;
	wire        [31:0] w_sys_tmp6;
	wire               w_sys_tmp7;
	wire        [31:0] w_sys_tmp8;
	wire        [31:0] w_sys_tmp9;
	wire        [31:0] w_sys_tmp11;
	wire        [31:0] w_sys_tmp12;
	wire signed [31:0] w_sys_tmp13;
	wire        [31:0] w_sys_tmp14;
	wire        [31:0] w_sys_tmp15;
	wire        [31:0] w_sys_tmp17;
	wire        [31:0] w_sys_tmp19;
	wire signed [31:0] w_sys_tmp21;
	wire        [31:0] w_sys_tmp22;
	wire signed [31:0] w_sys_tmp27;
	wire signed [31:0] w_sys_tmp30;
	wire        [31:0] w_sys_tmp31;
	wire signed [31:0] w_sys_tmp33;
	wire signed [31:0] w_sys_tmp36;
	wire signed [31:0] w_sys_tmp39;
	wire        [31:0] w_sys_tmp40;
	wire               w_sys_tmp41;
	wire signed [31:0] w_sys_tmp42;
	wire               w_sys_tmp43;
	wire signed [31:0] w_sys_tmp46;
	wire signed [31:0] w_sys_tmp47;
	wire signed [31:0] w_sys_tmp48;
	wire        [31:0] w_sys_tmp49;
	wire signed [31:0] w_sys_tmp50;
	wire               w_sys_tmp87;
	wire signed [31:0] w_sys_tmp90;
	wire signed [31:0] w_sys_tmp91;
	wire signed [31:0] w_sys_tmp92;
	wire        [31:0] w_sys_tmp93;
	wire signed [31:0] w_sys_tmp94;
	wire               w_sys_tmp95;
	wire signed [31:0] w_sys_tmp96;
	wire               w_sys_tmp97;
	wire signed [31:0] w_sys_tmp98;
	wire               w_sys_tmp99;
	wire        [31:0] w_sys_tmp100;
	wire        [31:0] w_sys_tmp101;
	wire signed [31:0] w_sys_tmp102;
	wire signed [31:0] w_sys_tmp103;
	wire signed [31:0] w_sys_tmp104;
	wire        [31:0] w_sys_tmp105;
	wire               w_sys_tmp109;
	wire               w_sys_tmp110;
	wire        [31:0] w_sys_tmp111;
	wire        [31:0] w_sys_tmp112;
	wire        [31:0] w_sys_tmp113;
	wire        [31:0] w_sys_tmp114;
	wire        [31:0] w_sys_tmp115;
	wire               w_sys_tmp116;
	wire               w_sys_tmp117;
	wire signed [31:0] w_sys_tmp118;
	wire signed [31:0] w_sys_tmp119;
	wire signed [31:0] w_sys_tmp120;
	wire               w_sys_tmp121;
	wire signed [31:0] w_sys_tmp122;
	wire               w_sys_tmp123;
	wire               w_sys_tmp124;
	wire        [31:0] w_sys_tmp125;
	wire signed [31:0] w_sys_tmp126;
	wire signed [31:0] w_sys_tmp127;
	wire signed [31:0] w_sys_tmp128;
	wire        [31:0] w_sys_tmp129;
	wire        [31:0] w_sys_tmp133;
	wire        [31:0] w_sys_tmp134;
	wire        [31:0] w_sys_tmp136;
	wire        [31:0] w_sys_tmp137;
	wire signed [31:0] w_sys_tmp138;
	wire signed [31:0] w_sys_tmp139;
	wire signed [31:0] w_sys_tmp140;
	wire        [31:0] w_sys_tmp144;
	wire        [31:0] w_sys_tmp146;
	wire        [31:0] w_sys_tmp147;
	wire        [31:0] w_sys_tmp148;
	wire signed [31:0] w_sys_tmp150;
	wire signed [31:0] w_sys_tmp151;
	wire signed [31:0] w_sys_tmp154;
	wire        [31:0] w_sys_tmp163;
	wire        [31:0] w_sys_tmp164;
	wire        [31:0] w_sys_tmp165;
	wire        [31:0] w_sys_tmp166;
	wire        [31:0] w_sys_tmp167;
	wire        [31:0] w_sys_tmp168;
	wire        [31:0] w_sys_tmp169;
	wire        [31:0] w_sys_tmp170;
	wire        [31:0] w_sys_tmp171;
	wire        [31:0] w_sys_tmp172;
	wire        [31:0] w_sys_tmp173;
	wire        [31:0] w_sys_tmp174;
	wire               w_sys_tmp175;
	wire        [31:0] w_sys_tmp177;
	wire        [31:0] w_sys_tmp178;
	wire signed [31:0] w_sys_tmp179;
	wire signed [31:0] w_sys_tmp180;
	wire signed [31:0] w_sys_tmp181;
	wire        [31:0] w_sys_tmp182;
	wire signed [31:0] w_sys_tmp184;
	wire signed [31:0] w_sys_tmp185;
	wire        [31:0] w_sys_tmp189;
	wire        [31:0] w_sys_tmp201;
	wire signed [31:0] w_sys_tmp207;
	wire               w_sys_tmp208;
	wire        [31:0] w_sys_tmp210;
	wire        [31:0] w_sys_tmp211;
	wire signed [31:0] w_sys_tmp212;
	wire signed [31:0] w_sys_tmp213;
	wire signed [31:0] w_sys_tmp214;
	wire        [31:0] w_sys_tmp215;
	wire signed [31:0] w_sys_tmp216;
	wire        [31:0] w_sys_tmp220;
	wire        [31:0] w_sys_tmp232;
	wire        [31:0] w_sys_tmp247;
	wire signed [31:0] w_sys_tmp265;
	wire        [31:0] w_sys_tmp266;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign w_sys_max_stage_p1 = (r_sys_max_stage + 2'h1);
	assign w_sys_max_step_p1 = (r_sys_max_step + 3'h1);
	assign w_sys_sqrt_stage_p1 = (r_sys_sqrt_stage + 2'h1);
	assign w_sys_sqrt_step_p1 = (r_sys_sqrt_step + 7'h1);
	assign o_run_busy = r_sys_run_busy;
	assign o_run_return = r_sys_run_return;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 4'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 6'h1);
	assign w_fld_a_0_addr_0 = 4'sh0;
	assign w_fld_a_0_datain_0 = 32'h0;
	assign w_fld_a_0_r_w_0 = 1'h0;
	assign w_fld_a_0_ce_0 = w_sys_ce;
	assign w_fld_a_0_ce_1 = w_sys_ce;
	assign w_fld_x_1_addr_0 = 4'sh0;
	assign w_fld_x_1_datain_0 = 32'h0;
	assign w_fld_x_1_r_w_0 = 1'h0;
	assign w_fld_x_1_ce_0 = w_sys_ce;
	assign w_fld_x_1_ce_1 = w_sys_ce;
	assign w_sys_tmp1 = w_ip_CompareFloatLT_result_0;
	assign w_sys_tmp2 = r_max_a_2;
	assign w_sys_tmp3 = r_max_b_3;
	assign w_sys_tmp4 = w_ip_DivFloat_quotient_0;
	assign w_sys_tmp5 = 32'h40000000;
	assign w_sys_tmp6 = 32'h0;
	assign w_sys_tmp7 = (r_sqrt_x_5 != r_sqrt_last_x_6);
	assign w_sys_tmp8 = w_ip_DivFloat_quotient_0;
	assign w_sys_tmp9 = w_ip_AddFloat_result_0;
	assign w_sys_tmp11 = 32'h40000000;
	assign w_sys_tmp12 = r_sqrt_x_5;
	assign w_sys_tmp13 = 32'sh00000003;
	assign w_sys_tmp14 = 32'h3089705f;
	assign w_sys_tmp15 = 32'h0;
	assign w_sys_tmp17 = 32'h3f800000;
	assign w_sys_tmp19 = 32'h40000000;
	assign w_sys_tmp21 = 32'sh00000002;
	assign w_sys_tmp22 = 32'h40400000;
	assign w_sys_tmp27 = 32'sh00000004;
	assign w_sys_tmp30 = 32'sh00000005;
	assign w_sys_tmp31 = 32'hc0000000;
	assign w_sys_tmp33 = 32'sh00000006;
	assign w_sys_tmp36 = 32'sh00000007;
	assign w_sys_tmp39 = 32'sh00000008;
	assign w_sys_tmp40 = 32'h40800000;
	assign w_sys_tmp41 = (r_run_i_7 < r_run_n_10);
	assign w_sys_tmp42 = (r_run_i_7 + w_sys_intOne);
	assign w_sys_tmp43 = (r_run_j_8 < r_run_n_10);
	assign w_sys_tmp46 = (w_sys_tmp47 + r_run_j_8);
	assign w_sys_tmp47 = (w_sys_tmp48 * r_run_i_7);
	assign w_sys_tmp48 = 32'sh00000003;
	assign w_sys_tmp49 = 32'h0;
	assign w_sys_tmp50 = (r_run_j_8 + w_sys_intOne);
	assign w_sys_tmp87 = (r_run_i_7 < r_run_n_10);
	assign w_sys_tmp90 = (w_sys_tmp91 + r_run_i_7);
	assign w_sys_tmp91 = (w_sys_tmp92 * r_run_i_7);
	assign w_sys_tmp92 = 32'sh00000003;
	assign w_sys_tmp93 = 32'h3f800000;
	assign w_sys_tmp94 = (r_run_i_7 + w_sys_intOne);
	assign w_sys_tmp95 = (r_run_i_7 < r_run_n_10);
	assign w_sys_tmp96 = (r_run_i_7 + w_sys_intOne);
	assign w_sys_tmp97 = (r_run_j_8 < r_run_n_10);
	assign w_sys_tmp98 = (r_run_j_8 + w_sys_intOne);
	assign w_sys_tmp99 = (r_run_i_7 != r_run_j_8);
	assign w_sys_tmp100 = w_ip_AddFloat_result_0;
	assign w_sys_tmp101 = w_ip_MultFloat_product_0;
	assign w_sys_tmp102 = (w_sys_tmp103 + r_run_j_8);
	assign w_sys_tmp103 = (w_sys_tmp104 * r_run_i_7);
	assign w_sys_tmp104 = 32'sh00000003;
	assign w_sys_tmp105 = w_fld_a_0_dataout_1;
	assign w_sys_tmp109 = ( !w_sys_tmp110 );
	assign w_sys_tmp110 = w_ip_CompareFloatLT_result_0;
	assign w_sys_tmp111 = 32'h0;
	assign w_sys_tmp112 = w_ip_DivFloat_quotient_0;
	assign w_sys_tmp113 = 32'h3f000000;
	assign w_sys_tmp114 = w_ip_MultFloat_product_0;
	assign w_sys_tmp115 = w_ip_FixedToFloat_floating_0;
	assign w_sys_tmp116 = w_ip_CompareFloatLT_result_0;
	assign w_sys_tmp117 = (r_run_i_7 < w_sys_tmp118);
	assign w_sys_tmp118 = (r_run_n_10 - w_sys_intOne);
	assign w_sys_tmp119 = (r_run_i_7 + w_sys_intOne);
	assign w_sys_tmp120 = (r_run_i_7 + w_sys_intOne);
	assign w_sys_tmp121 = (r_run_j_8 < r_run_n_10);
	assign w_sys_tmp122 = (r_run_j_8 + w_sys_intOne);
	assign w_sys_tmp123 = ( !w_sys_tmp124 );
	assign w_sys_tmp124 = w_ip_CompareFloatLT_result_0;
	assign w_sys_tmp125 = w_ip_MultFloat_product_0;
	assign w_sys_tmp126 = (w_sys_tmp127 + r_run_j_8);
	assign w_sys_tmp127 = (w_sys_tmp128 * r_run_i_7);
	assign w_sys_tmp128 = 32'sh00000003;
	assign w_sys_tmp129 = w_fld_a_0_dataout_1;
	assign w_sys_tmp133 = w_ip_AddFloat_result_0;
	assign w_sys_tmp134 = w_ip_MultFloat_product_0;
	assign w_sys_tmp136 = 32'h40000000;
	assign w_sys_tmp137 = w_fld_a_0_dataout_1;
	assign w_sys_tmp138 = (w_sys_tmp139 + r_run_j_8);
	assign w_sys_tmp139 = (w_sys_tmp140 * r_run_i_7);
	assign w_sys_tmp140 = 32'sh00000003;
	assign w_sys_tmp144 = w_ip_DivFloat_quotient_0;
	assign w_sys_tmp146 = 32'h3f000000;
	assign w_sys_tmp147 = w_sys_tmp133;
	assign w_sys_tmp148 = w_ip_FixedToFloat_floating_0;
	assign w_sys_tmp150 = (w_sys_tmp151 + r_run_j_8);
	assign w_sys_tmp151 = (w_sys_tmp140 * r_run_j_8);
	assign w_sys_tmp154 = (w_sys_tmp139 + r_run_i_7);
	assign w_sys_tmp163 = w_ip_AddFloat_result_0;
	assign w_sys_tmp164 = 32'h3f800000;
	assign w_sys_tmp165 = w_ip_MultFloat_product_0;
	assign w_sys_tmp166 = w_ip_DivFloat_quotient_0;
	assign w_sys_tmp167 = w_ip_MultFloat_product_0;
	assign w_sys_tmp168 = 32'h3f000000;
	assign w_sys_tmp169 = w_ip_AddFloat_result_0;
	assign w_sys_tmp170 = 32'h3f000000;
	assign w_sys_tmp171 = 32'h0;
	assign w_sys_tmp172 = w_ip_AddFloat_result_0;
	assign w_sys_tmp173 = 32'h3f000000;
	assign w_sys_tmp174 = 32'h0;
	assign w_sys_tmp175 = (r_run_k_9 < r_run_n_10);
	assign w_sys_tmp177 = w_ip_AddFloat_result_0;
	assign w_sys_tmp178 = w_fld_a_0_dataout_1;
	assign w_sys_tmp179 = (w_sys_tmp180 + r_run_k_9);
	assign w_sys_tmp180 = (w_sys_tmp181 * r_run_i_7);
	assign w_sys_tmp181 = 32'sh00000003;
	assign w_sys_tmp182 = w_ip_MultFloat_product_0;
	assign w_sys_tmp184 = (w_sys_tmp185 + r_run_k_9);
	assign w_sys_tmp185 = (w_sys_tmp181 * r_run_j_8);
	assign w_sys_tmp189 = 32'hbf800000;
	assign w_sys_tmp201 = w_sys_tmp177;
	assign w_sys_tmp207 = (r_run_k_9 + w_sys_intOne);
	assign w_sys_tmp208 = (r_run_k_9 < r_run_n_10);
	assign w_sys_tmp210 = w_ip_AddFloat_result_0;
	assign w_sys_tmp211 = w_fld_a_0_dataout_1;
	assign w_sys_tmp212 = (w_sys_tmp213 + r_run_i_7);
	assign w_sys_tmp213 = (w_sys_tmp214 * r_run_k_9);
	assign w_sys_tmp214 = 32'sh00000003;
	assign w_sys_tmp215 = w_ip_MultFloat_product_0;
	assign w_sys_tmp216 = (w_sys_tmp213 + r_run_j_8);
	assign w_sys_tmp220 = 32'hbf800000;
	assign w_sys_tmp232 = w_sys_tmp210;
	assign w_sys_tmp247 = ( -r_run_s_17 );
	assign w_sys_tmp265 = (r_run_k_9 + w_sys_intOne);
	assign w_sys_tmp266 = w_fld_a_0_dataout_1;


	DualPortRAM #(.DWIDTH(32), .AWIDTH(4), .WORDS(9) )
		dpram_a_0(
			.clk (clock),
			.ce_0 (w_fld_a_0_ce_0),
			.addr_0 (w_fld_a_0_addr_0),
			.datain_0 (w_fld_a_0_datain_0),
			.dataout_0 (w_fld_a_0_dataout_0),
			.r_w_0 (w_fld_a_0_r_w_0),
			.ce_1 (w_fld_a_0_ce_1),
			.addr_1 (r_fld_a_0_addr_1),
			.datain_1 (r_fld_a_0_datain_1),
			.dataout_1 (w_fld_a_0_dataout_1),
			.r_w_1 (r_fld_a_0_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(4), .WORDS(9) )
		dpram_x_1(
			.clk (clock),
			.ce_0 (w_fld_x_1_ce_0),
			.addr_0 (w_fld_x_1_addr_0),
			.datain_0 (w_fld_x_1_datain_0),
			.dataout_0 (w_fld_x_1_dataout_0),
			.r_w_0 (w_fld_x_1_r_w_0),
			.ce_1 (w_fld_x_1_ce_1),
			.addr_1 (r_fld_x_1_addr_1),
			.datain_1 (r_fld_x_1_datain_1),
			.dataout_1 (w_fld_x_1_dataout_1),
			.r_w_1 (r_fld_x_1_r_w_1)
		);

	AddFloat
		AddFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_AddFloat_portA_0),
			.b (r_ip_AddFloat_portB_0),
			.result (w_ip_AddFloat_result_0)
		);

	MultFloat
		MultFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_MultFloat_multiplicand_0),
			.b (r_ip_MultFloat_multiplier_0),
			.result (w_ip_MultFloat_product_0)
		);

	DivFloat
		DivFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_DivFloat_dividend_0),
			.b (r_ip_DivFloat_divisor_0),
			.result (w_ip_DivFloat_quotient_0)
		);

	CompareFloatLT
		CompareFloatLT_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_CompareFloatLT_portA_0),
			.b (r_ip_CompareFloatLT_portB_0),
			.result (w_ip_CompareFloatLT_result_0)
		);

	FixedToFloat
		FixedToFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_FixedToFloat_fixed_0),
			.result (w_ip_FixedToFloat_floating_0)
		);

	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_sqrt_phase) 
						4'h6: begin

							case(r_sys_sqrt_stage) 
								2'h0: begin
									if((r_sys_sqrt_step==7'h1e)) begin
										r_ip_AddFloat_portA_0 <= r_sqrt_x_5;

									end
								end

							endcase
						end

					endcase
				end

				3'h3: begin

					case(r_sys_run_phase) 
						7'h21: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_ip_AddFloat_portA_0 <= r_run_b2_12;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h5)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'hc)) begin
										r_ip_AddFloat_portA_0 <= r_run_b2_12;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h5)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp164;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp170;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp173;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8) || (r_sys_run_step==6'hb)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp0_float;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'he)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'hd)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp4_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_sqrt_phase) 
						4'h6: begin

							case(r_sys_sqrt_stage) 
								2'h0: begin
									if((r_sys_sqrt_step==7'h1e)) begin
										r_ip_AddFloat_portB_0 <= w_sys_tmp8;

									end
								end

							endcase
						end

					endcase
				end

				3'h3: begin

					case(r_sys_run_phase) 
						7'h21: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_ip_AddFloat_portB_0 <= w_sys_tmp101;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h5)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp137[31], w_sys_tmp137[30:0] };

									end
									else
									if((r_sys_run_step==6'hc)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp134[31], w_sys_tmp134[30:0] };

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h5)) begin
										r_ip_AddFloat_portB_0 <= w_sys_tmp165;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_ip_AddFloat_portB_0 <= r_run_coeff_15;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_ip_AddFloat_portB_0 <= { ~r_run_coeff_15[31], r_run_coeff_15[30:0] };

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8) || (r_sys_run_step==6'hb)) begin
										r_ip_AddFloat_portB_0 <= w_sys_tmp182;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he)) begin
										r_ip_AddFloat_portB_0 <= w_sys_tmp215;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h21: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp0_float;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp113;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp1_float;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h11)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp146;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h7)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp134;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h6)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp136;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_beta_14;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp168;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp189;

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp182;

									end
									else
									if((r_sys_run_step==6'h3)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_s_17;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h6)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_c_16;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h7)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp247;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp220;

									end
									else
									if((r_sys_run_step==6'h4) || (r_sys_run_step==6'h5)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_s_17;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h3) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h9)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_c_16;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h21: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp105;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp115;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_ip_MultFloat_multiplier_0 <= r_run_b2_12;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp129;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h7)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h6)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp137;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp148;

									end
									else
									if((r_sys_run_step==6'h11)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp147;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_ip_MultFloat_multiplier_0 <= r_run_beta_14;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_ip_MultFloat_multiplier_0 <= r_run_beta_14;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h3)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp178;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_ip_MultFloat_multiplier_0 <= r_run_s_17;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h5) || (r_sys_run_step==6'h9)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==6'h4) || (r_sys_run_step==6'h7)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp211;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_ip_MultFloat_multiplier_0 <= r_run_s_17;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_sqrt_phase) 
						4'h2: begin

							case(r_sys_sqrt_stage) 
								2'h0: begin
									if((r_sys_sqrt_step==7'h0)) begin
										r_ip_DivFloat_dividend_0 <= r_sqrt_s_4;

									end
								end

							endcase
						end

						4'h6: begin

							case(r_sys_sqrt_stage) 
								2'h0: begin
									if((r_sys_sqrt_step==7'h23)) begin
										r_ip_DivFloat_dividend_0 <= w_sys_tmp9;

									end
									else
									if((r_sys_sqrt_step==7'h0)) begin
										r_ip_DivFloat_dividend_0 <= r_sqrt_s_4;

									end
								end

							endcase
						end

					endcase
				end

				3'h3: begin

					case(r_sys_run_phase) 
						7'h26: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_ip_DivFloat_dividend_0 <= r_sys_tmp1_float;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'hb)) begin
										r_ip_DivFloat_dividend_0 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h16)) begin
										r_ip_DivFloat_dividend_0 <= w_sys_tmp134;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h5)) begin
										r_ip_DivFloat_dividend_0 <= w_sys_tmp167;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_sqrt_phase) 
						4'h2: begin

							case(r_sys_sqrt_stage) 
								2'h0: begin
									if((r_sys_sqrt_step==7'h0)) begin
										r_ip_DivFloat_divisor_0 <= w_sys_tmp5;

									end
								end

							endcase
						end

						4'h6: begin

							case(r_sys_sqrt_stage) 
								2'h0: begin
									if((r_sys_sqrt_step==7'h0)) begin
										r_ip_DivFloat_divisor_0 <= r_sqrt_x_5;

									end
									else
									if((r_sys_sqrt_step==7'h23)) begin
										r_ip_DivFloat_divisor_0 <= w_sys_tmp11;

									end
								end

							endcase
						end

					endcase
				end

				3'h3: begin

					case(r_sys_run_phase) 
						7'h26: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_ip_DivFloat_divisor_0 <= w_sys_tmp114;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h16)) begin
										r_ip_DivFloat_divisor_0 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'hb)) begin
										r_ip_DivFloat_divisor_0 <= w_sys_tmp134;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h5)) begin
										r_ip_DivFloat_divisor_0 <= r_run_tmp_20;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_max_phase) 
						4'h3: begin

							case(r_sys_max_stage) 
								2'h0: begin
									if((r_sys_max_step==3'h0)) begin
										r_ip_CompareFloatLT_portA_0 <= r_max_b_3;

									end
								end

							endcase
						end

					endcase
				end

				3'h3: begin

					case(r_sys_run_phase) 
						7'h23: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_ip_CompareFloatLT_portA_0 <= r_run_abserr_11;

									end
								end

							endcase
						end

						7'h28: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_ip_CompareFloatLT_portA_0 <= r_run_abserr_11;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_ip_CompareFloatLT_portA_0 <= r_run_bar_13;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_max_phase) 
						4'h3: begin

							case(r_sys_max_stage) 
								2'h0: begin
									if((r_sys_max_step==3'h0)) begin
										r_ip_CompareFloatLT_portB_0 <= r_max_a_2;

									end
								end

							endcase
						end

					endcase
				end

				3'h3: begin

					case(r_sys_run_phase) 
						7'h23: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_ip_CompareFloatLT_portB_0 <= r_run_b2_12;

									end
								end

							endcase
						end

						7'h28: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_ip_CompareFloatLT_portB_0 <= r_run_b2_12;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_ip_CompareFloatLT_portB_0 <= w_sys_tmp125;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h26: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1)) begin
										r_ip_FixedToFloat_fixed_0 <= r_run_n_10;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1)) begin
										r_ip_FixedToFloat_fixed_0 <= r_run_n_10;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 3'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 3'h3 : r_sys_processing_methodID);
				end

				3'h1: begin

					case(r_sys_max_phase) 
						4'h9: begin
							r_sys_processing_methodID <= r_sys_max_caller;
						end

					endcase
				end

				3'h2: begin

					case(r_sys_sqrt_phase) 
						4'ha: begin
							r_sys_processing_methodID <= r_sys_sqrt_caller;
						end

					endcase
				end

				3'h3: begin

					case(r_sys_run_phase) 
						7'h37: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'ha)) begin
										r_sys_processing_methodID <= 3'h2;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h5)) begin
										r_sys_processing_methodID <= 3'h1;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_processing_methodID <= 3'h2;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h5)) begin
										r_sys_processing_methodID <= 3'h1;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_processing_methodID <= 3'h2;

									end
								end

							endcase
						end

						7'h47: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_max_return <= 32'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_max_phase) 
						4'h4: begin
							r_sys_max_return <= w_sys_tmp2;
						end

						4'h6: begin
							r_sys_max_return <= w_sys_tmp3;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_max_caller <= 3'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h37: begin

							case(r_sys_run_stage) 
								4'h3: begin
									if((r_sys_run_step==6'h5)) begin
										r_sys_max_caller <= r_sys_processing_methodID;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h5)) begin
										r_sys_max_caller <= r_sys_processing_methodID;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_max_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_max_phase <= 4'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_max_phase) 
						4'h0: begin
							r_sys_max_phase <= 4'h3;
						end

						4'h3: begin

							case(r_sys_max_stage) 
								2'h0: begin
									if((r_sys_max_step==3'h3)) begin
										r_sys_max_phase <= ((w_sys_tmp1) ? 4'h5 : 4'h7);

									end
								end

							endcase
						end

						4'h4: begin
							r_sys_max_phase <= 4'h9;
						end

						4'h5: begin

							case(r_sys_max_stage) 
								2'h0: begin
									if((r_sys_max_step==3'h0)) begin
										r_sys_max_phase <= 4'h4;

									end
								end

							endcase
						end

						4'h6: begin
							r_sys_max_phase <= 4'h9;
						end

						4'h7: begin

							case(r_sys_max_stage) 
								2'h0: begin
									if((r_sys_max_step==3'h0)) begin
										r_sys_max_phase <= 4'h6;

									end
								end

							endcase
						end

						4'h9: begin
							r_sys_max_phase <= 4'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_max_stage <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_max_phase) 
						4'h3: begin

							case(r_sys_max_stage) 
								2'h0: begin
									if((r_sys_max_step==3'h3)) begin
										r_sys_max_stage <= 2'h0;

									end
								end

							endcase
						end

						4'h5: begin

							case(r_sys_max_stage) 
								2'h0: begin
									if((r_sys_max_step==3'h0)) begin
										r_sys_max_stage <= 2'h0;

									end
								end

							endcase
						end

						4'h7: begin

							case(r_sys_max_stage) 
								2'h0: begin
									if((r_sys_max_step==3'h0)) begin
										r_sys_max_stage <= 2'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_max_step <= 3'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_max_phase) 
						4'h3: begin

							case(r_sys_max_stage) 
								2'h0: begin
									if((r_sys_max_step==3'h3)) begin
										r_sys_max_step <= 3'h0;

									end
									else
									if((r_sys_max_step==3'h0) || (r_sys_max_step==3'h1) || (r_sys_max_step==3'h2)) begin
										r_sys_max_step <= w_sys_max_step_p1;

									end
								end

							endcase
						end

						4'h5: begin

							case(r_sys_max_stage) 
								2'h0: begin
									if((r_sys_max_step==3'h0)) begin
										r_sys_max_step <= 3'h0;

									end
								end

							endcase
						end

						4'h7: begin

							case(r_sys_max_stage) 
								2'h0: begin
									if((r_sys_max_step==3'h0)) begin
										r_sys_max_step <= 3'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_max_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_max_phase) 
						4'h0: begin
							r_sys_max_busy <= w_sys_boolTrue;
						end

						4'h9: begin
							r_sys_max_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_sqrt_return <= 32'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_sqrt_phase) 
						4'h7: begin
							r_sys_sqrt_return <= w_sys_tmp12;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_sqrt_caller <= 3'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h37: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'ha)) begin
										r_sys_sqrt_caller <= r_sys_processing_methodID;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_sqrt_caller <= r_sys_processing_methodID;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_sqrt_caller <= r_sys_processing_methodID;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_sqrt_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_sqrt_phase <= 4'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_sqrt_phase) 
						4'h0: begin
							r_sys_sqrt_phase <= 4'h2;
						end

						4'h2: begin

							case(r_sys_sqrt_stage) 
								2'h0: begin
									if((r_sys_sqrt_step==7'h1e)) begin
										r_sys_sqrt_phase <= 4'h4;

									end
								end

							endcase
						end

						4'h4: begin

							case(r_sys_sqrt_stage) 
								2'h0: begin
									if((r_sys_sqrt_step==7'h0)) begin
										r_sys_sqrt_phase <= ((w_sys_tmp7) ? 4'h6 : 4'h8);

									end
								end

							endcase
						end

						4'h6: begin

							case(r_sys_sqrt_stage) 
								2'h0: begin
									if((r_sys_sqrt_step==7'h41)) begin
										r_sys_sqrt_phase <= 4'h4;

									end
								end

							endcase
						end

						4'h7: begin
							r_sys_sqrt_phase <= 4'ha;
						end

						4'h8: begin

							case(r_sys_sqrt_stage) 
								2'h0: begin
									if((r_sys_sqrt_step==7'h0)) begin
										r_sys_sqrt_phase <= 4'h7;

									end
								end

							endcase
						end

						4'ha: begin
							r_sys_sqrt_phase <= 4'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_sqrt_stage <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_sqrt_phase) 
						4'h2: begin

							case(r_sys_sqrt_stage) 
								2'h0: begin
									if((r_sys_sqrt_step==7'h1e)) begin
										r_sys_sqrt_stage <= 2'h0;

									end
								end

							endcase
						end

						4'h4: begin

							case(r_sys_sqrt_stage) 
								2'h0: begin
									if((r_sys_sqrt_step==7'h0)) begin
										r_sys_sqrt_stage <= 2'h0;

									end
								end

							endcase
						end

						4'h6: begin

							case(r_sys_sqrt_stage) 
								2'h0: begin
									if((r_sys_sqrt_step==7'h41)) begin
										r_sys_sqrt_stage <= 2'h0;

									end
								end

							endcase
						end

						4'h8: begin

							case(r_sys_sqrt_stage) 
								2'h0: begin
									if((r_sys_sqrt_step==7'h0)) begin
										r_sys_sqrt_stage <= 2'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_sqrt_step <= 7'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_sqrt_phase) 
						4'h2: begin

							case(r_sys_sqrt_stage) 
								2'h0: begin
									if((7'h0<=r_sys_sqrt_step && r_sys_sqrt_step<=7'h1d)) begin
										r_sys_sqrt_step <= w_sys_sqrt_step_p1;

									end
									else
									if((r_sys_sqrt_step==7'h1e)) begin
										r_sys_sqrt_step <= 7'h0;

									end
								end

							endcase
						end

						4'h4: begin

							case(r_sys_sqrt_stage) 
								2'h0: begin
									if((r_sys_sqrt_step==7'h0)) begin
										r_sys_sqrt_step <= 7'h0;

									end
								end

							endcase
						end

						4'h6: begin

							case(r_sys_sqrt_stage) 
								2'h0: begin
									if((7'h0<=r_sys_sqrt_step && r_sys_sqrt_step<=7'h40)) begin
										r_sys_sqrt_step <= w_sys_sqrt_step_p1;

									end
									else
									if((r_sys_sqrt_step==7'h41)) begin
										r_sys_sqrt_step <= 7'h0;

									end
								end

							endcase
						end

						4'h8: begin

							case(r_sys_sqrt_stage) 
								2'h0: begin
									if((r_sys_sqrt_step==7'h0)) begin
										r_sys_sqrt_step <= 7'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_sqrt_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_sqrt_phase) 
						4'h0: begin
							r_sys_sqrt_busy <= w_sys_boolTrue;
						end

						4'ha: begin
							r_sys_sqrt_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_return <= 32'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h24: begin
							r_sys_run_return <= w_sys_tmp111;
						end

						7'h44: begin
							r_sys_run_return <= r_sys_tmp2_float;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 3'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 7'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h0: begin
							r_sys_run_phase <= 7'h2;
						end

						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 7'h4;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h5;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp41) ? 7'h9 : 7'hf);

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h5;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'ha;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp43) ? 7'hd : 7'h6);

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sys_run_phase <= 7'ha;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h10;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp87) ? 7'h13 : 7'h15);

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h10;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h16;

									end
								end

							endcase
						end

						7'h16: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp95) ? 7'h1a : 7'h23);

									end
								end

							endcase
						end

						7'h17: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h16;

									end
								end

							endcase
						end

						7'h1a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h1b;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp97) ? 7'h1f : 7'h17);

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h1b;

									end
								end

							endcase
						end

						7'h1f: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp99) ? 7'h21 : 7'h1c);

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_phase <= 7'h1c;

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_run_phase <= ((w_sys_tmp109) ? 7'h25 : 7'h26);

									end
								end

							endcase
						end

						7'h24: begin
							r_sys_run_phase <= 7'h47;
						end

						7'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h24;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2b)) begin
										r_sys_run_phase <= 7'h28;

									end
								end

							endcase
						end

						7'h28: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_run_phase <= ((w_sys_tmp116) ? 7'h2b : 7'h45);

									end
								end

							endcase
						end

						7'h2b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h2c;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp117) ? 7'h30 : 7'h28);

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h2c;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h31;

									end
								end

							endcase
						end

						7'h31: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp121) ? 7'h35 : 7'h2d);

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h31;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'hb)) begin
										r_sys_run_phase <= ((w_sys_tmp123) ? 7'h36 : 7'h37);

									end
								end

							endcase
						end

						7'h36: begin
							r_sys_run_phase <= 7'h32;
						end

						7'h37: begin

							case(r_sys_run_stage) 
								4'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_phase <= 7'h39;

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h3a;

									end
								end

							endcase
						end

						7'h3a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp175) ? 7'h3d : 7'h3f);

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h10)) begin
										r_sys_run_phase <= 7'h3a;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h40;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp208) ? 7'h43 : 7'h32);

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h13)) begin
										r_sys_run_phase <= 7'h40;

									end
								end

							endcase
						end

						7'h44: begin
							r_sys_run_phase <= 7'h47;
						end

						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_run_phase <= 7'h44;

									end
								end

							endcase
						end

						7'h47: begin
							r_sys_run_phase <= 7'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 4'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h16: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h17: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h1a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h1f: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2b)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h28: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h2b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h31: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'hb)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h34)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'hb)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h23)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h6)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h6)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h3a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h10)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h13)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 6'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h5)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h16: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h17: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h1a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h1f: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'hc)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h3)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h2a)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h2b)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h28: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h3)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h2b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h31: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'hb)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'ha)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h34)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h33)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								4'h1: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'ha)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'hb)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								4'h2: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h22)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h23)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								4'h3: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h5)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								4'h5: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h5)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h3a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'hf)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h10)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h12)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h13)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				3'h3: begin

					case(r_sys_run_phase) 
						7'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						7'h47: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_a_0_addr_1 <= 4'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp21[3:0] );

									end
									else
									if((r_sys_run_step==6'h4)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp27[3:0] );

									end
									else
									if((r_sys_run_step==6'h7)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp36[3:0] );

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp30[3:0] );

									end
									else
									if((r_sys_run_step==6'h3)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp13[3:0] );

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_intOne[3:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_intZero[3:0] );

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp39[3:0] );

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp33[3:0] );

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp102[3:0] );

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp126[3:0] );

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp154[3:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h4)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp138[3:0] );

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp150[3:0] );

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h2) || (r_sys_run_step==6'hd)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp179[3:0] );

									end
									else
									if((r_sys_run_step==6'h1) || (r_sys_run_step==6'h3) || (r_sys_run_step==6'h10)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp184[3:0] );

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h1) || (r_sys_run_step==6'h3) || (r_sys_run_step==6'h12)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp216[3:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h2) || (r_sys_run_step==6'he)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_tmp212[3:0] );

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_fld_a_0_addr_1 <= $signed( w_sys_intZero[3:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_fld_a_0_datain_1 <= w_sys_tmp17;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h7)) begin
										r_fld_a_0_datain_1 <= w_sys_tmp31;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h6)) begin
										r_fld_a_0_datain_1 <= w_sys_tmp22;

									end
									else
									if((r_sys_run_step==6'h1) || (r_sys_run_step==6'h3) || (r_sys_run_step==6'h4)) begin
										r_fld_a_0_datain_1 <= w_sys_tmp19;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_fld_a_0_datain_1 <= w_sys_tmp40;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h10)) begin
										r_fld_a_0_datain_1 <= w_sys_tmp201;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h12)) begin
										r_fld_a_0_datain_1 <= w_sys_tmp232;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_a_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_max_phase) 
						4'h9: begin
							r_fld_a_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

				3'h2: begin

					case(r_sys_sqrt_phase) 
						4'ha: begin
							r_fld_a_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

				3'h3: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_a_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1)) begin
										r_fld_a_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1)) begin
										r_fld_a_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h4)) begin
										r_fld_a_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3)) begin
										r_fld_a_0_r_w_1 <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h10)) begin
										r_fld_a_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3)) begin
										r_fld_a_0_r_w_1 <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h12)) begin
										r_fld_a_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_fld_a_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h47: begin
							r_fld_a_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_x_1_addr_1 <= 4'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_x_1_addr_1 <= $signed( w_sys_tmp46[3:0] );

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_fld_x_1_addr_1 <= $signed( w_sys_tmp90[3:0] );

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h1) || (r_sys_run_step==6'h3) || (r_sys_run_step==6'h13)) begin
										r_fld_x_1_addr_1 <= $signed( w_sys_tmp216[3:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h2) || (r_sys_run_step==6'hf)) begin
										r_fld_x_1_addr_1 <= $signed( w_sys_tmp212[3:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_x_1_datain_1 <= w_sys_tmp49;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_fld_x_1_datain_1 <= w_sys_tmp93;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'hf) || (r_sys_run_step==6'h13)) begin
										r_fld_x_1_datain_1 <= w_sys_tmp232;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_x_1_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_max_phase) 
						4'h9: begin
							r_fld_x_1_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

				3'h2: begin

					case(r_sys_sqrt_phase) 
						4'ha: begin
							r_fld_x_1_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

				3'h3: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_x_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_fld_x_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3)) begin
										r_fld_x_1_r_w_1 <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hf) || (r_sys_run_step==6'h13)) begin
										r_fld_x_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h47: begin
							r_fld_x_1_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h37: begin

							case(r_sys_run_stage) 
								4'h3: begin
									if((r_sys_run_step==6'h5)) begin
										r_max_a_2 <= w_sys_tmp169;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h5)) begin
										r_max_a_2 <= w_sys_tmp172;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h37: begin

							case(r_sys_run_stage) 
								4'h3: begin
									if((r_sys_run_step==6'h5)) begin
										r_max_b_3 <= w_sys_tmp171;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h5)) begin
										r_max_b_3 <= w_sys_tmp174;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h37: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'ha)) begin
										r_sqrt_s_4 <= w_sys_tmp163;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sqrt_s_4 <= r_run_tmp_20;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sqrt_s_4 <= r_run_tmp_20;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_sqrt_phase) 
						4'h2: begin

							case(r_sys_sqrt_stage) 
								2'h0: begin
									if((r_sys_sqrt_step==7'h1e)) begin
										r_sqrt_x_5 <= w_sys_tmp4;

									end
								end

							endcase
						end

						4'h6: begin

							case(r_sys_sqrt_stage) 
								2'h0: begin
									if((r_sys_sqrt_step==7'h41)) begin
										r_sqrt_x_5 <= w_sys_tmp8;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_sqrt_phase) 
						4'h2: begin

							case(r_sys_sqrt_stage) 
								2'h0: begin
									if((r_sys_sqrt_step==7'h0)) begin
										r_sqrt_last_x_6 <= w_sys_tmp6;

									end
								end

							endcase
						end

						4'h6: begin

							case(r_sys_sqrt_stage) 
								2'h0: begin
									if((r_sys_sqrt_step==7'h0)) begin
										r_sqrt_last_x_6 <= r_sqrt_x_5;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h4: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_i_7 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_i_7 <= w_sys_tmp42;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_i_7 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_i_7 <= w_sys_tmp94;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_i_7 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h17: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_i_7 <= w_sys_tmp96;

									end
								end

							endcase
						end

						7'h2b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_i_7 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_i_7 <= w_sys_tmp119;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_8 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_8 <= w_sys_tmp50;

									end
								end

							endcase
						end

						7'h1a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_8 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_8 <= w_sys_tmp98;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_8 <= w_sys_tmp120;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_8 <= w_sys_tmp122;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h39: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_9 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h10)) begin
										r_run_k_9 <= w_sys_tmp207;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_9 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h13)) begin
										r_run_k_9 <= w_sys_tmp265;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_n_10 <= w_sys_tmp13;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_abserr_11 <= w_sys_tmp14;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_b2_12 <= w_sys_tmp15;

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_run_b2_12 <= w_sys_tmp100;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h11)) begin
										r_run_b2_12 <= w_sys_tmp133;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h26: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2b)) begin
										r_run_bar_13 <= w_sys_tmp112;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h34)) begin
										r_run_bar_13 <= w_sys_tmp144;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h37: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h29)) begin
										r_run_beta_14 <= w_sys_tmp144;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h37: begin

							case(r_sys_run_stage) 
								4'h2: begin
									if((r_sys_run_step==6'h23)) begin
										r_run_coeff_15 <= w_sys_tmp166;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h37: begin

							case(r_sys_run_stage) 
								4'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_run_c_16 <= r_sys_sqrt_return;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h37: begin

							case(r_sys_run_stage) 
								4'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_run_s_17 <= r_sys_sqrt_return;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_run_cs_18 <= w_sys_tmp177;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'hf)) begin
										r_run_cs_18 <= w_sys_tmp210;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h10)) begin
										r_run_sc_19 <= w_sys_tmp177;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h12) || (r_sys_run_step==6'h13)) begin
										r_run_sc_19 <= w_sys_tmp210;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h37: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'hb)) begin
										r_run_tmp_20 <= r_sys_sqrt_return;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h6)) begin
										r_run_tmp_20 <= r_sys_max_return;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h6)) begin
										r_run_tmp_20 <= r_sys_max_return;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h21: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_fld_a_0_dataout_1;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h7)) begin
										r_sys_tmp0_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp0_float <= w_fld_a_0_dataout_1;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h4) || (r_sys_run_step==6'h5)) begin
										r_sys_tmp0_float <= w_fld_a_0_dataout_1;

									end
									else
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'ha)) begin
										r_sys_tmp0_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h4)) begin
										r_sys_tmp0_float <= w_fld_x_1_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h26: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h5)) begin
										r_sys_tmp1_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_fld_a_0_dataout_1;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h7)) begin
										r_sys_tmp1_float <= w_ip_FixedToFloat_floating_0;

									end
									else
									if((r_sys_run_step==6'h4)) begin
										r_sys_tmp1_float <= w_fld_a_0_dataout_1;

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_sys_tmp1_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_sys_tmp1_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h5)) begin
										r_sys_tmp1_float <= w_fld_a_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h43: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'hb)) begin
										r_sys_tmp2_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp2_float <= w_sys_tmp266;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h43: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h3) || (r_sys_run_step==6'h5)) begin
										r_sys_tmp3_float <= w_fld_x_1_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_run_phase) 
						7'h43: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h4)) begin
										r_sys_tmp4_float <= w_fld_a_0_dataout_1;

									end
									else
									if((r_sys_run_step==6'h8) || (r_sys_run_step==6'hc)) begin
										r_sys_tmp4_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
