/*
TimeStamp:	2016/9/5		15:35
*/


module c1_test(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy	
);

	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 6:0] r_sys_run_phase;
	reg         [ 1:0] r_sys_run_stage;
	reg         [ 6:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 1:0] w_sys_run_stage_p1;
	wire        [ 6:0] w_sys_run_step_p1;
	wire signed [14:0] w_fld_u_0_addr_0;
	wire        [31:0] w_fld_u_0_datain_0;
	wire        [31:0] w_fld_u_0_dataout_0;
	wire               w_fld_u_0_r_w_0;
	wire               w_fld_u_0_ce_0;
	reg  signed [14:0] r_fld_u_0_addr_1;
	reg         [31:0] r_fld_u_0_datain_1;
	wire        [31:0] w_fld_u_0_dataout_1;
	reg                r_fld_u_0_r_w_1;
	wire               w_fld_u_0_ce_1;
	wire signed [14:0] w_fld_uu_1_addr_0;
	wire        [31:0] w_fld_uu_1_datain_0;
	wire        [31:0] w_fld_uu_1_dataout_0;
	wire               w_fld_uu_1_r_w_0;
	wire               w_fld_uu_1_ce_0;
	reg  signed [14:0] r_fld_uu_1_addr_1;
	reg         [31:0] r_fld_uu_1_datain_1;
	wire        [31:0] w_fld_uu_1_dataout_1;
	reg                r_fld_uu_1_r_w_1;
	wire               w_fld_uu_1_ce_1;
	wire signed [14:0] w_fld_q_2_addr_0;
	wire        [31:0] w_fld_q_2_datain_0;
	wire        [31:0] w_fld_q_2_dataout_0;
	wire               w_fld_q_2_r_w_0;
	wire               w_fld_q_2_ce_0;
	reg  signed [14:0] r_fld_q_2_addr_1;
	reg         [31:0] r_fld_q_2_datain_1;
	wire        [31:0] w_fld_q_2_dataout_1;
	reg                r_fld_q_2_r_w_1;
	wire               w_fld_q_2_ce_1;
	reg  signed [31:0] r_run_k_5;
	reg  signed [31:0] r_run_j_6;
	reg  signed [31:0] r_run_n_7;
	reg  signed [31:0] r_run_mx_8;
	reg  signed [31:0] r_run_my_9;
	reg  signed [31:0] r_run_nlast_10;
	reg         [31:0] r_run_dx_11;
	reg         [31:0] r_run_dy_12;
	reg         [31:0] r_run_r1_13;
	reg         [31:0] r_run_r2_14;
	reg         [31:0] r_run_dt_15;
	reg  signed [31:0] r_run_copy0_j_16;
	reg  signed [31:0] r_run_copy0_j_17;
	reg  signed [31:0] r_run_copy1_j_18;
	reg  signed [31:0] r_run_copy2_j_19;
	reg  signed [31:0] r_run_copy0_j_20;
	reg  signed [31:0] r_run_copy0_j_21;
	reg  signed [31:0] r_run_copy0_j_22;
	reg  signed [31:0] r_run_copy0_j_23;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [14:0] w_sub01_u_addr;
	reg  signed [14:0] r_sub01_u_addr;
	wire        [31:0] w_sub01_u_datain;
	reg         [31:0] r_sub01_u_datain;
	wire        [31:0] w_sub01_u_dataout;
	wire               w_sub01_u_r_w;
	reg                r_sub01_u_r_w;
	wire signed [14:0] w_sub01_q_addr;
	reg  signed [14:0] r_sub01_q_addr;
	wire        [31:0] w_sub01_q_datain;
	reg         [31:0] r_sub01_q_datain;
	wire        [31:0] w_sub01_q_dataout;
	wire               w_sub01_q_r_w;
	reg                r_sub01_q_r_w;
	wire signed [14:0] w_sub01_result_addr;
	reg  signed [14:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [14:0] w_sub00_u_addr;
	reg  signed [14:0] r_sub00_u_addr;
	wire        [31:0] w_sub00_u_datain;
	reg         [31:0] r_sub00_u_datain;
	wire        [31:0] w_sub00_u_dataout;
	wire               w_sub00_u_r_w;
	reg                r_sub00_u_r_w;
	wire signed [14:0] w_sub00_q_addr;
	reg  signed [14:0] r_sub00_q_addr;
	wire        [31:0] w_sub00_q_datain;
	reg         [31:0] r_sub00_q_datain;
	wire        [31:0] w_sub00_q_dataout;
	wire               w_sub00_q_r_w;
	reg                r_sub00_q_r_w;
	wire signed [14:0] w_sub00_result_addr;
	reg  signed [14:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	wire signed [31:0] w_sys_tmp1;
	wire        [31:0] w_sys_tmp3;
	wire        [31:0] w_sys_tmp5;
	wire        [31:0] w_sys_tmp6;
	wire               w_sys_tmp8;
	wire               w_sys_tmp9;
	wire signed [31:0] w_sys_tmp10;
	wire               w_sys_tmp11;
	wire               w_sys_tmp12;
	wire signed [31:0] w_sys_tmp15;
	wire signed [31:0] w_sys_tmp16;
	wire signed [31:0] w_sys_tmp17;
	wire        [31:0] w_sys_tmp18;
	wire signed [31:0] w_sys_tmp20;
	wire signed [31:0] w_sys_tmp21;
	wire signed [31:0] w_sys_tmp24;
	wire signed [31:0] w_sys_tmp25;
	wire               w_sys_tmp254;
	wire               w_sys_tmp255;
	wire signed [31:0] w_sys_tmp256;
	wire               w_sys_tmp257;
	wire               w_sys_tmp258;
	wire signed [31:0] w_sys_tmp261;
	wire signed [31:0] w_sys_tmp262;
	wire        [31:0] w_sys_tmp263;
	wire signed [31:0] w_sys_tmp265;
	wire signed [31:0] w_sys_tmp266;
	wire        [31:0] w_sys_tmp268;
	wire signed [31:0] w_sys_tmp270;
	wire signed [31:0] w_sys_tmp271;
	wire        [31:0] w_sys_tmp273;
	wire signed [31:0] w_sys_tmp275;
	wire signed [31:0] w_sys_tmp276;
	wire signed [31:0] w_sys_tmp279;
	wire signed [31:0] w_sys_tmp280;
	wire signed [31:0] w_sys_tmp281;
	wire signed [31:0] w_sys_tmp282;
	wire               w_sys_tmp720;
	wire               w_sys_tmp721;
	wire signed [31:0] w_sys_tmp722;
	wire signed [31:0] w_sys_tmp723;
	wire               w_sys_tmp724;
	wire               w_sys_tmp725;
	wire signed [31:0] w_sys_tmp726;
	wire signed [31:0] w_sys_tmp729;
	wire signed [31:0] w_sys_tmp730;
	wire signed [31:0] w_sys_tmp731;
	wire        [31:0] w_sys_tmp732;
	wire signed [31:0] w_sys_tmp733;
	wire signed [31:0] w_sys_tmp734;
	wire signed [31:0] w_sys_tmp736;
	wire signed [31:0] w_sys_tmp737;
	wire signed [31:0] w_sys_tmp928;
	wire               w_sys_tmp929;
	wire               w_sys_tmp930;
	wire signed [31:0] w_sys_tmp931;
	wire signed [31:0] w_sys_tmp932;
	wire               w_sys_tmp933;
	wire               w_sys_tmp934;
	wire signed [31:0] w_sys_tmp935;
	wire signed [31:0] w_sys_tmp938;
	wire signed [31:0] w_sys_tmp939;
	wire signed [31:0] w_sys_tmp940;
	wire        [31:0] w_sys_tmp941;
	wire signed [31:0] w_sys_tmp942;
	wire signed [31:0] w_sys_tmp943;
	wire signed [31:0] w_sys_tmp945;
	wire signed [31:0] w_sys_tmp946;
	wire signed [31:0] w_sys_tmp1137;
	wire               w_sys_tmp1138;
	wire               w_sys_tmp1139;
	wire signed [31:0] w_sys_tmp1140;
	wire signed [31:0] w_sys_tmp1141;
	wire signed [31:0] w_sys_tmp1142;
	wire               w_sys_tmp1143;
	wire               w_sys_tmp1144;
	wire signed [31:0] w_sys_tmp1145;
	wire signed [31:0] w_sys_tmp1148;
	wire signed [31:0] w_sys_tmp1149;
	wire signed [31:0] w_sys_tmp1150;
	wire        [31:0] w_sys_tmp1151;
	wire signed [31:0] w_sys_tmp1152;
	wire signed [31:0] w_sys_tmp1153;
	wire signed [31:0] w_sys_tmp1155;
	wire signed [31:0] w_sys_tmp1156;
	wire signed [31:0] w_sys_tmp1347;
	wire               w_sys_tmp1348;
	wire               w_sys_tmp1349;
	wire signed [31:0] w_sys_tmp1350;
	wire signed [31:0] w_sys_tmp1351;
	wire signed [31:0] w_sys_tmp1352;
	wire               w_sys_tmp1353;
	wire               w_sys_tmp1354;
	wire signed [31:0] w_sys_tmp1355;
	wire signed [31:0] w_sys_tmp1358;
	wire signed [31:0] w_sys_tmp1359;
	wire signed [31:0] w_sys_tmp1360;
	wire        [31:0] w_sys_tmp1361;
	wire signed [31:0] w_sys_tmp1362;
	wire signed [31:0] w_sys_tmp1363;
	wire signed [31:0] w_sys_tmp1365;
	wire signed [31:0] w_sys_tmp1366;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 2'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 7'h1);
	assign w_fld_u_0_addr_0 = 15'sh0;
	assign w_fld_u_0_datain_0 = 32'h0;
	assign w_fld_u_0_r_w_0 = 1'h0;
	assign w_fld_u_0_ce_0 = w_sys_ce;
	assign w_fld_u_0_ce_1 = w_sys_ce;
	assign w_fld_uu_1_addr_0 = 15'sh0;
	assign w_fld_uu_1_datain_0 = 32'h0;
	assign w_fld_uu_1_r_w_0 = 1'h0;
	assign w_fld_uu_1_ce_0 = w_sys_ce;
	assign w_fld_uu_1_ce_1 = w_sys_ce;
	assign w_fld_q_2_addr_0 = 15'sh0;
	assign w_fld_q_2_datain_0 = 32'h0;
	assign w_fld_q_2_r_w_0 = 1'h0;
	assign w_fld_q_2_ce_0 = w_sys_ce;
	assign w_fld_q_2_ce_1 = w_sys_ce;
	assign w_sub01_u_addr = ( (|r_sys_processing_methodID) ? r_sub01_u_addr : 15'sh0 ) ;
	assign w_sub01_u_datain = ( (|r_sys_processing_methodID) ? r_sub01_u_datain : 32'h0 ) ;
	assign w_sub01_u_r_w = ( (|r_sys_processing_methodID) ? r_sub01_u_r_w : 1'h0 ) ;
	assign w_sub01_q_addr = ( (|r_sys_processing_methodID) ? r_sub01_q_addr : 15'sh0 ) ;
	assign w_sub01_q_datain = ( (|r_sys_processing_methodID) ? r_sub01_q_datain : 32'h0 ) ;
	assign w_sub01_q_r_w = ( (|r_sys_processing_methodID) ? r_sub01_q_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 15'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub00_u_addr = ( (|r_sys_processing_methodID) ? r_sub00_u_addr : 15'sh0 ) ;
	assign w_sub00_u_datain = ( (|r_sys_processing_methodID) ? r_sub00_u_datain : 32'h0 ) ;
	assign w_sub00_u_r_w = ( (|r_sys_processing_methodID) ? r_sub00_u_r_w : 1'h0 ) ;
	assign w_sub00_q_addr = ( (|r_sys_processing_methodID) ? r_sub00_q_addr : 15'sh0 ) ;
	assign w_sub00_q_datain = ( (|r_sys_processing_methodID) ? r_sub00_q_datain : 32'h0 ) ;
	assign w_sub00_q_r_w = ( (|r_sys_processing_methodID) ? r_sub00_q_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 15'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh00000081;
	assign w_sys_tmp3 = 32'h3c000000;
	assign w_sys_tmp5 = 32'h3ba3d70a;
	assign w_sys_tmp6 = 32'h42a3d70a;
	assign w_sys_tmp8 = ( !w_sys_tmp9 );
	assign w_sys_tmp9 = (r_run_my_9 < r_run_k_5);
	assign w_sys_tmp10 = (r_run_k_5 + w_sys_intOne);
	assign w_sys_tmp11 = ( !w_sys_tmp12 );
	assign w_sys_tmp12 = (r_run_mx_8 < r_run_j_6);
	assign w_sys_tmp15 = (w_sys_tmp16 + r_run_k_5);
	assign w_sys_tmp16 = (r_run_j_6 * w_sys_tmp17);
	assign w_sys_tmp17 = 32'sh00000081;
	assign w_sys_tmp18 = 32'h0;
	assign w_sys_tmp20 = (w_sys_tmp21 + r_run_k_5);
	assign w_sys_tmp21 = (r_run_copy0_j_16 * w_sys_tmp17);
	assign w_sys_tmp24 = (r_run_copy0_j_16 + w_sys_intOne);
	assign w_sys_tmp25 = (r_run_j_6 + w_sys_intOne);
	assign w_sys_tmp254 = ( !w_sys_tmp255 );
	assign w_sys_tmp255 = (r_run_nlast_10 < r_run_n_7);
	assign w_sys_tmp256 = (r_run_n_7 + w_sys_intOne);
	assign w_sys_tmp257 = ( !w_sys_tmp258 );
	assign w_sys_tmp258 = (r_run_my_9 < r_run_j_6);
	assign w_sys_tmp261 = (w_sys_tmp262 + r_run_j_6);
	assign w_sys_tmp262 = 32'sh00000081;
	assign w_sys_tmp263 = 32'h3f000000;
	assign w_sys_tmp265 = (w_sys_tmp266 + r_run_copy2_j_19);
	assign w_sys_tmp266 = (r_run_mx_8 * w_sys_tmp262);
	assign w_sys_tmp268 = 32'h0;
	assign w_sys_tmp270 = (w_sys_tmp271 + w_sys_intOne);
	assign w_sys_tmp271 = (r_run_copy1_j_18 * w_sys_tmp262);
	assign w_sys_tmp273 = 32'h3f800000;
	assign w_sys_tmp275 = (w_sys_tmp276 + r_run_my_9);
	assign w_sys_tmp276 = (r_run_copy0_j_17 * w_sys_tmp262);
	assign w_sys_tmp279 = (r_run_copy0_j_17 + w_sys_intOne);
	assign w_sys_tmp280 = (r_run_copy1_j_18 + w_sys_intOne);
	assign w_sys_tmp281 = (r_run_copy2_j_19 + w_sys_intOne);
	assign w_sys_tmp282 = (r_run_j_6 + w_sys_intOne);
	assign w_sys_tmp720 = ( !w_sys_tmp721 );
	assign w_sys_tmp721 = (w_sys_tmp722 < r_run_k_5);
	assign w_sys_tmp722 = 32'sh00000041;
	assign w_sys_tmp723 = (r_run_k_5 + w_sys_intOne);
	assign w_sys_tmp724 = ( !w_sys_tmp725 );
	assign w_sys_tmp725 = (w_sys_tmp726 < r_run_j_6);
	assign w_sys_tmp726 = 32'sh00000081;
	assign w_sys_tmp729 = (w_sys_tmp730 + r_run_k_5);
	assign w_sys_tmp730 = (r_run_j_6 * w_sys_tmp731);
	assign w_sys_tmp731 = 32'sh00000081;
	assign w_sys_tmp732 = w_fld_u_0_dataout_1;
	assign w_sys_tmp733 = (w_sys_tmp734 + r_run_k_5);
	assign w_sys_tmp734 = (r_run_copy0_j_20 * w_sys_tmp731);
	assign w_sys_tmp736 = (r_run_copy0_j_20 + w_sys_intOne);
	assign w_sys_tmp737 = (r_run_j_6 + w_sys_intOne);
	assign w_sys_tmp928 = 32'sh00000040;
	assign w_sys_tmp929 = ( !w_sys_tmp930 );
	assign w_sys_tmp930 = (w_sys_tmp931 < r_run_k_5);
	assign w_sys_tmp931 = 32'sh00000081;
	assign w_sys_tmp932 = (r_run_k_5 + w_sys_intOne);
	assign w_sys_tmp933 = ( !w_sys_tmp934 );
	assign w_sys_tmp934 = (w_sys_tmp935 < r_run_j_6);
	assign w_sys_tmp935 = 32'sh00000081;
	assign w_sys_tmp938 = (w_sys_tmp939 + r_run_k_5);
	assign w_sys_tmp939 = (r_run_j_6 * w_sys_tmp940);
	assign w_sys_tmp940 = 32'sh00000081;
	assign w_sys_tmp941 = w_fld_u_0_dataout_1;
	assign w_sys_tmp942 = (w_sys_tmp943 + r_run_k_5);
	assign w_sys_tmp943 = (r_run_copy0_j_21 * w_sys_tmp940);
	assign w_sys_tmp945 = (r_run_copy0_j_21 + w_sys_intOne);
	assign w_sys_tmp946 = (r_run_j_6 + w_sys_intOne);
	assign w_sys_tmp1137 = 32'sh00000002;
	assign w_sys_tmp1138 = ( !w_sys_tmp1139 );
	assign w_sys_tmp1139 = (w_sys_tmp1140 < r_run_k_5);
	assign w_sys_tmp1140 = 32'sh00000040;
	assign w_sys_tmp1141 = (r_run_k_5 + w_sys_intOne);
	assign w_sys_tmp1142 = 32'sh00000002;
	assign w_sys_tmp1143 = ( !w_sys_tmp1144 );
	assign w_sys_tmp1144 = (w_sys_tmp1145 < r_run_j_6);
	assign w_sys_tmp1145 = 32'sh00000080;
	assign w_sys_tmp1148 = (w_sys_tmp1149 + r_run_k_5);
	assign w_sys_tmp1149 = (r_run_j_6 * w_sys_tmp1150);
	assign w_sys_tmp1150 = 32'sh00000081;
	assign w_sys_tmp1151 = w_sub00_result_dataout;
	assign w_sys_tmp1152 = (w_sys_tmp1153 + r_run_k_5);
	assign w_sys_tmp1153 = (r_run_copy0_j_22 * w_sys_tmp1150);
	assign w_sys_tmp1155 = (r_run_copy0_j_22 + w_sys_intOne);
	assign w_sys_tmp1156 = (r_run_j_6 + w_sys_intOne);
	assign w_sys_tmp1347 = 32'sh00000041;
	assign w_sys_tmp1348 = ( !w_sys_tmp1349 );
	assign w_sys_tmp1349 = (w_sys_tmp1350 < r_run_k_5);
	assign w_sys_tmp1350 = 32'sh00000080;
	assign w_sys_tmp1351 = (r_run_k_5 + w_sys_intOne);
	assign w_sys_tmp1352 = 32'sh00000002;
	assign w_sys_tmp1353 = ( !w_sys_tmp1354 );
	assign w_sys_tmp1354 = (w_sys_tmp1355 < r_run_j_6);
	assign w_sys_tmp1355 = 32'sh00000080;
	assign w_sys_tmp1358 = (w_sys_tmp1359 + r_run_k_5);
	assign w_sys_tmp1359 = (r_run_j_6 * w_sys_tmp1360);
	assign w_sys_tmp1360 = 32'sh00000081;
	assign w_sys_tmp1361 = w_sub01_result_dataout;
	assign w_sys_tmp1362 = (w_sys_tmp1363 + r_run_k_5);
	assign w_sys_tmp1363 = (r_run_copy0_j_23 * w_sys_tmp1360);
	assign w_sys_tmp1365 = (r_run_copy0_j_23 + w_sys_intOne);
	assign w_sys_tmp1366 = (r_run_j_6 + w_sys_intOne);


	subunder
		sub01_inst(
			.i_fld_q_1_addr_0 (w_sub01_q_addr),
			.i_fld_q_1_datain_0 (w_sub01_q_datain),
			.o_fld_q_1_dataout_0 (w_sub01_q_dataout),
			.i_fld_q_1_r_w_0 (w_sub01_q_r_w),
			.i_fld_result_2_addr_0 (w_sub01_result_addr),
			.i_fld_result_2_datain_0 (w_sub01_result_datain),
			.o_fld_result_2_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub01_result_r_w),
			.i_fld_u_0_addr_0 (w_sub01_u_addr),
			.i_fld_u_0_datain_0 (w_sub01_u_datain),
			.o_fld_u_0_dataout_0 (w_sub01_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub01_u_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	subup
		sub00_inst(
			.i_fld_q_1_addr_0 (w_sub00_q_addr),
			.i_fld_q_1_datain_0 (w_sub00_q_datain),
			.o_fld_q_1_dataout_0 (w_sub00_q_dataout),
			.i_fld_q_1_r_w_0 (w_sub00_q_r_w),
			.i_fld_result_2_addr_0 (w_sub00_result_addr),
			.i_fld_result_2_datain_0 (w_sub00_result_datain),
			.o_fld_result_2_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub00_result_r_w),
			.i_fld_u_0_addr_0 (w_sub00_u_addr),
			.i_fld_u_0_datain_0 (w_sub00_u_datain),
			.o_fld_u_0_dataout_0 (w_sub00_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub00_u_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_u_0(
			.clk (clock),
			.ce_0 (w_fld_u_0_ce_0),
			.addr_0 (w_fld_u_0_addr_0),
			.datain_0 (w_fld_u_0_datain_0),
			.dataout_0 (w_fld_u_0_dataout_0),
			.r_w_0 (w_fld_u_0_r_w_0),
			.ce_1 (w_fld_u_0_ce_1),
			.addr_1 (r_fld_u_0_addr_1),
			.datain_1 (r_fld_u_0_datain_1),
			.dataout_1 (w_fld_u_0_dataout_1),
			.r_w_1 (r_fld_u_0_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_uu_1(
			.clk (clock),
			.ce_0 (w_fld_uu_1_ce_0),
			.addr_0 (w_fld_uu_1_addr_0),
			.datain_0 (w_fld_uu_1_datain_0),
			.dataout_0 (w_fld_uu_1_dataout_0),
			.r_w_0 (w_fld_uu_1_r_w_0),
			.ce_1 (w_fld_uu_1_ce_1),
			.addr_1 (r_fld_uu_1_addr_1),
			.datain_1 (r_fld_uu_1_datain_1),
			.dataout_1 (w_fld_uu_1_dataout_1),
			.r_w_1 (r_fld_uu_1_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_q_2(
			.clk (clock),
			.ce_0 (w_fld_q_2_ce_0),
			.addr_0 (w_fld_q_2_addr_0),
			.datain_0 (w_fld_q_2_datain_0),
			.dataout_0 (w_fld_q_2_dataout_0),
			.r_w_0 (w_fld_q_2_r_w_0),
			.ce_1 (w_fld_q_2_ce_1),
			.addr_1 (r_fld_q_2_addr_1),
			.datain_1 (r_fld_q_2_datain_1),
			.dataout_1 (w_fld_q_2_dataout_1),
			.r_w_1 (r_fld_q_2_r_w_1)
		);

	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						7'h49: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 7'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h0: begin
							r_sys_run_phase <= 7'h2;
						end

						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h4;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h5;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp8) ? 7'h9 : 7'hf);

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h5;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'ha;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp11) ? 7'hd : 7'h6);

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h13)) begin
										r_sys_run_phase <= 7'ha;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h10;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp254) ? 7'h14 : 7'h49);

									end
								end

							endcase
						end

						7'h11: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h10;

									end
								end

							endcase
						end

						7'h14: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h15;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp257) ? 7'h18 : 7'h1a);

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h4f)) begin
										r_sys_run_phase <= 7'h15;

									end
								end

							endcase
						end

						7'h1a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h1b;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp720) ? 7'h1f : 7'h25);

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h1b;

									end
								end

							endcase
						end

						7'h1f: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h20;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp724) ? 7'h23 : 7'h1c);

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h15)) begin
										r_sys_run_phase <= 7'h20;

									end
								end

							endcase
						end

						7'h25: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h26;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp929) ? 7'h2a : 7'h2f);

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h26;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h2b;

									end
								end

							endcase
						end

						7'h2b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp933) ? 7'h2e : 7'h27);

									end
								end

							endcase
						end

						7'h2e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h15)) begin
										r_sys_run_phase <= 7'h2b;

									end
								end

							endcase
						end

						7'h2f: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_phase <= 7'h31;

									end
								end

							endcase
						end

						7'h31: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_phase <= 7'h33;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h34;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1138) ? 7'h38 : 7'h3e);

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h34;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h39;

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1143) ? 7'h3c : 7'h35);

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h15)) begin
										r_sys_run_phase <= 7'h39;

									end
								end

							endcase
						end

						7'h3e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h3f;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1348) ? 7'h43 : 7'h11);

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h3f;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h44;

									end
								end

							endcase
						end

						7'h44: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1353) ? 7'h47 : 7'h40);

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h15)) begin
										r_sys_run_phase <= 7'h44;

									end
								end

							endcase
						end

						7'h49: begin
							r_sys_run_phase <= 7'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h13)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h11: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h14: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h4f)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h1a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h1f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h15)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h25: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h2b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h2e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h15)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h31: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h15)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h3e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h44: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h15)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 7'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h12)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h11: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h14: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h4e)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h4f)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h1a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h1f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h14)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h25: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h2b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h2e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h14)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h31: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub00_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub01_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h14)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h3e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h44: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h14)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						7'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						7'h49: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp15[14:0] );

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h4) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h38) || (r_sys_run_step==7'h3c) || (r_sys_run_step==7'h40) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h48) || (r_sys_run_step==7'h4c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp261[14:0] );

									end
									else
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h2b) || (r_sys_run_step==7'h2f) || (r_sys_run_step==7'h33) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h3b) || (r_sys_run_step==7'h3f) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h47) || (r_sys_run_step==7'h4b) || (r_sys_run_step==7'h4f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp275[14:0] );

									end
									else
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h3e) || (r_sys_run_step==7'h42) || (r_sys_run_step==7'h46) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h4e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp270[14:0] );

									end
									else
									if((r_sys_run_step==7'h1) || (r_sys_run_step==7'h5) || (r_sys_run_step==7'h9) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h45) || (r_sys_run_step==7'h49) || (r_sys_run_step==7'h4d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp265[14:0] );

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp733[14:0] );

									end
								end

							endcase
						end

						7'h2e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp942[14:0] );

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h15)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1148[14:0] );

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h15)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1358[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp18;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1) || (r_sys_run_step==7'h3) || (r_sys_run_step==7'h5) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'h9) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h2b) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h2f) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h33) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h3b) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h3f) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h45) || (r_sys_run_step==7'h47) || (r_sys_run_step==7'h49) || (r_sys_run_step==7'h4b) || (r_sys_run_step==7'h4d) || (r_sys_run_step==7'h4f)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp268;

									end
									else
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h3e) || (r_sys_run_step==7'h42) || (r_sys_run_step==7'h46) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h4e)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp273;

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h4) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h38) || (r_sys_run_step==7'h3c) || (r_sys_run_step==7'h40) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h48) || (r_sys_run_step==7'h4c)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp263;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h15)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp1151;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h15)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp1361;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h4f)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h2e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h15)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h15)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h49: begin
							r_fld_u_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_uu_1_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_fld_uu_1_addr_1 <= $signed( w_sys_tmp20[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_fld_uu_1_datain_1 <= w_sys_tmp18;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_uu_1_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_fld_uu_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h49: begin
							r_fld_uu_1_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_q_2_addr_1 <= 15'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_q_2_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h49: begin
							r_fld_q_2_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_5 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_5 <= w_sys_tmp10;

									end
								end

							endcase
						end

						7'h1a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_5 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_5 <= w_sys_tmp723;

									end
								end

							endcase
						end

						7'h25: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_5 <= w_sys_tmp928;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_5 <= w_sys_tmp932;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_5 <= w_sys_tmp1137;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_5 <= w_sys_tmp1141;

									end
								end

							endcase
						end

						7'h3e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_5 <= w_sys_tmp1347;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_5 <= w_sys_tmp1351;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_6 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_run_j_6 <= w_sys_tmp25;

									end
								end

							endcase
						end

						7'h14: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_6 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h4) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h38) || (r_sys_run_step==7'h3c) || (r_sys_run_step==7'h40) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h48) || (r_sys_run_step==7'h4c)) begin
										r_run_j_6 <= w_sys_tmp282;

									end
								end

							endcase
						end

						7'h1f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_6 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h15)) begin
										r_run_j_6 <= w_sys_tmp737;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_6 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h2e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h15)) begin
										r_run_j_6 <= w_sys_tmp946;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_6 <= w_sys_tmp1142;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h15)) begin
										r_run_j_6 <= w_sys_tmp1156;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_6 <= w_sys_tmp1352;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h15)) begin
										r_run_j_6 <= w_sys_tmp1366;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hf: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_n_7 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h11: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_n_7 <= w_sys_tmp256;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_mx_8 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_my_9 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_nlast_10 <= w_sys_intOne;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_dx_11 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_dy_12 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_r1_13 <= w_sys_tmp6;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_r2_14 <= w_sys_tmp6;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_dt_15 <= w_sys_tmp5;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_16 <= r_run_j_6;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_run_copy0_j_16 <= w_sys_tmp24;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h14: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_17 <= r_run_j_6;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h2b) || (r_sys_run_step==7'h2f) || (r_sys_run_step==7'h33) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h3b) || (r_sys_run_step==7'h3f) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h47) || (r_sys_run_step==7'h4b) || (r_sys_run_step==7'h4f)) begin
										r_run_copy0_j_17 <= w_sys_tmp279;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h14: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_18 <= r_run_j_6;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h3e) || (r_sys_run_step==7'h42) || (r_sys_run_step==7'h46) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h4e)) begin
										r_run_copy1_j_18 <= w_sys_tmp280;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h14: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy2_j_19 <= r_run_j_6;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1) || (r_sys_run_step==7'h5) || (r_sys_run_step==7'h9) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h45) || (r_sys_run_step==7'h49) || (r_sys_run_step==7'h4d)) begin
										r_run_copy2_j_19 <= w_sys_tmp281;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h1f: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_20 <= r_run_j_6;

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_run_copy0_j_20 <= w_sys_tmp736;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2a: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_21 <= r_run_j_6;

									end
								end

							endcase
						end

						7'h2e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_run_copy0_j_21 <= w_sys_tmp945;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h38: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_22 <= r_run_j_6;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_run_copy0_j_22 <= w_sys_tmp1155;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h43: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_23 <= r_run_j_6;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_run_copy0_j_23 <= w_sys_tmp1365;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2f: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h15)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp938[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h15)) begin
										r_sub01_u_datain <= w_sys_tmp941;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h15)) begin
										r_sub01_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h49: begin
							r_sub01_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_q_addr <= 15'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_q_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_q_r_w <= w_sys_boolFalse;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_q_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h49: begin
							r_sub01_q_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h47: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1362[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h49: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h23: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h15)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp729[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h23: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h15)) begin
										r_sub00_u_datain <= w_sys_tmp732;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h23: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h15)) begin
										r_sub00_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h49: begin
							r_sub00_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_q_addr <= 15'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_q_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_q_r_w <= w_sys_boolFalse;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_q_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h49: begin
							r_sub00_q_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1152[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h13)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h49: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


endmodule
