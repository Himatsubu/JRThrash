/*
TimeStamp:	2017/1/5		15:28
*/


module TopClass(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_mainRoutine_req,	
	output                o_mainRoutine_busy,	
	output signed  [31:0] o_mainRoutine_return,	
	output signed  [31:0] o_mainRoutine_arrayY_4_addr,	
	output signed  [31:0] o_mainRoutine_arrayY_4_datain,	
	input  signed  [31:0] i_mainRoutine_arrayY_4_dataout,	
	output                o_mainRoutine_arrayY_4_r_w,	
	output                o_mainRoutine_arrayY_4_ce,	
	input                 i_mainRoutine_arrayY_4_cacheHit,	
	input  signed  [31:0] i_mainRoutine_dataNum_5	
);

	reg                r_sys_setValueToChildArray_arbiter0;
	reg                r_sys_subAprocess_arbiter1;
	reg                r_sys_subBprocess_arbiter2;
	reg                r_sys_subRoutine_arbiter3;
	reg  signed [31:0] r_ip_FixedToFloat_fixed_0;
	wire        [31:0] w_ip_FixedToFloat_floating_0;
	reg         [ 2:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [31:0] r_sys_mainRoutine_return;
	reg         [ 2:0] r_sys_mainRoutine_caller;
	reg                r_sys_mainRoutine_req;
	reg         [ 2:0] r_sys_mainRoutine_phase;
	reg         [ 2:0] r_sys_mainRoutine_stage;
	reg         [ 3:0] r_sys_mainRoutine_step;
	reg                r_sys_mainRoutine_busy;
	wire        [ 2:0] w_sys_mainRoutine_stage_p1;
	wire        [ 3:0] w_sys_mainRoutine_step_p1;
	reg  signed [31:0] r_sys_setValueToChildArray_return;
	reg         [ 2:0] r_sys_setValueToChildArray_caller;
	reg                r_sys_setValueToChildArray_req;
	reg         [ 3:0] r_sys_setValueToChildArray_phase;
	reg         [ 1:0] r_sys_setValueToChildArray_stage;
	reg         [ 2:0] r_sys_setValueToChildArray_step;
	reg                r_sys_setValueToChildArray_busy;
	wire        [ 1:0] w_sys_setValueToChildArray_stage_p1;
	wire        [ 2:0] w_sys_setValueToChildArray_step_p1;
	reg  signed [31:0] r_sys_subRoutine_return;
	reg         [ 2:0] r_sys_subRoutine_caller;
	reg                r_sys_subRoutine_req;
	reg         [ 4:0] r_sys_subRoutine_phase;
	reg         [ 1:0] r_sys_subRoutine_stage;
	reg         [ 2:0] r_sys_subRoutine_step;
	reg                r_sys_subRoutine_busy;
	wire        [ 1:0] w_sys_subRoutine_stage_p1;
	wire        [ 2:0] w_sys_subRoutine_step_p1;
	wire signed [ 4:0] w_fld_arrayX_3_addr_0;
	wire signed [31:0] w_fld_arrayX_3_datain_0;
	wire signed [31:0] w_fld_arrayX_3_dataout_0;
	wire               w_fld_arrayX_3_r_w_0;
	wire               w_fld_arrayX_3_ce_0;
	reg  signed [ 4:0] r_fld_arrayX_3_addr_1;
	reg  signed [31:0] r_fld_arrayX_3_datain_1;
	wire signed [31:0] w_fld_arrayX_3_dataout_1;
	reg                r_fld_arrayX_3_r_w_1;
	wire               w_fld_arrayX_3_ce_1;
	reg  signed [31:0] r_mainRoutine_arrayY_4_addr;
	reg  signed [31:0] r_mainRoutine_arrayY_4_datain;
	wire signed [31:0] w_mainRoutine_arrayY_4_dataout;
	reg                r_mainRoutine_arrayY_4_r_w;
	wire signed [31:0] w_mainRoutine_arrayY_4_addr;
	wire signed [31:0] w_mainRoutine_arrayY_4_datain;
	wire               w_mainRoutine_arrayY_4_r_w;
	wire               w_mainRoutine_arrayY_4_ce;
	wire               w_mainRoutine_arrayY_4_cacheHit;
	reg  signed [31:0] r_mainRoutine_dataNum_5;
	reg  signed [31:0] r_mainRoutine_subARet_6;
	reg  signed [31:0] r_mainRoutine_subBRet_7;
	reg  signed [31:0] r_mainRoutine_subXRet_8;
	reg  signed [31:0] r_setValueToChildArray_ax_9_addr;
	reg  signed [31:0] r_setValueToChildArray_ax_9_datain;
	wire signed [31:0] w_setValueToChildArray_ax_9_dataout;
	reg                r_setValueToChildArray_ax_9_r_w;
	wire signed [31:0] w_setValueToChildArray_ax_9_addr;
	wire signed [31:0] w_setValueToChildArray_ax_9_datain;
	wire               w_setValueToChildArray_ax_9_r_w;
	wire               w_setValueToChildArray_ax_9_ce;
	wire               w_setValueToChildArray_ax_9_cacheHit;
	reg  signed [31:0] r_setValueToChildArray_bx_10_addr;
	reg  signed [31:0] r_setValueToChildArray_bx_10_datain;
	wire signed [31:0] w_setValueToChildArray_bx_10_dataout;
	reg                r_setValueToChildArray_bx_10_r_w;
	wire signed [31:0] w_setValueToChildArray_bx_10_addr;
	wire signed [31:0] w_setValueToChildArray_bx_10_datain;
	wire               w_setValueToChildArray_bx_10_r_w;
	wire               w_setValueToChildArray_bx_10_ce;
	wire               w_setValueToChildArray_bx_10_cacheHit;
	reg  signed [31:0] r_setValueToChildArray_dataNum_11;
	reg  signed [31:0] r_setValueToChildArray_i_12;
	reg  signed [31:0] r_subRoutine_ax_13_addr;
	reg  signed [31:0] r_subRoutine_ax_13_datain;
	wire signed [31:0] w_subRoutine_ax_13_dataout;
	reg                r_subRoutine_ax_13_r_w;
	wire signed [31:0] w_subRoutine_ax_13_addr;
	wire signed [31:0] w_subRoutine_ax_13_datain;
	wire               w_subRoutine_ax_13_r_w;
	wire               w_subRoutine_ax_13_ce;
	wire               w_subRoutine_ax_13_cacheHit;
	reg  signed [31:0] r_subRoutine_bx_14_addr;
	reg  signed [31:0] r_subRoutine_bx_14_datain;
	wire signed [31:0] w_subRoutine_bx_14_dataout;
	reg                r_subRoutine_bx_14_r_w;
	wire signed [31:0] w_subRoutine_bx_14_addr;
	wire signed [31:0] w_subRoutine_bx_14_datain;
	wire               w_subRoutine_bx_14_r_w;
	wire               w_subRoutine_bx_14_ce;
	wire               w_subRoutine_bx_14_cacheHit;
	reg  signed [31:0] r_subRoutine_dataNum_15;
	reg  signed [31:0] r_subRoutine_i_16;
	reg  signed [31:0] r_subRoutine_ret_17;
	reg  signed [31:0] r_subRoutine_copy0_i_18;
	reg  signed [31:0] r_subRoutine_copy1_i_19;
	reg  signed [31:0] r_subRoutine_copy2_i_20;
	reg  signed [31:0] r_subRoutine_copy3_i_21;
	reg  signed [31:0] r_subRoutine_copy4_i_22;
	reg  signed [31:0] r_subRoutine_copy0_i_23;
	reg                r_subClassAX_subAprocess_req;
	wire               w_subClassAX_subAprocess_busy;
	wire signed [31:0] w_subClassAX_subAprocess_return;
	wire signed [ 4:0] w_subClassAX_arrayA_addr;
	reg  signed [ 4:0] r_subClassAX_arrayA_addr;
	wire signed [31:0] w_subClassAX_arrayA_datain;
	reg  signed [31:0] r_subClassAX_arrayA_datain;
	wire signed [31:0] w_subClassAX_arrayA_dataout;
	wire               w_subClassAX_arrayA_r_w;
	reg                r_subClassAX_arrayA_r_w;
	wire signed [31:0] w_subClassAX_subAprocess_ax_addr;
	wire signed [31:0] w_subClassAX_subAprocess_ax_datain;
	wire signed [31:0] w_subClassAX_subAprocess_ax_dataout;
	wire               w_subClassAX_subAprocess_ax_r_w;
	wire               w_subClassAX_subAprocess_ax_ce;
	wire signed [31:0] w_subClassAX_subAprocess_bx_addr;
	wire signed [31:0] w_subClassAX_subAprocess_bx_datain;
	wire signed [31:0] w_subClassAX_subAprocess_bx_dataout;
	wire               w_subClassAX_subAprocess_bx_r_w;
	wire               w_subClassAX_subAprocess_bx_ce;
	wire               w_subClassAX_subAprocess_bx_cacheHit;
	reg  signed [31:0] r_subClassAX_subAprocess_dataNum;
	reg                r_subClassA_subAprocess_req;
	wire               w_subClassA_subAprocess_busy;
	wire signed [31:0] w_subClassA_subAprocess_return;
	wire signed [ 4:0] w_subClassA_arrayA_addr;
	reg  signed [ 4:0] r_subClassA_arrayA_addr;
	wire signed [31:0] w_subClassA_arrayA_datain;
	reg  signed [31:0] r_subClassA_arrayA_datain;
	wire signed [31:0] w_subClassA_arrayA_dataout;
	wire               w_subClassA_arrayA_r_w;
	reg                r_subClassA_arrayA_r_w;
	wire signed [31:0] w_subClassA_subAprocess_ax_addr;
	wire signed [31:0] w_subClassA_subAprocess_ax_datain;
	wire signed [31:0] w_subClassA_subAprocess_ax_dataout;
	wire               w_subClassA_subAprocess_ax_r_w;
	wire               w_subClassA_subAprocess_ax_ce;
	wire signed [31:0] w_subClassA_subAprocess_bx_addr;
	wire signed [31:0] w_subClassA_subAprocess_bx_datain;
	wire signed [31:0] w_subClassA_subAprocess_bx_dataout;
	wire               w_subClassA_subAprocess_bx_r_w;
	wire               w_subClassA_subAprocess_bx_ce;
	wire               w_subClassA_subAprocess_bx_cacheHit;
	reg  signed [31:0] r_subClassA_subAprocess_dataNum;
	reg                r_subClassB_subBprocess_req;
	wire               w_subClassB_subBprocess_busy;
	wire signed [31:0] w_subClassB_subBprocess_return;
	wire signed [ 4:0] w_subClassB_arrayB_addr;
	reg  signed [ 4:0] r_subClassB_arrayB_addr;
	wire signed [31:0] w_subClassB_arrayB_datain;
	reg  signed [31:0] r_subClassB_arrayB_datain;
	wire signed [31:0] w_subClassB_arrayB_dataout;
	wire               w_subClassB_arrayB_r_w;
	reg                r_subClassB_arrayB_r_w;
	wire signed [31:0] w_subClassB_subBprocess_ax_addr;
	wire signed [31:0] w_subClassB_subBprocess_ax_datain;
	wire signed [31:0] w_subClassB_subBprocess_ax_dataout;
	wire               w_subClassB_subBprocess_ax_r_w;
	wire               w_subClassB_subBprocess_ax_ce;
	wire               w_subClassB_subBprocess_ax_cacheHit;
	wire signed [31:0] w_subClassB_subBprocess_bx_addr;
	wire signed [31:0] w_subClassB_subBprocess_bx_datain;
	wire signed [31:0] w_subClassB_subBprocess_bx_dataout;
	wire               w_subClassB_subBprocess_bx_r_w;
	wire               w_subClassB_subBprocess_bx_ce;
	reg  signed [31:0] r_subClassB_subBprocess_dataNum;
	reg  signed [31:0] r_sys_tmp0_int;
	reg  signed [31:0] r_sys_tmp1_int;
	reg  signed [31:0] r_sys_tmp2_int;
	reg  signed [31:0] r_sys_tmp3_int;
	wire        [31:0] w_sys_tmp1;
	wire signed [31:0] w_sys_tmp2;
	wire signed [31:0] w_sys_tmp3;
	wire               w_sys_tmp4;
	wire signed [31:0] w_sys_tmp7;
	wire signed [31:0] w_sys_tmp8;
	wire signed [31:0] w_sys_tmp10;
	wire signed [31:0] w_sys_tmp12;
	wire signed [31:0] w_sys_tmp13;
	wire signed [31:0] w_sys_tmp14;
	wire               w_sys_tmp15;
	wire signed [31:0] w_sys_tmp18;
	wire signed [31:0] w_sys_tmp19;
	wire signed [31:0] w_sys_tmp20;
	wire signed [31:0] w_sys_tmp22;
	wire signed [31:0] w_sys_tmp23;
	wire signed [31:0] w_sys_tmp24;
	wire signed [31:0] w_sys_tmp25;
	wire signed [31:0] w_sys_tmp26;
	wire signed [31:0] w_sys_tmp27;
	wire signed [31:0] w_sys_tmp28;
	wire signed [31:0] w_sys_tmp29;
	wire signed [31:0] w_sys_tmp30;
	wire signed [31:0] w_sys_tmp31;
	wire signed [31:0] w_sys_tmp33;
	wire signed [31:0] w_sys_tmp34;
	wire signed [31:0] w_sys_tmp35;
	wire signed [31:0] w_sys_tmp36;
	wire signed [31:0] w_sys_tmp38;
	wire signed [31:0] w_sys_tmp39;
	wire signed [31:0] w_sys_tmp40;
	wire signed [31:0] w_sys_tmp41;
	wire signed [31:0] w_sys_tmp42;
	wire               w_sys_tmp83;
	wire signed [31:0] w_sys_tmp85;
	wire signed [31:0] w_sys_tmp86;
	wire signed [31:0] w_sys_tmp87;
	wire signed [31:0] w_sys_tmp88;
	wire signed [31:0] w_sys_tmp89;
	wire signed [31:0] w_sys_tmp90;
	wire signed [31:0] w_sys_tmp109;
	wire signed [31:0] w_sys_tmp110;
	wire signed [31:0] w_sys_tmp111;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce & w_mainRoutine_arrayY_4_cacheHit & w_setValueToChildArray_ax_9_cacheHit & w_setValueToChildArray_bx_10_cacheHit & w_subRoutine_ax_13_cacheHit & w_subRoutine_bx_14_cacheHit;
	assign o_mainRoutine_busy = r_sys_mainRoutine_busy;
	assign o_mainRoutine_return = r_sys_mainRoutine_return;
	assign w_sys_mainRoutine_stage_p1 = (r_sys_mainRoutine_stage + 3'h1);
	assign w_sys_mainRoutine_step_p1 = (r_sys_mainRoutine_step + 4'h1);
	assign w_sys_setValueToChildArray_stage_p1 = (r_sys_setValueToChildArray_stage + 2'h1);
	assign w_sys_setValueToChildArray_step_p1 = (r_sys_setValueToChildArray_step + 3'h1);
	assign w_sys_subRoutine_stage_p1 = (r_sys_subRoutine_stage + 2'h1);
	assign w_sys_subRoutine_step_p1 = (r_sys_subRoutine_step + 3'h1);
	assign w_fld_arrayX_3_addr_0 = ( r_sys_subAprocess_arbiter1 ? $signed( w_subClassA_subAprocess_ax_addr[4:0] ) : ( r_sys_subBprocess_arbiter2 ? $signed( w_subClassB_subBprocess_bx_addr[4:0] ) : ( r_sys_setValueToChildArray_arbiter0 ? $signed( w_setValueToChildArray_bx_10_addr[4:0] ) : 5'sh0 )  )  ) ;
	assign w_fld_arrayX_3_datain_0 = ( r_sys_subAprocess_arbiter1 ? w_subClassA_subAprocess_ax_datain : ( r_sys_subBprocess_arbiter2 ? w_subClassB_subBprocess_bx_datain : ( r_sys_setValueToChildArray_arbiter0 ? w_setValueToChildArray_bx_10_datain : 32'sh0 )  )  ) ;
	assign w_fld_arrayX_3_r_w_0 = ( r_sys_subAprocess_arbiter1 ? w_subClassA_subAprocess_ax_r_w : ( r_sys_subBprocess_arbiter2 ? w_subClassB_subBprocess_bx_r_w : ( r_sys_setValueToChildArray_arbiter0 ? w_setValueToChildArray_bx_10_r_w : 1'h0 )  )  ) ;
	assign w_fld_arrayX_3_ce_0 = ( r_sys_subAprocess_arbiter1 ? w_subClassA_subAprocess_ax_ce : ( r_sys_subBprocess_arbiter2 ? w_subClassB_subBprocess_bx_ce : w_sys_ce )  ) ;
	assign w_fld_arrayX_3_ce_1 = w_sys_ce;
	assign w_mainRoutine_arrayY_4_dataout = i_mainRoutine_arrayY_4_dataout;
	assign w_mainRoutine_arrayY_4_addr = ( r_sys_subAprocess_arbiter1 ? w_subClassA_subAprocess_bx_addr : ( r_sys_subBprocess_arbiter2 ? w_subClassB_subBprocess_ax_addr : ( r_sys_setValueToChildArray_arbiter0 ? w_setValueToChildArray_ax_9_addr : r_mainRoutine_arrayY_4_addr )  )  ) ;
	assign w_mainRoutine_arrayY_4_datain = ( r_sys_subAprocess_arbiter1 ? w_subClassA_subAprocess_bx_datain : ( r_sys_subBprocess_arbiter2 ? w_subClassB_subBprocess_ax_datain : ( r_sys_setValueToChildArray_arbiter0 ? w_setValueToChildArray_ax_9_datain : r_mainRoutine_arrayY_4_datain )  )  ) ;
	assign w_mainRoutine_arrayY_4_r_w = ( r_sys_subAprocess_arbiter1 ? w_subClassA_subAprocess_bx_r_w : ( r_sys_subBprocess_arbiter2 ? w_subClassB_subBprocess_ax_r_w : ( r_sys_setValueToChildArray_arbiter0 ? w_setValueToChildArray_ax_9_r_w : r_mainRoutine_arrayY_4_r_w )  )  ) ;
	assign w_mainRoutine_arrayY_4_ce = ( r_sys_subAprocess_arbiter1 ? w_subClassA_subAprocess_bx_ce : ( r_sys_subBprocess_arbiter2 ? w_subClassB_subBprocess_ax_ce : w_sys_ce )  ) ;
	assign w_mainRoutine_arrayY_4_cacheHit = i_mainRoutine_arrayY_4_cacheHit;
	assign o_mainRoutine_arrayY_4_addr = w_mainRoutine_arrayY_4_addr;
	assign o_mainRoutine_arrayY_4_datain = w_mainRoutine_arrayY_4_datain;
	assign o_mainRoutine_arrayY_4_r_w = w_mainRoutine_arrayY_4_r_w;
	assign o_mainRoutine_arrayY_4_ce = w_mainRoutine_arrayY_4_ce;
	assign w_setValueToChildArray_ax_9_dataout = ( r_sys_setValueToChildArray_arbiter0 ? w_mainRoutine_arrayY_4_dataout : 32'sh0 ) ;
	assign w_setValueToChildArray_ax_9_addr = ( r_sys_subRoutine_arbiter3 ? w_subRoutine_ax_13_addr : r_setValueToChildArray_ax_9_addr ) ;
	assign w_setValueToChildArray_ax_9_datain = ( r_sys_subRoutine_arbiter3 ? w_subRoutine_ax_13_datain : r_setValueToChildArray_ax_9_datain ) ;
	assign w_setValueToChildArray_ax_9_r_w = ( r_sys_subRoutine_arbiter3 ? w_subRoutine_ax_13_r_w : r_setValueToChildArray_ax_9_r_w ) ;
	assign w_setValueToChildArray_ax_9_ce = w_sys_ce;
	assign w_setValueToChildArray_ax_9_cacheHit = ( r_sys_setValueToChildArray_arbiter0 ? w_mainRoutine_arrayY_4_cacheHit : w_sys_boolTrue ) ;
	assign w_setValueToChildArray_bx_10_dataout = ( r_sys_setValueToChildArray_arbiter0 ? w_fld_arrayX_3_dataout_0 : 32'sh0 ) ;
	assign w_setValueToChildArray_bx_10_addr = ( r_sys_subRoutine_arbiter3 ? w_subRoutine_bx_14_addr : r_setValueToChildArray_bx_10_addr ) ;
	assign w_setValueToChildArray_bx_10_datain = ( r_sys_subRoutine_arbiter3 ? w_subRoutine_bx_14_datain : r_setValueToChildArray_bx_10_datain ) ;
	assign w_setValueToChildArray_bx_10_r_w = ( r_sys_subRoutine_arbiter3 ? w_subRoutine_bx_14_r_w : r_setValueToChildArray_bx_10_r_w ) ;
	assign w_setValueToChildArray_bx_10_ce = w_sys_ce;
	assign w_setValueToChildArray_bx_10_cacheHit = ( r_sys_setValueToChildArray_arbiter0 ? w_sys_boolTrue : w_sys_boolTrue ) ;
	assign w_subRoutine_ax_13_dataout = ( r_sys_subRoutine_arbiter3 ? w_setValueToChildArray_ax_9_dataout : 32'sh0 ) ;
	assign w_subRoutine_ax_13_addr = r_subRoutine_ax_13_addr;
	assign w_subRoutine_ax_13_datain = r_subRoutine_ax_13_datain;
	assign w_subRoutine_ax_13_r_w = r_subRoutine_ax_13_r_w;
	assign w_subRoutine_ax_13_ce = w_sys_ce;
	assign w_subRoutine_ax_13_cacheHit = ( r_sys_subRoutine_arbiter3 ? w_setValueToChildArray_ax_9_cacheHit : w_sys_boolTrue ) ;
	assign w_subRoutine_bx_14_dataout = ( r_sys_subRoutine_arbiter3 ? w_setValueToChildArray_bx_10_dataout : 32'sh0 ) ;
	assign w_subRoutine_bx_14_addr = r_subRoutine_bx_14_addr;
	assign w_subRoutine_bx_14_datain = r_subRoutine_bx_14_datain;
	assign w_subRoutine_bx_14_r_w = r_subRoutine_bx_14_r_w;
	assign w_subRoutine_bx_14_ce = w_sys_ce;
	assign w_subRoutine_bx_14_cacheHit = ( r_sys_subRoutine_arbiter3 ? w_setValueToChildArray_bx_10_cacheHit : w_sys_boolTrue ) ;
	assign w_subClassAX_arrayA_addr = ( (|r_sys_processing_methodID) ? r_subClassAX_arrayA_addr : 5'sh0 ) ;
	assign w_subClassAX_arrayA_datain = ( (|r_sys_processing_methodID) ? r_subClassAX_arrayA_datain : 32'sh0 ) ;
	assign w_subClassAX_arrayA_r_w = ( (|r_sys_processing_methodID) ? r_subClassAX_arrayA_r_w : 1'h0 ) ;
	assign w_subClassAX_subAprocess_ax_dataout = 32'sh0;
	assign w_subClassAX_subAprocess_bx_dataout = 32'sh0;
	assign w_subClassAX_subAprocess_bx_cacheHit = 1'b1;
	assign w_subClassA_arrayA_addr = ( (|r_sys_processing_methodID) ? r_subClassA_arrayA_addr : 5'sh0 ) ;
	assign w_subClassA_arrayA_datain = ( (|r_sys_processing_methodID) ? r_subClassA_arrayA_datain : 32'sh0 ) ;
	assign w_subClassA_arrayA_r_w = ( (|r_sys_processing_methodID) ? r_subClassA_arrayA_r_w : 1'h0 ) ;
	assign w_subClassA_subAprocess_ax_dataout = ( r_sys_subAprocess_arbiter1 ? w_fld_arrayX_3_dataout_0 : 32'sh0 ) ;
	assign w_subClassA_subAprocess_bx_dataout = ( r_sys_subAprocess_arbiter1 ? w_mainRoutine_arrayY_4_dataout : 32'sh0 ) ;
	assign w_subClassA_subAprocess_bx_cacheHit = ( r_sys_subAprocess_arbiter1 ? w_mainRoutine_arrayY_4_cacheHit : 1'b1 ) ;
	assign w_subClassB_arrayB_addr = ( (|r_sys_processing_methodID) ? r_subClassB_arrayB_addr : 5'sh0 ) ;
	assign w_subClassB_arrayB_datain = ( (|r_sys_processing_methodID) ? r_subClassB_arrayB_datain : 32'sh0 ) ;
	assign w_subClassB_arrayB_r_w = ( (|r_sys_processing_methodID) ? r_subClassB_arrayB_r_w : 1'h0 ) ;
	assign w_subClassB_subBprocess_ax_dataout = ( r_sys_subBprocess_arbiter2 ? w_mainRoutine_arrayY_4_dataout : 32'sh0 ) ;
	assign w_subClassB_subBprocess_ax_cacheHit = ( r_sys_subBprocess_arbiter2 ? w_mainRoutine_arrayY_4_cacheHit : 1'b1 ) ;
	assign w_subClassB_subBprocess_bx_dataout = ( r_sys_subBprocess_arbiter2 ? w_fld_arrayX_3_dataout_0 : 32'sh0 ) ;
	assign w_sys_tmp1 = w_ip_FixedToFloat_floating_0;
	assign w_sys_tmp2 = (w_sys_tmp3 + r_mainRoutine_subXRet_8);
	assign w_sys_tmp3 = (r_mainRoutine_subARet_6 + r_mainRoutine_subBRet_7);
	assign w_sys_tmp4 = (r_setValueToChildArray_i_12 < r_setValueToChildArray_dataNum_11);
	assign w_sys_tmp7 = (w_sys_tmp8 + w_sys_intOne);
	assign w_sys_tmp8 = (r_setValueToChildArray_i_12 + r_setValueToChildArray_i_12);
	assign w_sys_tmp10 = 32'sh0000000a;
	assign w_sys_tmp12 = w_subClassA_arrayA_dataout;
	assign w_sys_tmp13 = (r_setValueToChildArray_i_12 + w_sys_intOne);
	assign w_sys_tmp14 = r_sys_subRoutine_return;
	assign w_sys_tmp15 = (r_subRoutine_i_16 < r_subRoutine_dataNum_15);
	assign w_sys_tmp18 = (w_sys_tmp19 * w_sys_tmp20);
	assign w_sys_tmp19 = (r_subRoutine_copy4_i_22 - r_subRoutine_dataNum_15);
	assign w_sys_tmp20 = (r_subRoutine_copy3_i_21 - r_subRoutine_dataNum_15);
	assign w_sys_tmp22 = (w_sys_tmp23 / w_sys_tmp25);
	assign w_sys_tmp23 = (w_sys_tmp24 + r_subRoutine_dataNum_15);
	assign w_sys_tmp24 = (r_subRoutine_copy1_i_19 + r_subRoutine_dataNum_15);
	assign w_sys_tmp25 = (r_subRoutine_copy0_i_18 - r_subRoutine_dataNum_15);
	assign w_sys_tmp26 = (r_subRoutine_copy0_i_18 + w_sys_intOne);
	assign w_sys_tmp27 = (r_subRoutine_copy1_i_19 + w_sys_intOne);
	assign w_sys_tmp28 = (r_subRoutine_copy2_i_20 + w_sys_intOne);
	assign w_sys_tmp29 = (r_subRoutine_copy3_i_21 + w_sys_intOne);
	assign w_sys_tmp30 = (r_subRoutine_copy4_i_22 + w_sys_intOne);
	assign w_sys_tmp31 = (r_subRoutine_i_16 + w_sys_intOne);
	assign w_sys_tmp33 = (w_sys_tmp34 - r_subRoutine_dataNum_15);
	assign w_sys_tmp34 = w_sys_tmp30;
	assign w_sys_tmp35 = (w_sys_tmp36 - r_subRoutine_dataNum_15);
	assign w_sys_tmp36 = w_sys_tmp29;
	assign w_sys_tmp38 = (w_sys_tmp39 + r_subRoutine_dataNum_15);
	assign w_sys_tmp39 = (w_sys_tmp40 + r_subRoutine_dataNum_15);
	assign w_sys_tmp40 = w_sys_tmp27;
	assign w_sys_tmp41 = (w_sys_tmp42 - r_subRoutine_dataNum_15);
	assign w_sys_tmp42 = w_sys_tmp26;
	assign w_sys_tmp83 = (r_subRoutine_i_16 < r_subRoutine_dataNum_15);
	assign w_sys_tmp85 = (r_subRoutine_ret_17 + w_sys_tmp86);
	assign w_sys_tmp86 = (w_sys_tmp87 + w_sys_tmp88);
	assign w_sys_tmp87 = w_subRoutine_ax_13_dataout;
	assign w_sys_tmp88 = w_subRoutine_bx_14_dataout;
	assign w_sys_tmp89 = (r_subRoutine_copy0_i_23 + w_sys_intOne);
	assign w_sys_tmp90 = (r_subRoutine_i_16 + w_sys_intOne);
	assign w_sys_tmp109 = r_subRoutine_ret_17;
	assign w_sys_tmp110 = (w_sys_tmp33 * w_sys_tmp35);
	assign w_sys_tmp111 = (w_sys_tmp38 / w_sys_tmp41);


	SubClassA
		subClassAX_inst(
			.i_fld_arrayA_0_addr_0 (w_subClassAX_arrayA_addr),
			.i_fld_arrayA_0_datain_0 (w_subClassAX_arrayA_datain),
			.o_fld_arrayA_0_dataout_0 (w_subClassAX_arrayA_dataout),
			.i_fld_arrayA_0_r_w_0 (w_subClassAX_arrayA_r_w),
			.o_subAprocess_ax_1_addr (w_subClassAX_subAprocess_ax_addr),
			.o_subAprocess_ax_1_ce (w_subClassAX_subAprocess_ax_ce),
			.o_subAprocess_ax_1_datain (w_subClassAX_subAprocess_ax_datain),
			.i_subAprocess_ax_1_dataout (w_subClassAX_subAprocess_ax_dataout),
			.o_subAprocess_ax_1_r_w (w_subClassAX_subAprocess_ax_r_w),
			.o_subAprocess_busy (w_subClassAX_subAprocess_busy),
			.o_subAprocess_bx_2_addr (w_subClassAX_subAprocess_bx_addr),
			.i_subAprocess_bx_2_cacheHit (w_subClassAX_subAprocess_bx_cacheHit),
			.o_subAprocess_bx_2_ce (w_subClassAX_subAprocess_bx_ce),
			.o_subAprocess_bx_2_datain (w_subClassAX_subAprocess_bx_datain),
			.i_subAprocess_bx_2_dataout (w_subClassAX_subAprocess_bx_dataout),
			.o_subAprocess_bx_2_r_w (w_subClassAX_subAprocess_bx_r_w),
			.i_subAprocess_dataNum_3 (r_subClassAX_subAprocess_dataNum),
			.i_subAprocess_req (r_subClassAX_subAprocess_req),
			.o_subAprocess_return (w_subClassAX_subAprocess_return),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	SubClassA
		subClassA_inst(
			.i_fld_arrayA_0_addr_0 (w_subClassA_arrayA_addr),
			.i_fld_arrayA_0_datain_0 (w_subClassA_arrayA_datain),
			.o_fld_arrayA_0_dataout_0 (w_subClassA_arrayA_dataout),
			.i_fld_arrayA_0_r_w_0 (w_subClassA_arrayA_r_w),
			.o_subAprocess_ax_1_addr (w_subClassA_subAprocess_ax_addr),
			.o_subAprocess_ax_1_ce (w_subClassA_subAprocess_ax_ce),
			.o_subAprocess_ax_1_datain (w_subClassA_subAprocess_ax_datain),
			.i_subAprocess_ax_1_dataout (w_subClassA_subAprocess_ax_dataout),
			.o_subAprocess_ax_1_r_w (w_subClassA_subAprocess_ax_r_w),
			.o_subAprocess_busy (w_subClassA_subAprocess_busy),
			.o_subAprocess_bx_2_addr (w_subClassA_subAprocess_bx_addr),
			.i_subAprocess_bx_2_cacheHit (w_subClassA_subAprocess_bx_cacheHit),
			.o_subAprocess_bx_2_ce (w_subClassA_subAprocess_bx_ce),
			.o_subAprocess_bx_2_datain (w_subClassA_subAprocess_bx_datain),
			.i_subAprocess_bx_2_dataout (w_subClassA_subAprocess_bx_dataout),
			.o_subAprocess_bx_2_r_w (w_subClassA_subAprocess_bx_r_w),
			.i_subAprocess_dataNum_3 (r_subClassA_subAprocess_dataNum),
			.i_subAprocess_req (r_subClassA_subAprocess_req),
			.o_subAprocess_return (w_subClassA_subAprocess_return),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	SubClassB
		subClassB_inst(
			.i_fld_arrayB_0_addr_0 (w_subClassB_arrayB_addr),
			.i_fld_arrayB_0_datain_0 (w_subClassB_arrayB_datain),
			.o_fld_arrayB_0_dataout_0 (w_subClassB_arrayB_dataout),
			.i_fld_arrayB_0_r_w_0 (w_subClassB_arrayB_r_w),
			.o_subBprocess_ax_1_addr (w_subClassB_subBprocess_ax_addr),
			.i_subBprocess_ax_1_cacheHit (w_subClassB_subBprocess_ax_cacheHit),
			.o_subBprocess_ax_1_ce (w_subClassB_subBprocess_ax_ce),
			.o_subBprocess_ax_1_datain (w_subClassB_subBprocess_ax_datain),
			.i_subBprocess_ax_1_dataout (w_subClassB_subBprocess_ax_dataout),
			.o_subBprocess_ax_1_r_w (w_subClassB_subBprocess_ax_r_w),
			.o_subBprocess_busy (w_subClassB_subBprocess_busy),
			.o_subBprocess_bx_2_addr (w_subClassB_subBprocess_bx_addr),
			.o_subBprocess_bx_2_ce (w_subClassB_subBprocess_bx_ce),
			.o_subBprocess_bx_2_datain (w_subClassB_subBprocess_bx_datain),
			.i_subBprocess_bx_2_dataout (w_subClassB_subBprocess_bx_dataout),
			.o_subBprocess_bx_2_r_w (w_subClassB_subBprocess_bx_r_w),
			.i_subBprocess_dataNum_3 (r_subClassB_subBprocess_dataNum),
			.i_subBprocess_req (r_subClassB_subBprocess_req),
			.o_subBprocess_return (w_subClassB_subBprocess_return),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(5), .WORDS(32) )
		dpram_arrayX_3(
			.clk (clock),
			.ce_0 (w_fld_arrayX_3_ce_0),
			.addr_0 (w_fld_arrayX_3_addr_0),
			.datain_0 (w_fld_arrayX_3_datain_0),
			.dataout_0 (w_fld_arrayX_3_dataout_0),
			.r_w_0 (w_fld_arrayX_3_r_w_0),
			.ce_1 (w_fld_arrayX_3_ce_1),
			.addr_1 (r_fld_arrayX_3_addr_1),
			.datain_1 (r_fld_arrayX_3_datain_1),
			.dataout_1 (w_fld_arrayX_3_dataout_1),
			.r_w_1 (r_fld_arrayX_3_r_w_1)
		);

	FixedToFloat
		FixedToFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_FixedToFloat_fixed_0),
			.result (w_ip_FixedToFloat_floating_0)
		);

	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_setValueToChildArray_arbiter0 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_mainRoutine_phase) 
						3'h2: begin

							case(r_sys_mainRoutine_stage) 
								3'h1: begin
									if((r_sys_mainRoutine_step==4'h1)) begin
										r_sys_setValueToChildArray_arbiter0 <= w_sys_boolFalse;

									end
									else
									if((r_sys_mainRoutine_step==4'h0)) begin
										r_sys_setValueToChildArray_arbiter0 <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_subAprocess_arbiter1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_mainRoutine_phase) 
						3'h2: begin

							case(r_sys_mainRoutine_stage) 
								3'h2: begin
									if((r_sys_mainRoutine_step==4'h0)) begin
										r_sys_subAprocess_arbiter1 <= w_sys_boolTrue;

									end
									else
									if((r_sys_mainRoutine_step==4'h2)) begin
										r_sys_subAprocess_arbiter1 <= ((w_subClassA_subAprocess_busy) ? w_sys_boolTrue : w_sys_boolFalse);

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_subBprocess_arbiter2 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_mainRoutine_phase) 
						3'h2: begin

							case(r_sys_mainRoutine_stage) 
								3'h3: begin
									if((r_sys_mainRoutine_step==4'h0)) begin
										r_sys_subBprocess_arbiter2 <= w_sys_boolTrue;

									end
									else
									if((r_sys_mainRoutine_step==4'h2)) begin
										r_sys_subBprocess_arbiter2 <= ((w_subClassB_subBprocess_busy) ? w_sys_boolTrue : w_sys_boolFalse);

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_subRoutine_arbiter3 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h9: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h1)) begin
										r_sys_subRoutine_arbiter3 <= w_sys_boolFalse;

									end
									else
									if((r_sys_setValueToChildArray_step==3'h0)) begin
										r_sys_subRoutine_arbiter3 <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_mainRoutine_phase) 
						3'h4: begin

							case(r_sys_mainRoutine_stage) 
								3'h0: begin
									if((r_sys_mainRoutine_step==4'h0)) begin
										r_ip_FixedToFloat_fixed_0 <= w_sys_tmp2;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 3'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h0: begin
					r_sys_processing_methodID <= ((i_mainRoutine_req) ? 3'h1 : r_sys_processing_methodID);
				end

				3'h1: begin

					case(r_sys_mainRoutine_phase) 
						3'h2: begin

							case(r_sys_mainRoutine_stage) 
								3'h1: begin
									if((r_sys_mainRoutine_step==4'h0)) begin
										r_sys_processing_methodID <= 3'h2;

									end
								end

							endcase
						end

						3'h6: begin
							r_sys_processing_methodID <= r_sys_mainRoutine_caller;
						end

					endcase
				end

				3'h2: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h9: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h0)) begin
										r_sys_processing_methodID <= 3'h3;

									end
								end

							endcase
						end

						4'hb: begin
							r_sys_processing_methodID <= r_sys_setValueToChildArray_caller;
						end

					endcase
				end

				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h13: begin
							r_sys_processing_methodID <= r_sys_subRoutine_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_mainRoutine_return <= 32'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_mainRoutine_phase) 
						3'h3: begin
							r_sys_mainRoutine_return <= w_sys_tmp1;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_mainRoutine_caller <= 3'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_mainRoutine_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_mainRoutine_phase <= 3'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_mainRoutine_phase) 
						3'h0: begin
							r_sys_mainRoutine_phase <= 3'h2;
						end

						3'h2: begin

							case(r_sys_mainRoutine_stage) 
								3'h3: begin
									if((r_sys_mainRoutine_step==4'h3)) begin
										r_sys_mainRoutine_phase <= 3'h4;

									end
								end

							endcase
						end

						3'h3: begin
							r_sys_mainRoutine_phase <= 3'h6;
						end

						3'h4: begin

							case(r_sys_mainRoutine_stage) 
								3'h0: begin
									if((r_sys_mainRoutine_step==4'h7)) begin
										r_sys_mainRoutine_phase <= 3'h3;

									end
								end

							endcase
						end

						3'h6: begin
							r_sys_mainRoutine_phase <= 3'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_mainRoutine_stage <= 3'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_mainRoutine_phase) 
						3'h2: begin

							case(r_sys_mainRoutine_stage) 
								3'h0: begin
									if((r_sys_mainRoutine_step==4'h0)) begin
										r_sys_mainRoutine_stage <= w_sys_mainRoutine_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_mainRoutine_step==4'h1)) begin
										r_sys_mainRoutine_stage <= w_sys_mainRoutine_stage_p1;

									end
								end

								3'h2: begin
									if((r_sys_mainRoutine_step==4'h3)) begin
										r_sys_mainRoutine_stage <= w_sys_mainRoutine_stage_p1;

									end
								end

								3'h3: begin
									if((r_sys_mainRoutine_step==4'h3)) begin
										r_sys_mainRoutine_stage <= 3'h0;

									end
								end

							endcase
						end

						3'h4: begin

							case(r_sys_mainRoutine_stage) 
								3'h0: begin
									if((r_sys_mainRoutine_step==4'h7)) begin
										r_sys_mainRoutine_stage <= 3'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_mainRoutine_step <= 4'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_mainRoutine_phase) 
						3'h2: begin

							case(r_sys_mainRoutine_stage) 
								3'h0: begin
									if((r_sys_mainRoutine_step==4'h0)) begin
										r_sys_mainRoutine_step <= 4'h0;

									end
								end

								3'h1: begin
									if((r_sys_mainRoutine_step==4'h0)) begin
										r_sys_mainRoutine_step <= w_sys_mainRoutine_step_p1;

									end
									else
									if((r_sys_mainRoutine_step==4'h1)) begin
										r_sys_mainRoutine_step <= 4'h0;

									end
								end

								3'h2: begin
									if((r_sys_mainRoutine_step==4'h2)) begin
										r_sys_mainRoutine_step <= ((w_subClassA_subAprocess_busy) ? r_sys_mainRoutine_step : w_sys_mainRoutine_step_p1);

									end
									else
									if((r_sys_mainRoutine_step==4'h3)) begin
										r_sys_mainRoutine_step <= 4'h0;

									end
									else
									if((r_sys_mainRoutine_step==4'h0) || (r_sys_mainRoutine_step==4'h1)) begin
										r_sys_mainRoutine_step <= w_sys_mainRoutine_step_p1;

									end
								end

								3'h3: begin
									if((r_sys_mainRoutine_step==4'h3)) begin
										r_sys_mainRoutine_step <= 4'h0;

									end
									else
									if((r_sys_mainRoutine_step==4'h0) || (r_sys_mainRoutine_step==4'h1)) begin
										r_sys_mainRoutine_step <= w_sys_mainRoutine_step_p1;

									end
									else
									if((r_sys_mainRoutine_step==4'h2)) begin
										r_sys_mainRoutine_step <= ((w_subClassB_subBprocess_busy) ? r_sys_mainRoutine_step : w_sys_mainRoutine_step_p1);

									end
								end

							endcase
						end

						3'h4: begin

							case(r_sys_mainRoutine_stage) 
								3'h0: begin
									if((r_sys_mainRoutine_step==4'h7)) begin
										r_sys_mainRoutine_step <= 4'h0;

									end
									else
									if((4'h0<=r_sys_mainRoutine_step && r_sys_mainRoutine_step<=4'h6)) begin
										r_sys_mainRoutine_step <= w_sys_mainRoutine_step_p1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_mainRoutine_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h0: begin
					r_sys_mainRoutine_busy <= ((i_mainRoutine_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				3'h1: begin

					case(r_sys_mainRoutine_phase) 
						3'h0: begin
							r_sys_mainRoutine_busy <= w_sys_boolTrue;
						end

						3'h6: begin
							r_sys_mainRoutine_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_setValueToChildArray_return <= 32'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h8: begin
							r_sys_setValueToChildArray_return <= w_sys_tmp14;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_setValueToChildArray_caller <= 3'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_mainRoutine_phase) 
						3'h2: begin

							case(r_sys_mainRoutine_stage) 
								3'h1: begin
									if((r_sys_mainRoutine_step==4'h0)) begin
										r_sys_setValueToChildArray_caller <= r_sys_processing_methodID;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_setValueToChildArray_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_setValueToChildArray_phase <= 4'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h0: begin
							r_sys_setValueToChildArray_phase <= 4'h3;
						end

						4'h3: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h0)) begin
										r_sys_setValueToChildArray_phase <= 4'h4;

									end
								end

							endcase
						end

						4'h4: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h0)) begin
										r_sys_setValueToChildArray_phase <= ((w_sys_tmp4) ? 4'h7 : 4'h9);

									end
								end

							endcase
						end

						4'h7: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h3)) begin
										r_sys_setValueToChildArray_phase <= 4'h4;

									end
								end

							endcase
						end

						4'h8: begin
							r_sys_setValueToChildArray_phase <= 4'hb;
						end

						4'h9: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h1)) begin
										r_sys_setValueToChildArray_phase <= 4'h8;

									end
								end

							endcase
						end

						4'hb: begin
							r_sys_setValueToChildArray_phase <= 4'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_setValueToChildArray_stage <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h3: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h0)) begin
										r_sys_setValueToChildArray_stage <= 2'h0;

									end
								end

							endcase
						end

						4'h4: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h0)) begin
										r_sys_setValueToChildArray_stage <= 2'h0;

									end
								end

							endcase
						end

						4'h7: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h3)) begin
										r_sys_setValueToChildArray_stage <= 2'h0;

									end
								end

							endcase
						end

						4'h9: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h1)) begin
										r_sys_setValueToChildArray_stage <= 2'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_setValueToChildArray_step <= 3'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h3: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h0)) begin
										r_sys_setValueToChildArray_step <= 3'h0;

									end
								end

							endcase
						end

						4'h4: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h0)) begin
										r_sys_setValueToChildArray_step <= 3'h0;

									end
								end

							endcase
						end

						4'h7: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h0) || (r_sys_setValueToChildArray_step==3'h1) || (r_sys_setValueToChildArray_step==3'h2)) begin
										r_sys_setValueToChildArray_step <= w_sys_setValueToChildArray_step_p1;

									end
									else
									if((r_sys_setValueToChildArray_step==3'h3)) begin
										r_sys_setValueToChildArray_step <= 3'h0;

									end
								end

							endcase
						end

						4'h9: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h1)) begin
										r_sys_setValueToChildArray_step <= 3'h0;

									end
									else
									if((r_sys_setValueToChildArray_step==3'h0)) begin
										r_sys_setValueToChildArray_step <= w_sys_setValueToChildArray_step_p1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_setValueToChildArray_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h0: begin
							r_sys_setValueToChildArray_busy <= w_sys_boolTrue;
						end

						4'hb: begin
							r_sys_setValueToChildArray_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_subRoutine_return <= 32'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h10: begin
							r_sys_subRoutine_return <= w_sys_tmp109;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_subRoutine_caller <= 3'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h9: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h0)) begin
										r_sys_subRoutine_caller <= r_sys_processing_methodID;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_subRoutine_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_subRoutine_phase <= 5'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h0: begin
							r_sys_subRoutine_phase <= 5'h2;
						end

						5'h2: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_sys_subRoutine_phase <= 5'h4;

									end
								end

							endcase
						end

						5'h4: begin

							case(r_sys_subRoutine_stage) 
								2'h1: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_sys_subRoutine_phase <= 5'h5;

									end
								end

							endcase
						end

						5'h5: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_sys_subRoutine_phase <= ((w_sys_tmp15) ? 5'h8 : 5'h9);

									end
								end

							endcase
						end

						5'h8: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h3)) begin
										r_sys_subRoutine_phase <= 5'h5;

									end
								end

							endcase
						end

						5'h9: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_sys_subRoutine_phase <= 5'hb;

									end
								end

							endcase
						end

						5'hb: begin

							case(r_sys_subRoutine_stage) 
								2'h1: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_sys_subRoutine_phase <= 5'hc;

									end
								end

							endcase
						end

						5'hc: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_sys_subRoutine_phase <= ((w_sys_tmp83) ? 5'hf : 5'h11);

									end
								end

							endcase
						end

						5'hf: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h5)) begin
										r_sys_subRoutine_phase <= 5'hc;

									end
								end

							endcase
						end

						5'h10: begin
							r_sys_subRoutine_phase <= 5'h13;
						end

						5'h11: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_sys_subRoutine_phase <= 5'h10;

									end
								end

							endcase
						end

						5'h13: begin
							r_sys_subRoutine_phase <= 5'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_subRoutine_stage <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h2: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_sys_subRoutine_stage <= 2'h0;

									end
								end

							endcase
						end

						5'h4: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_sys_subRoutine_stage <= w_sys_subRoutine_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_sys_subRoutine_stage <= 2'h0;

									end
								end

							endcase
						end

						5'h5: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_sys_subRoutine_stage <= 2'h0;

									end
								end

							endcase
						end

						5'h8: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h3)) begin
										r_sys_subRoutine_stage <= 2'h0;

									end
								end

							endcase
						end

						5'h9: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_sys_subRoutine_stage <= 2'h0;

									end
								end

							endcase
						end

						5'hb: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_sys_subRoutine_stage <= w_sys_subRoutine_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_sys_subRoutine_stage <= 2'h0;

									end
								end

							endcase
						end

						5'hc: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_sys_subRoutine_stage <= 2'h0;

									end
								end

							endcase
						end

						5'hf: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h5)) begin
										r_sys_subRoutine_stage <= 2'h0;

									end
								end

							endcase
						end

						5'h11: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_sys_subRoutine_stage <= 2'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_subRoutine_step <= 3'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h2: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_sys_subRoutine_step <= 3'h0;

									end
								end

							endcase
						end

						5'h4: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_sys_subRoutine_step <= 3'h0;

									end
								end

								2'h1: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_sys_subRoutine_step <= 3'h0;

									end
								end

							endcase
						end

						5'h5: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_sys_subRoutine_step <= 3'h0;

									end
								end

							endcase
						end

						5'h8: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h3)) begin
										r_sys_subRoutine_step <= 3'h0;

									end
									else
									if((r_sys_subRoutine_step==3'h0) || (r_sys_subRoutine_step==3'h1) || (r_sys_subRoutine_step==3'h2)) begin
										r_sys_subRoutine_step <= w_sys_subRoutine_step_p1;

									end
								end

							endcase
						end

						5'h9: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_sys_subRoutine_step <= 3'h0;

									end
								end

							endcase
						end

						5'hb: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_sys_subRoutine_step <= 3'h0;

									end
								end

								2'h1: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_sys_subRoutine_step <= 3'h0;

									end
								end

							endcase
						end

						5'hc: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_sys_subRoutine_step <= 3'h0;

									end
								end

							endcase
						end

						5'hf: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h5)) begin
										r_sys_subRoutine_step <= 3'h0;

									end
									else
									if((3'h0<=r_sys_subRoutine_step && r_sys_subRoutine_step<=3'h4)) begin
										r_sys_subRoutine_step <= w_sys_subRoutine_step_p1;

									end
								end

							endcase
						end

						5'h11: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_sys_subRoutine_step <= 3'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_subRoutine_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h0: begin
							r_sys_subRoutine_busy <= w_sys_boolTrue;
						end

						5'h13: begin
							r_sys_subRoutine_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_arrayX_3_addr_1 <= 5'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_arrayX_3_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_mainRoutine_phase) 
						3'h6: begin
							r_fld_arrayX_3_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

				3'h2: begin

					case(r_sys_setValueToChildArray_phase) 
						4'hb: begin
							r_fld_arrayX_3_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h13: begin
							r_fld_arrayX_3_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_mainRoutine_arrayY_4_addr <= 32'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_mainRoutine_arrayY_4_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_mainRoutine_phase) 
						3'h6: begin
							r_mainRoutine_arrayY_4_r_w <= w_sys_boolFalse;
						end

					endcase
				end

				3'h2: begin

					case(r_sys_setValueToChildArray_phase) 
						4'hb: begin
							r_mainRoutine_arrayY_4_r_w <= w_sys_boolFalse;
						end

					endcase
				end

				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h13: begin
							r_mainRoutine_arrayY_4_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h0: begin
					r_mainRoutine_dataNum_5 <= ((i_mainRoutine_req) ? i_mainRoutine_dataNum_5 : r_mainRoutine_dataNum_5);
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_mainRoutine_phase) 
						3'h2: begin

							case(r_sys_mainRoutine_stage) 
								3'h0: begin
									if((r_sys_mainRoutine_step==4'h0)) begin
										r_mainRoutine_subARet_6 <= w_sys_intZero;

									end
								end

								3'h2: begin
									if((r_sys_mainRoutine_step==4'h3)) begin
										r_mainRoutine_subARet_6 <= w_subClassA_subAprocess_return;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_mainRoutine_phase) 
						3'h2: begin

							case(r_sys_mainRoutine_stage) 
								3'h0: begin
									if((r_sys_mainRoutine_step==4'h0)) begin
										r_mainRoutine_subBRet_7 <= w_sys_intZero;

									end
								end

								3'h3: begin
									if((r_sys_mainRoutine_step==4'h3)) begin
										r_mainRoutine_subBRet_7 <= w_subClassB_subBprocess_return;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_mainRoutine_phase) 
						3'h2: begin

							case(r_sys_mainRoutine_stage) 
								3'h0: begin
									if((r_sys_mainRoutine_step==4'h0)) begin
										r_mainRoutine_subXRet_8 <= w_sys_intZero;

									end
								end

								3'h1: begin
									if((r_sys_mainRoutine_step==4'h1)) begin
										r_mainRoutine_subXRet_8 <= r_sys_setValueToChildArray_return;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_setValueToChildArray_ax_9_addr <= 32'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_setValueToChildArray_ax_9_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_mainRoutine_phase) 
						3'h6: begin
							r_setValueToChildArray_ax_9_r_w <= w_sys_boolFalse;
						end

					endcase
				end

				3'h2: begin

					case(r_sys_setValueToChildArray_phase) 
						4'hb: begin
							r_setValueToChildArray_ax_9_r_w <= w_sys_boolFalse;
						end

					endcase
				end

				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h13: begin
							r_setValueToChildArray_ax_9_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_setValueToChildArray_bx_10_addr <= 32'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_setValueToChildArray_bx_10_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_mainRoutine_phase) 
						3'h6: begin
							r_setValueToChildArray_bx_10_r_w <= w_sys_boolFalse;
						end

					endcase
				end

				3'h2: begin

					case(r_sys_setValueToChildArray_phase) 
						4'hb: begin
							r_setValueToChildArray_bx_10_r_w <= w_sys_boolFalse;
						end

					endcase
				end

				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h13: begin
							r_setValueToChildArray_bx_10_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_mainRoutine_phase) 
						3'h2: begin

							case(r_sys_mainRoutine_stage) 
								3'h1: begin
									if((r_sys_mainRoutine_step==4'h0)) begin
										r_setValueToChildArray_dataNum_11 <= r_mainRoutine_dataNum_5;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h3: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h0)) begin
										r_setValueToChildArray_i_12 <= w_sys_intZero;

									end
								end

							endcase
						end

						4'h7: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h0)) begin
										r_setValueToChildArray_i_12 <= w_sys_tmp13;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_subRoutine_ax_13_addr <= 32'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h8: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_subRoutine_ax_13_addr <= r_subRoutine_i_16;

									end
									else
									if((r_sys_subRoutine_step==3'h1) || (r_sys_subRoutine_step==3'h2) || (r_sys_subRoutine_step==3'h3)) begin
										r_subRoutine_ax_13_addr <= r_sys_tmp1_int;

									end
								end

							endcase
						end

						5'hf: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h1) || (r_sys_subRoutine_step==3'h2) || (r_sys_subRoutine_step==3'h3)) begin
										r_subRoutine_ax_13_addr <= r_sys_tmp3_int;

									end
									else
									if((r_sys_subRoutine_step==3'h0)) begin
										r_subRoutine_ax_13_addr <= r_subRoutine_i_16;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h8: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_subRoutine_ax_13_datain <= w_sys_tmp18;

									end
									else
									if((r_sys_subRoutine_step==3'h1) || (r_sys_subRoutine_step==3'h2) || (r_sys_subRoutine_step==3'h3)) begin
										r_subRoutine_ax_13_datain <= r_sys_tmp0_int;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_subRoutine_ax_13_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_mainRoutine_phase) 
						3'h6: begin
							r_subRoutine_ax_13_r_w <= w_sys_boolFalse;
						end

					endcase
				end

				3'h2: begin

					case(r_sys_setValueToChildArray_phase) 
						4'hb: begin
							r_subRoutine_ax_13_r_w <= w_sys_boolFalse;
						end

					endcase
				end

				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h8: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((3'h0<=r_sys_subRoutine_step && r_sys_subRoutine_step<=3'h3)) begin
										r_subRoutine_ax_13_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						5'hf: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((3'h0<=r_sys_subRoutine_step && r_sys_subRoutine_step<=3'h3)) begin
										r_subRoutine_ax_13_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						5'h13: begin
							r_subRoutine_ax_13_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_subRoutine_bx_14_addr <= 32'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h8: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h1) || (r_sys_subRoutine_step==3'h2) || (r_sys_subRoutine_step==3'h3)) begin
										r_subRoutine_bx_14_addr <= r_sys_tmp2_int;

									end
									else
									if((r_sys_subRoutine_step==3'h0)) begin
										r_subRoutine_bx_14_addr <= r_subRoutine_copy2_i_20;

									end
								end

							endcase
						end

						5'hf: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h1) || (r_sys_subRoutine_step==3'h2) || (r_sys_subRoutine_step==3'h3)) begin
										r_subRoutine_bx_14_addr <= r_sys_tmp2_int;

									end
									else
									if((r_sys_subRoutine_step==3'h0)) begin
										r_subRoutine_bx_14_addr <= r_subRoutine_copy0_i_23;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h8: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h1) || (r_sys_subRoutine_step==3'h2) || (r_sys_subRoutine_step==3'h3)) begin
										r_subRoutine_bx_14_datain <= r_sys_tmp3_int;

									end
									else
									if((r_sys_subRoutine_step==3'h0)) begin
										r_subRoutine_bx_14_datain <= w_sys_tmp22;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_subRoutine_bx_14_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_mainRoutine_phase) 
						3'h6: begin
							r_subRoutine_bx_14_r_w <= w_sys_boolFalse;
						end

					endcase
				end

				3'h2: begin

					case(r_sys_setValueToChildArray_phase) 
						4'hb: begin
							r_subRoutine_bx_14_r_w <= w_sys_boolFalse;
						end

					endcase
				end

				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h8: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((3'h0<=r_sys_subRoutine_step && r_sys_subRoutine_step<=3'h3)) begin
										r_subRoutine_bx_14_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						5'hf: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((3'h0<=r_sys_subRoutine_step && r_sys_subRoutine_step<=3'h3)) begin
										r_subRoutine_bx_14_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						5'h13: begin
							r_subRoutine_bx_14_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h9: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h0)) begin
										r_subRoutine_dataNum_15 <= r_setValueToChildArray_dataNum_11;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h2: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_subRoutine_i_16 <= w_sys_intZero;

									end
								end

							endcase
						end

						5'h4: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_subRoutine_i_16 <= w_sys_intZero;

									end
								end

							endcase
						end

						5'h8: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((3'h0<=r_sys_subRoutine_step && r_sys_subRoutine_step<=3'h3)) begin
										r_subRoutine_i_16 <= w_sys_tmp31;

									end
								end

							endcase
						end

						5'hb: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_subRoutine_i_16 <= w_sys_intZero;

									end
								end

							endcase
						end

						5'hf: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((3'h0<=r_sys_subRoutine_step && r_sys_subRoutine_step<=3'h3)) begin
										r_subRoutine_i_16 <= w_sys_tmp90;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h9: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_subRoutine_ret_17 <= w_sys_intZero;

									end
								end

							endcase
						end

						5'hf: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((3'h2<=r_sys_subRoutine_step && r_sys_subRoutine_step<=3'h5)) begin
										r_subRoutine_ret_17 <= w_sys_tmp85;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h4: begin

							case(r_sys_subRoutine_stage) 
								2'h1: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_subRoutine_copy0_i_18 <= r_subRoutine_i_16;

									end
								end

							endcase
						end

						5'h8: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((3'h0<=r_sys_subRoutine_step && r_sys_subRoutine_step<=3'h3)) begin
										r_subRoutine_copy0_i_18 <= w_sys_tmp26;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h4: begin

							case(r_sys_subRoutine_stage) 
								2'h1: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_subRoutine_copy1_i_19 <= r_subRoutine_i_16;

									end
								end

							endcase
						end

						5'h8: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((3'h0<=r_sys_subRoutine_step && r_sys_subRoutine_step<=3'h3)) begin
										r_subRoutine_copy1_i_19 <= w_sys_tmp27;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h4: begin

							case(r_sys_subRoutine_stage) 
								2'h1: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_subRoutine_copy2_i_20 <= r_subRoutine_i_16;

									end
								end

							endcase
						end

						5'h8: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((3'h0<=r_sys_subRoutine_step && r_sys_subRoutine_step<=3'h3)) begin
										r_subRoutine_copy2_i_20 <= w_sys_tmp28;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h4: begin

							case(r_sys_subRoutine_stage) 
								2'h1: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_subRoutine_copy3_i_21 <= r_subRoutine_i_16;

									end
								end

							endcase
						end

						5'h8: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((3'h0<=r_sys_subRoutine_step && r_sys_subRoutine_step<=3'h3)) begin
										r_subRoutine_copy3_i_21 <= w_sys_tmp29;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h4: begin

							case(r_sys_subRoutine_stage) 
								2'h1: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_subRoutine_copy4_i_22 <= r_subRoutine_i_16;

									end
								end

							endcase
						end

						5'h8: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((3'h0<=r_sys_subRoutine_step && r_sys_subRoutine_step<=3'h3)) begin
										r_subRoutine_copy4_i_22 <= w_sys_tmp30;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'hb: begin

							case(r_sys_subRoutine_stage) 
								2'h1: begin
									if((r_sys_subRoutine_step==3'h0)) begin
										r_subRoutine_copy0_i_23 <= r_subRoutine_i_16;

									end
								end

							endcase
						end

						5'hf: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((3'h0<=r_sys_subRoutine_step && r_sys_subRoutine_step<=3'h3)) begin
										r_subRoutine_copy0_i_23 <= w_sys_tmp89;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_subClassAX_subAprocess_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_subClassAX_arrayA_addr <= 5'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h7: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h0)) begin
										r_subClassAX_arrayA_addr <= $signed( r_setValueToChildArray_i_12[4:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h7: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h0)) begin
										r_subClassAX_arrayA_datain <= w_sys_tmp10;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_subClassAX_arrayA_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_mainRoutine_phase) 
						3'h2: begin

							case(r_sys_mainRoutine_stage) 
								3'h1: begin
									if((r_sys_mainRoutine_step==4'h0)) begin
										r_subClassAX_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_mainRoutine_step==4'h0)) begin
										r_subClassAX_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_mainRoutine_step==4'h0)) begin
										r_subClassAX_arrayA_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_subClassAX_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

				3'h2: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h7: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h0)) begin
										r_subClassAX_arrayA_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						4'h9: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h0)) begin
										r_subClassAX_arrayA_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						4'hb: begin
							r_subClassAX_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h13: begin
							r_subClassAX_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_subClassA_subAprocess_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_mainRoutine_phase) 
						3'h2: begin

							case(r_sys_mainRoutine_stage) 
								3'h2: begin
									if((r_sys_mainRoutine_step==4'h1)) begin
										r_subClassA_subAprocess_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_mainRoutine_step==4'h0)) begin
										r_subClassA_subAprocess_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_subClassA_arrayA_addr <= 5'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h7: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h0)) begin
										r_subClassA_arrayA_addr <= $signed( r_setValueToChildArray_i_12[4:0] );

									end
									else
									if((r_sys_setValueToChildArray_step==3'h1)) begin
										r_subClassA_arrayA_addr <= $signed( r_sys_tmp0_int[4:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h7: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h0)) begin
										r_subClassA_arrayA_datain <= w_sys_tmp7;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_subClassA_arrayA_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_mainRoutine_phase) 
						3'h2: begin

							case(r_sys_mainRoutine_stage) 
								3'h1: begin
									if((r_sys_mainRoutine_step==4'h0)) begin
										r_subClassA_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_mainRoutine_step==4'h0)) begin
										r_subClassA_arrayA_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_mainRoutine_step==4'h0)) begin
										r_subClassA_arrayA_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_subClassA_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

				3'h2: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h7: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h1)) begin
										r_subClassA_arrayA_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_setValueToChildArray_step==3'h0)) begin
										r_subClassA_arrayA_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						4'h9: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h0)) begin
										r_subClassA_arrayA_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						4'hb: begin
							r_subClassA_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h13: begin
							r_subClassA_arrayA_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_mainRoutine_phase) 
						3'h2: begin

							case(r_sys_mainRoutine_stage) 
								3'h2: begin
									if((r_sys_mainRoutine_step==4'h0)) begin
										r_subClassA_subAprocess_dataNum <= r_mainRoutine_dataNum_5;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_subClassB_subBprocess_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_mainRoutine_phase) 
						3'h2: begin

							case(r_sys_mainRoutine_stage) 
								3'h3: begin
									if((r_sys_mainRoutine_step==4'h1)) begin
										r_subClassB_subBprocess_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_mainRoutine_step==4'h0)) begin
										r_subClassB_subBprocess_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_subClassB_arrayB_addr <= 5'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h7: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h3)) begin
										r_subClassB_arrayB_addr <= $signed( r_sys_tmp1_int[4:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h7: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h3)) begin
										r_subClassB_arrayB_datain <= w_sys_tmp12;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_subClassB_arrayB_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_mainRoutine_phase) 
						3'h2: begin

							case(r_sys_mainRoutine_stage) 
								3'h1: begin
									if((r_sys_mainRoutine_step==4'h0)) begin
										r_subClassB_arrayB_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_mainRoutine_step==4'h0)) begin
										r_subClassB_arrayB_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_mainRoutine_step==4'h0)) begin
										r_subClassB_arrayB_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						3'h6: begin
							r_subClassB_arrayB_r_w <= w_sys_boolFalse;
						end

					endcase
				end

				3'h2: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h7: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h3)) begin
										r_subClassB_arrayB_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						4'h9: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h0)) begin
										r_subClassB_arrayB_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						4'hb: begin
							r_subClassB_arrayB_r_w <= w_sys_boolFalse;
						end

					endcase
				end

				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h13: begin
							r_subClassB_arrayB_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h1: begin

					case(r_sys_mainRoutine_phase) 
						3'h2: begin

							case(r_sys_mainRoutine_stage) 
								3'h3: begin
									if((r_sys_mainRoutine_step==4'h0)) begin
										r_subClassB_subBprocess_dataNum <= r_mainRoutine_dataNum_5;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h7: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h0)) begin
										r_sys_tmp0_int <= r_setValueToChildArray_i_12;

									end
								end

							endcase
						end

					endcase
				end

				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h8: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0) || (r_sys_subRoutine_step==3'h1) || (r_sys_subRoutine_step==3'h2)) begin
										r_sys_tmp0_int <= w_sys_tmp110;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h2: begin

					case(r_sys_setValueToChildArray_phase) 
						4'h7: begin

							case(r_sys_setValueToChildArray_stage) 
								2'h0: begin
									if((r_sys_setValueToChildArray_step==3'h0)) begin
										r_sys_tmp1_int <= r_setValueToChildArray_i_12;

									end
								end

							endcase
						end

					endcase
				end

				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h8: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0) || (r_sys_subRoutine_step==3'h1) || (r_sys_subRoutine_step==3'h2)) begin
										r_sys_tmp1_int <= w_sys_tmp31;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h8: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0) || (r_sys_subRoutine_step==3'h1) || (r_sys_subRoutine_step==3'h2)) begin
										r_sys_tmp2_int <= w_sys_tmp28;

									end
								end

							endcase
						end

						5'hf: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0) || (r_sys_subRoutine_step==3'h1) || (r_sys_subRoutine_step==3'h2)) begin
										r_sys_tmp2_int <= w_sys_tmp89;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				3'h3: begin

					case(r_sys_subRoutine_phase) 
						5'h8: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0) || (r_sys_subRoutine_step==3'h1) || (r_sys_subRoutine_step==3'h2)) begin
										r_sys_tmp3_int <= w_sys_tmp111;

									end
								end

							endcase
						end

						5'hf: begin

							case(r_sys_subRoutine_stage) 
								2'h0: begin
									if((r_sys_subRoutine_step==3'h0) || (r_sys_subRoutine_step==3'h1) || (r_sys_subRoutine_step==3'h2)) begin
										r_sys_tmp3_int <= w_sys_tmp90;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
