/*
TimeStamp:	2016/9/6		15:33
*/


module c1(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy	
);

	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 6:0] r_sys_run_phase;
	reg         [ 2:0] r_sys_run_stage;
	reg         [ 4:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 2:0] w_sys_run_stage_p1;
	wire        [ 4:0] w_sys_run_step_p1;
	wire signed [14:0] w_fld_u_0_addr_0;
	wire        [31:0] w_fld_u_0_datain_0;
	wire        [31:0] w_fld_u_0_dataout_0;
	wire               w_fld_u_0_r_w_0;
	wire               w_fld_u_0_ce_0;
	reg  signed [14:0] r_fld_u_0_addr_1;
	reg         [31:0] r_fld_u_0_datain_1;
	wire        [31:0] w_fld_u_0_dataout_1;
	reg                r_fld_u_0_r_w_1;
	wire               w_fld_u_0_ce_1;
	wire signed [14:0] w_fld_uu_1_addr_0;
	wire        [31:0] w_fld_uu_1_datain_0;
	wire        [31:0] w_fld_uu_1_dataout_0;
	wire               w_fld_uu_1_r_w_0;
	wire               w_fld_uu_1_ce_0;
	reg  signed [14:0] r_fld_uu_1_addr_1;
	reg         [31:0] r_fld_uu_1_datain_1;
	wire        [31:0] w_fld_uu_1_dataout_1;
	reg                r_fld_uu_1_r_w_1;
	wire               w_fld_uu_1_ce_1;
	wire signed [14:0] w_fld_q_2_addr_0;
	wire        [31:0] w_fld_q_2_datain_0;
	wire        [31:0] w_fld_q_2_dataout_0;
	wire               w_fld_q_2_r_w_0;
	wire               w_fld_q_2_ce_0;
	reg  signed [14:0] r_fld_q_2_addr_1;
	reg         [31:0] r_fld_q_2_datain_1;
	wire        [31:0] w_fld_q_2_dataout_1;
	reg                r_fld_q_2_r_w_1;
	wire               w_fld_q_2_ce_1;
	reg  signed [31:0] r_run_k_7;
	reg  signed [31:0] r_run_j_8;
	reg  signed [31:0] r_run_n_9;
	reg  signed [31:0] r_run_mx_10;
	reg  signed [31:0] r_run_my_11;
	reg  signed [31:0] r_run_nlast_12;
	reg         [31:0] r_run_dx_13;
	reg         [31:0] r_run_dy_14;
	reg         [31:0] r_run_r1_15;
	reg         [31:0] r_run_r2_16;
	reg         [31:0] r_run_dt_17;
	reg  signed [31:0] r_run_copy0_j_18;
	reg  signed [31:0] r_run_copy0_j_19;
	reg  signed [31:0] r_run_copy1_j_20;
	reg  signed [31:0] r_run_copy2_j_21;
	reg  signed [31:0] r_run_copy0_j_22;
	reg  signed [31:0] r_run_copy0_j_23;
	reg  signed [31:0] r_run_copy0_j_24;
	reg  signed [31:0] r_run_copy0_j_25;
	reg  signed [31:0] r_run_copy0_j_26;
	reg  signed [31:0] r_run_copy0_j_27;
	reg  signed [31:0] r_run_copy0_j_28;
	reg  signed [31:0] r_run_copy0_j_29;
	reg                r_sub03_run_req;
	wire               w_sub03_run_busy;
	wire signed [14:0] w_sub03_u_addr;
	reg  signed [14:0] r_sub03_u_addr;
	wire        [31:0] w_sub03_u_datain;
	reg         [31:0] r_sub03_u_datain;
	wire        [31:0] w_sub03_u_dataout;
	wire               w_sub03_u_r_w;
	reg                r_sub03_u_r_w;
	wire signed [14:0] w_sub03_q_addr;
	reg  signed [14:0] r_sub03_q_addr;
	wire        [31:0] w_sub03_q_datain;
	reg         [31:0] r_sub03_q_datain;
	wire        [31:0] w_sub03_q_dataout;
	wire               w_sub03_q_r_w;
	reg                r_sub03_q_r_w;
	wire signed [14:0] w_sub03_result_addr;
	reg  signed [14:0] r_sub03_result_addr;
	wire        [31:0] w_sub03_result_datain;
	reg         [31:0] r_sub03_result_datain;
	wire        [31:0] w_sub03_result_dataout;
	wire               w_sub03_result_r_w;
	reg                r_sub03_result_r_w;
	reg                r_sub02_run_req;
	wire               w_sub02_run_busy;
	wire signed [14:0] w_sub02_u_addr;
	reg  signed [14:0] r_sub02_u_addr;
	wire        [31:0] w_sub02_u_datain;
	reg         [31:0] r_sub02_u_datain;
	wire        [31:0] w_sub02_u_dataout;
	wire               w_sub02_u_r_w;
	reg                r_sub02_u_r_w;
	wire signed [14:0] w_sub02_q_addr;
	reg  signed [14:0] r_sub02_q_addr;
	wire        [31:0] w_sub02_q_datain;
	reg         [31:0] r_sub02_q_datain;
	wire        [31:0] w_sub02_q_dataout;
	wire               w_sub02_q_r_w;
	reg                r_sub02_q_r_w;
	wire signed [14:0] w_sub02_result_addr;
	reg  signed [14:0] r_sub02_result_addr;
	wire        [31:0] w_sub02_result_datain;
	reg         [31:0] r_sub02_result_datain;
	wire        [31:0] w_sub02_result_dataout;
	wire               w_sub02_result_r_w;
	reg                r_sub02_result_r_w;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [14:0] w_sub01_u_addr;
	reg  signed [14:0] r_sub01_u_addr;
	wire        [31:0] w_sub01_u_datain;
	reg         [31:0] r_sub01_u_datain;
	wire        [31:0] w_sub01_u_dataout;
	wire               w_sub01_u_r_w;
	reg                r_sub01_u_r_w;
	wire signed [14:0] w_sub01_q_addr;
	reg  signed [14:0] r_sub01_q_addr;
	wire        [31:0] w_sub01_q_datain;
	reg         [31:0] r_sub01_q_datain;
	wire        [31:0] w_sub01_q_dataout;
	wire               w_sub01_q_r_w;
	reg                r_sub01_q_r_w;
	wire signed [14:0] w_sub01_result_addr;
	reg  signed [14:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [14:0] w_sub00_u_addr;
	reg  signed [14:0] r_sub00_u_addr;
	wire        [31:0] w_sub00_u_datain;
	reg         [31:0] r_sub00_u_datain;
	wire        [31:0] w_sub00_u_dataout;
	wire               w_sub00_u_r_w;
	reg                r_sub00_u_r_w;
	wire signed [14:0] w_sub00_q_addr;
	reg  signed [14:0] r_sub00_q_addr;
	wire        [31:0] w_sub00_q_datain;
	reg         [31:0] r_sub00_q_datain;
	wire        [31:0] w_sub00_q_dataout;
	wire               w_sub00_q_r_w;
	reg                r_sub00_q_r_w;
	wire signed [14:0] w_sub00_result_addr;
	reg  signed [14:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	wire signed [31:0] w_sys_tmp1;
	wire        [31:0] w_sys_tmp3;
	wire        [31:0] w_sys_tmp4;
	wire        [31:0] w_sys_tmp6;
	wire               w_sys_tmp8;
	wire               w_sys_tmp9;
	wire signed [31:0] w_sys_tmp10;
	wire               w_sys_tmp11;
	wire               w_sys_tmp12;
	wire signed [31:0] w_sys_tmp15;
	wire signed [31:0] w_sys_tmp16;
	wire signed [31:0] w_sys_tmp17;
	wire        [31:0] w_sys_tmp18;
	wire signed [31:0] w_sys_tmp20;
	wire signed [31:0] w_sys_tmp21;
	wire signed [31:0] w_sys_tmp24;
	wire signed [31:0] w_sys_tmp25;
	wire               w_sys_tmp98;
	wire               w_sys_tmp99;
	wire signed [31:0] w_sys_tmp100;
	wire               w_sys_tmp101;
	wire               w_sys_tmp102;
	wire signed [31:0] w_sys_tmp105;
	wire signed [31:0] w_sys_tmp106;
	wire        [31:0] w_sys_tmp107;
	wire signed [31:0] w_sys_tmp109;
	wire signed [31:0] w_sys_tmp110;
	wire        [31:0] w_sys_tmp112;
	wire signed [31:0] w_sys_tmp114;
	wire signed [31:0] w_sys_tmp115;
	wire        [31:0] w_sys_tmp117;
	wire signed [31:0] w_sys_tmp119;
	wire signed [31:0] w_sys_tmp120;
	wire signed [31:0] w_sys_tmp123;
	wire signed [31:0] w_sys_tmp124;
	wire signed [31:0] w_sys_tmp125;
	wire signed [31:0] w_sys_tmp126;
	wire               w_sys_tmp265;
	wire               w_sys_tmp266;
	wire signed [31:0] w_sys_tmp267;
	wire signed [31:0] w_sys_tmp268;
	wire               w_sys_tmp269;
	wire               w_sys_tmp270;
	wire signed [31:0] w_sys_tmp271;
	wire signed [31:0] w_sys_tmp274;
	wire signed [31:0] w_sys_tmp275;
	wire signed [31:0] w_sys_tmp276;
	wire        [31:0] w_sys_tmp277;
	wire signed [31:0] w_sys_tmp278;
	wire signed [31:0] w_sys_tmp279;
	wire signed [31:0] w_sys_tmp281;
	wire signed [31:0] w_sys_tmp282;
	wire signed [31:0] w_sys_tmp343;
	wire               w_sys_tmp344;
	wire               w_sys_tmp345;
	wire signed [31:0] w_sys_tmp346;
	wire signed [31:0] w_sys_tmp349;
	wire signed [31:0] w_sys_tmp350;
	wire signed [31:0] w_sys_tmp351;
	wire        [31:0] w_sys_tmp352;
	wire signed [31:0] w_sys_tmp353;
	wire signed [31:0] w_sys_tmp354;
	wire signed [31:0] w_sys_tmp356;
	wire signed [31:0] w_sys_tmp357;
	wire signed [31:0] w_sys_tmp418;
	wire               w_sys_tmp419;
	wire               w_sys_tmp420;
	wire signed [31:0] w_sys_tmp421;
	wire signed [31:0] w_sys_tmp422;
	wire               w_sys_tmp423;
	wire               w_sys_tmp424;
	wire signed [31:0] w_sys_tmp425;
	wire signed [31:0] w_sys_tmp428;
	wire signed [31:0] w_sys_tmp429;
	wire signed [31:0] w_sys_tmp430;
	wire        [31:0] w_sys_tmp431;
	wire signed [31:0] w_sys_tmp432;
	wire signed [31:0] w_sys_tmp433;
	wire signed [31:0] w_sys_tmp435;
	wire signed [31:0] w_sys_tmp436;
	wire signed [31:0] w_sys_tmp497;
	wire               w_sys_tmp498;
	wire               w_sys_tmp499;
	wire signed [31:0] w_sys_tmp500;
	wire signed [31:0] w_sys_tmp503;
	wire signed [31:0] w_sys_tmp504;
	wire signed [31:0] w_sys_tmp505;
	wire        [31:0] w_sys_tmp506;
	wire signed [31:0] w_sys_tmp507;
	wire signed [31:0] w_sys_tmp508;
	wire signed [31:0] w_sys_tmp510;
	wire signed [31:0] w_sys_tmp511;
	wire signed [31:0] w_sys_tmp572;
	wire               w_sys_tmp573;
	wire               w_sys_tmp574;
	wire signed [31:0] w_sys_tmp575;
	wire signed [31:0] w_sys_tmp576;
	wire signed [31:0] w_sys_tmp577;
	wire               w_sys_tmp578;
	wire               w_sys_tmp579;
	wire signed [31:0] w_sys_tmp580;
	wire signed [31:0] w_sys_tmp583;
	wire signed [31:0] w_sys_tmp584;
	wire signed [31:0] w_sys_tmp585;
	wire        [31:0] w_sys_tmp586;
	wire signed [31:0] w_sys_tmp587;
	wire signed [31:0] w_sys_tmp588;
	wire signed [31:0] w_sys_tmp590;
	wire signed [31:0] w_sys_tmp591;
	wire signed [31:0] w_sys_tmp652;
	wire               w_sys_tmp653;
	wire               w_sys_tmp654;
	wire signed [31:0] w_sys_tmp655;
	wire signed [31:0] w_sys_tmp658;
	wire signed [31:0] w_sys_tmp659;
	wire signed [31:0] w_sys_tmp660;
	wire        [31:0] w_sys_tmp661;
	wire signed [31:0] w_sys_tmp662;
	wire signed [31:0] w_sys_tmp663;
	wire signed [31:0] w_sys_tmp665;
	wire signed [31:0] w_sys_tmp666;
	wire signed [31:0] w_sys_tmp727;
	wire               w_sys_tmp728;
	wire               w_sys_tmp729;
	wire signed [31:0] w_sys_tmp730;
	wire signed [31:0] w_sys_tmp731;
	wire signed [31:0] w_sys_tmp732;
	wire               w_sys_tmp733;
	wire               w_sys_tmp734;
	wire signed [31:0] w_sys_tmp735;
	wire signed [31:0] w_sys_tmp738;
	wire signed [31:0] w_sys_tmp739;
	wire signed [31:0] w_sys_tmp740;
	wire        [31:0] w_sys_tmp741;
	wire signed [31:0] w_sys_tmp742;
	wire signed [31:0] w_sys_tmp743;
	wire signed [31:0] w_sys_tmp745;
	wire signed [31:0] w_sys_tmp746;
	wire signed [31:0] w_sys_tmp807;
	wire               w_sys_tmp808;
	wire               w_sys_tmp809;
	wire signed [31:0] w_sys_tmp810;
	wire signed [31:0] w_sys_tmp813;
	wire signed [31:0] w_sys_tmp814;
	wire signed [31:0] w_sys_tmp815;
	wire        [31:0] w_sys_tmp816;
	wire signed [31:0] w_sys_tmp817;
	wire signed [31:0] w_sys_tmp818;
	wire signed [31:0] w_sys_tmp820;
	wire signed [31:0] w_sys_tmp821;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 3'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 5'h1);
	assign w_fld_u_0_addr_0 = 15'sh0;
	assign w_fld_u_0_datain_0 = 32'h0;
	assign w_fld_u_0_r_w_0 = 1'h0;
	assign w_fld_u_0_ce_0 = w_sys_ce;
	assign w_fld_u_0_ce_1 = w_sys_ce;
	assign w_fld_uu_1_addr_0 = 15'sh0;
	assign w_fld_uu_1_datain_0 = 32'h0;
	assign w_fld_uu_1_r_w_0 = 1'h0;
	assign w_fld_uu_1_ce_0 = w_sys_ce;
	assign w_fld_uu_1_ce_1 = w_sys_ce;
	assign w_fld_q_2_addr_0 = 15'sh0;
	assign w_fld_q_2_datain_0 = 32'h0;
	assign w_fld_q_2_r_w_0 = 1'h0;
	assign w_fld_q_2_ce_0 = w_sys_ce;
	assign w_fld_q_2_ce_1 = w_sys_ce;
	assign w_sub03_u_addr = ( (|r_sys_processing_methodID) ? r_sub03_u_addr : 15'sh0 ) ;
	assign w_sub03_u_datain = ( (|r_sys_processing_methodID) ? r_sub03_u_datain : 32'h0 ) ;
	assign w_sub03_u_r_w = ( (|r_sys_processing_methodID) ? r_sub03_u_r_w : 1'h0 ) ;
	assign w_sub03_q_addr = ( (|r_sys_processing_methodID) ? r_sub03_q_addr : 15'sh0 ) ;
	assign w_sub03_q_datain = ( (|r_sys_processing_methodID) ? r_sub03_q_datain : 32'h0 ) ;
	assign w_sub03_q_r_w = ( (|r_sys_processing_methodID) ? r_sub03_q_r_w : 1'h0 ) ;
	assign w_sub03_result_addr = ( (|r_sys_processing_methodID) ? r_sub03_result_addr : 15'sh0 ) ;
	assign w_sub03_result_datain = ( (|r_sys_processing_methodID) ? r_sub03_result_datain : 32'h0 ) ;
	assign w_sub03_result_r_w = ( (|r_sys_processing_methodID) ? r_sub03_result_r_w : 1'h0 ) ;
	assign w_sub02_u_addr = ( (|r_sys_processing_methodID) ? r_sub02_u_addr : 15'sh0 ) ;
	assign w_sub02_u_datain = ( (|r_sys_processing_methodID) ? r_sub02_u_datain : 32'h0 ) ;
	assign w_sub02_u_r_w = ( (|r_sys_processing_methodID) ? r_sub02_u_r_w : 1'h0 ) ;
	assign w_sub02_q_addr = ( (|r_sys_processing_methodID) ? r_sub02_q_addr : 15'sh0 ) ;
	assign w_sub02_q_datain = ( (|r_sys_processing_methodID) ? r_sub02_q_datain : 32'h0 ) ;
	assign w_sub02_q_r_w = ( (|r_sys_processing_methodID) ? r_sub02_q_r_w : 1'h0 ) ;
	assign w_sub02_result_addr = ( (|r_sys_processing_methodID) ? r_sub02_result_addr : 15'sh0 ) ;
	assign w_sub02_result_datain = ( (|r_sys_processing_methodID) ? r_sub02_result_datain : 32'h0 ) ;
	assign w_sub02_result_r_w = ( (|r_sys_processing_methodID) ? r_sub02_result_r_w : 1'h0 ) ;
	assign w_sub01_u_addr = ( (|r_sys_processing_methodID) ? r_sub01_u_addr : 15'sh0 ) ;
	assign w_sub01_u_datain = ( (|r_sys_processing_methodID) ? r_sub01_u_datain : 32'h0 ) ;
	assign w_sub01_u_r_w = ( (|r_sys_processing_methodID) ? r_sub01_u_r_w : 1'h0 ) ;
	assign w_sub01_q_addr = ( (|r_sys_processing_methodID) ? r_sub01_q_addr : 15'sh0 ) ;
	assign w_sub01_q_datain = ( (|r_sys_processing_methodID) ? r_sub01_q_datain : 32'h0 ) ;
	assign w_sub01_q_r_w = ( (|r_sys_processing_methodID) ? r_sub01_q_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 15'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub00_u_addr = ( (|r_sys_processing_methodID) ? r_sub00_u_addr : 15'sh0 ) ;
	assign w_sub00_u_datain = ( (|r_sys_processing_methodID) ? r_sub00_u_datain : 32'h0 ) ;
	assign w_sub00_u_r_w = ( (|r_sys_processing_methodID) ? r_sub00_u_r_w : 1'h0 ) ;
	assign w_sub00_q_addr = ( (|r_sys_processing_methodID) ? r_sub00_q_addr : 15'sh0 ) ;
	assign w_sub00_q_datain = ( (|r_sys_processing_methodID) ? r_sub00_q_datain : 32'h0 ) ;
	assign w_sub00_q_r_w = ( (|r_sys_processing_methodID) ? r_sub00_q_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 15'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh00000081;
	assign w_sys_tmp3 = 32'h3a03126f;
	assign w_sys_tmp4 = 32'h3c000000;
	assign w_sys_tmp6 = 32'h4103126f;
	assign w_sys_tmp8 = ( !w_sys_tmp9 );
	assign w_sys_tmp9 = (r_run_my_11 < r_run_k_7);
	assign w_sys_tmp10 = (r_run_k_7 + w_sys_intOne);
	assign w_sys_tmp11 = ( !w_sys_tmp12 );
	assign w_sys_tmp12 = (r_run_mx_10 < r_run_j_8);
	assign w_sys_tmp15 = (w_sys_tmp16 + r_run_k_7);
	assign w_sys_tmp16 = (r_run_j_8 * w_sys_tmp17);
	assign w_sys_tmp17 = 32'sh00000081;
	assign w_sys_tmp18 = 32'h0;
	assign w_sys_tmp20 = (w_sys_tmp21 + r_run_k_7);
	assign w_sys_tmp21 = (r_run_copy0_j_18 * w_sys_tmp17);
	assign w_sys_tmp24 = (r_run_copy0_j_18 + w_sys_intOne);
	assign w_sys_tmp25 = (r_run_j_8 + w_sys_intOne);
	assign w_sys_tmp98 = ( !w_sys_tmp99 );
	assign w_sys_tmp99 = (r_run_nlast_12 < r_run_n_9);
	assign w_sys_tmp100 = (r_run_n_9 + w_sys_intOne);
	assign w_sys_tmp101 = ( !w_sys_tmp102 );
	assign w_sys_tmp102 = (r_run_my_11 < r_run_j_8);
	assign w_sys_tmp105 = (w_sys_tmp106 + r_run_j_8);
	assign w_sys_tmp106 = 32'sh00000081;
	assign w_sys_tmp107 = 32'h3f000000;
	assign w_sys_tmp109 = (w_sys_tmp110 + r_run_copy2_j_21);
	assign w_sys_tmp110 = (r_run_mx_10 * w_sys_tmp106);
	assign w_sys_tmp112 = 32'h0;
	assign w_sys_tmp114 = (w_sys_tmp115 + w_sys_intOne);
	assign w_sys_tmp115 = (r_run_copy1_j_20 * w_sys_tmp106);
	assign w_sys_tmp117 = 32'h3f800000;
	assign w_sys_tmp119 = (w_sys_tmp120 + r_run_my_11);
	assign w_sys_tmp120 = (r_run_copy0_j_19 * w_sys_tmp106);
	assign w_sys_tmp123 = (r_run_copy0_j_19 + w_sys_intOne);
	assign w_sys_tmp124 = (r_run_copy1_j_20 + w_sys_intOne);
	assign w_sys_tmp125 = (r_run_copy2_j_21 + w_sys_intOne);
	assign w_sys_tmp126 = (r_run_j_8 + w_sys_intOne);
	assign w_sys_tmp265 = ( !w_sys_tmp266 );
	assign w_sys_tmp266 = (w_sys_tmp267 < r_run_k_7);
	assign w_sys_tmp267 = 32'sh00000041;
	assign w_sys_tmp268 = (r_run_k_7 + w_sys_intOne);
	assign w_sys_tmp269 = ( !w_sys_tmp270 );
	assign w_sys_tmp270 = (w_sys_tmp271 < r_run_j_8);
	assign w_sys_tmp271 = 32'sh00000041;
	assign w_sys_tmp274 = (w_sys_tmp275 + r_run_k_7);
	assign w_sys_tmp275 = (r_run_j_8 * w_sys_tmp276);
	assign w_sys_tmp276 = 32'sh00000081;
	assign w_sys_tmp277 = w_fld_u_0_dataout_1;
	assign w_sys_tmp278 = (w_sys_tmp279 + r_run_k_7);
	assign w_sys_tmp279 = (r_run_copy0_j_22 * w_sys_tmp276);
	assign w_sys_tmp281 = (r_run_copy0_j_22 + w_sys_intOne);
	assign w_sys_tmp282 = (r_run_j_8 + w_sys_intOne);
	assign w_sys_tmp343 = 32'sh00000041;
	assign w_sys_tmp344 = ( !w_sys_tmp345 );
	assign w_sys_tmp345 = (w_sys_tmp346 < r_run_j_8);
	assign w_sys_tmp346 = 32'sh00000081;
	assign w_sys_tmp349 = (w_sys_tmp350 + r_run_k_7);
	assign w_sys_tmp350 = (r_run_j_8 * w_sys_tmp351);
	assign w_sys_tmp351 = 32'sh00000081;
	assign w_sys_tmp352 = w_fld_u_0_dataout_1;
	assign w_sys_tmp353 = (w_sys_tmp354 + r_run_k_7);
	assign w_sys_tmp354 = (r_run_copy0_j_23 * w_sys_tmp351);
	assign w_sys_tmp356 = (r_run_copy0_j_23 + w_sys_intOne);
	assign w_sys_tmp357 = (r_run_j_8 + w_sys_intOne);
	assign w_sys_tmp418 = 32'sh00000040;
	assign w_sys_tmp419 = ( !w_sys_tmp420 );
	assign w_sys_tmp420 = (w_sys_tmp421 < r_run_k_7);
	assign w_sys_tmp421 = 32'sh00000081;
	assign w_sys_tmp422 = (r_run_k_7 + w_sys_intOne);
	assign w_sys_tmp423 = ( !w_sys_tmp424 );
	assign w_sys_tmp424 = (w_sys_tmp425 < r_run_j_8);
	assign w_sys_tmp425 = 32'sh00000041;
	assign w_sys_tmp428 = (w_sys_tmp429 + r_run_k_7);
	assign w_sys_tmp429 = (r_run_j_8 * w_sys_tmp430);
	assign w_sys_tmp430 = 32'sh00000081;
	assign w_sys_tmp431 = w_fld_u_0_dataout_1;
	assign w_sys_tmp432 = (w_sys_tmp433 + r_run_k_7);
	assign w_sys_tmp433 = (r_run_copy0_j_24 * w_sys_tmp430);
	assign w_sys_tmp435 = (r_run_copy0_j_24 + w_sys_intOne);
	assign w_sys_tmp436 = (r_run_j_8 + w_sys_intOne);
	assign w_sys_tmp497 = 32'sh00000041;
	assign w_sys_tmp498 = ( !w_sys_tmp499 );
	assign w_sys_tmp499 = (w_sys_tmp500 < r_run_j_8);
	assign w_sys_tmp500 = 32'sh00000081;
	assign w_sys_tmp503 = (w_sys_tmp504 + r_run_k_7);
	assign w_sys_tmp504 = (r_run_j_8 * w_sys_tmp505);
	assign w_sys_tmp505 = 32'sh00000081;
	assign w_sys_tmp506 = w_fld_u_0_dataout_1;
	assign w_sys_tmp507 = (w_sys_tmp508 + r_run_k_7);
	assign w_sys_tmp508 = (r_run_copy0_j_25 * w_sys_tmp505);
	assign w_sys_tmp510 = (r_run_copy0_j_25 + w_sys_intOne);
	assign w_sys_tmp511 = (r_run_j_8 + w_sys_intOne);
	assign w_sys_tmp572 = 32'sh00000002;
	assign w_sys_tmp573 = ( !w_sys_tmp574 );
	assign w_sys_tmp574 = (w_sys_tmp575 < r_run_k_7);
	assign w_sys_tmp575 = 32'sh00000040;
	assign w_sys_tmp576 = (r_run_k_7 + w_sys_intOne);
	assign w_sys_tmp577 = 32'sh00000002;
	assign w_sys_tmp578 = ( !w_sys_tmp579 );
	assign w_sys_tmp579 = (w_sys_tmp580 < r_run_j_8);
	assign w_sys_tmp580 = 32'sh00000040;
	assign w_sys_tmp583 = (w_sys_tmp584 + r_run_k_7);
	assign w_sys_tmp584 = (r_run_j_8 * w_sys_tmp585);
	assign w_sys_tmp585 = 32'sh00000081;
	assign w_sys_tmp586 = w_sub00_result_dataout;
	assign w_sys_tmp587 = (w_sys_tmp588 + r_run_k_7);
	assign w_sys_tmp588 = (r_run_copy0_j_26 * w_sys_tmp585);
	assign w_sys_tmp590 = (r_run_copy0_j_26 + w_sys_intOne);
	assign w_sys_tmp591 = (r_run_j_8 + w_sys_intOne);
	assign w_sys_tmp652 = 32'sh00000041;
	assign w_sys_tmp653 = ( !w_sys_tmp654 );
	assign w_sys_tmp654 = (w_sys_tmp655 < r_run_j_8);
	assign w_sys_tmp655 = 32'sh00000080;
	assign w_sys_tmp658 = (w_sys_tmp659 + r_run_k_7);
	assign w_sys_tmp659 = (r_run_j_8 * w_sys_tmp660);
	assign w_sys_tmp660 = 32'sh00000081;
	assign w_sys_tmp661 = w_sub01_result_dataout;
	assign w_sys_tmp662 = (w_sys_tmp663 + r_run_k_7);
	assign w_sys_tmp663 = (r_run_copy0_j_27 * w_sys_tmp660);
	assign w_sys_tmp665 = (r_run_copy0_j_27 + w_sys_intOne);
	assign w_sys_tmp666 = (r_run_j_8 + w_sys_intOne);
	assign w_sys_tmp727 = 32'sh00000041;
	assign w_sys_tmp728 = ( !w_sys_tmp729 );
	assign w_sys_tmp729 = (w_sys_tmp730 < r_run_k_7);
	assign w_sys_tmp730 = 32'sh00000080;
	assign w_sys_tmp731 = (r_run_k_7 + w_sys_intOne);
	assign w_sys_tmp732 = 32'sh00000002;
	assign w_sys_tmp733 = ( !w_sys_tmp734 );
	assign w_sys_tmp734 = (w_sys_tmp735 < r_run_j_8);
	assign w_sys_tmp735 = 32'sh00000040;
	assign w_sys_tmp738 = (w_sys_tmp739 + r_run_k_7);
	assign w_sys_tmp739 = (r_run_j_8 * w_sys_tmp740);
	assign w_sys_tmp740 = 32'sh00000081;
	assign w_sys_tmp741 = w_sub02_result_dataout;
	assign w_sys_tmp742 = (w_sys_tmp743 + r_run_k_7);
	assign w_sys_tmp743 = (r_run_copy0_j_28 * w_sys_tmp740);
	assign w_sys_tmp745 = (r_run_copy0_j_28 + w_sys_intOne);
	assign w_sys_tmp746 = (r_run_j_8 + w_sys_intOne);
	assign w_sys_tmp807 = 32'sh00000041;
	assign w_sys_tmp808 = ( !w_sys_tmp809 );
	assign w_sys_tmp809 = (w_sys_tmp810 < r_run_j_8);
	assign w_sys_tmp810 = 32'sh00000080;
	assign w_sys_tmp813 = (w_sys_tmp814 + r_run_k_7);
	assign w_sys_tmp814 = (r_run_j_8 * w_sys_tmp815);
	assign w_sys_tmp815 = 32'sh00000081;
	assign w_sys_tmp816 = w_sub03_result_dataout;
	assign w_sys_tmp817 = (w_sys_tmp818 + r_run_k_7);
	assign w_sys_tmp818 = (r_run_copy0_j_29 * w_sys_tmp815);
	assign w_sys_tmp820 = (r_run_copy0_j_29 + w_sys_intOne);
	assign w_sys_tmp821 = (r_run_j_8 + w_sys_intOne);


	sub03
		sub03_inst(
			.i_fld_q_1_addr_0 (w_sub03_q_addr),
			.i_fld_q_1_datain_0 (w_sub03_q_datain),
			.o_fld_q_1_dataout_0 (w_sub03_q_dataout),
			.i_fld_q_1_r_w_0 (w_sub03_q_r_w),
			.i_fld_result_2_addr_0 (w_sub03_result_addr),
			.i_fld_result_2_datain_0 (w_sub03_result_datain),
			.o_fld_result_2_dataout_0 (w_sub03_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub03_result_r_w),
			.i_fld_u_0_addr_0 (w_sub03_u_addr),
			.i_fld_u_0_datain_0 (w_sub03_u_datain),
			.o_fld_u_0_dataout_0 (w_sub03_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub03_u_r_w),
			.o_run_busy (w_sub03_run_busy),
			.i_run_req (r_sub03_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub02
		sub02_inst(
			.i_fld_q_1_addr_0 (w_sub02_q_addr),
			.i_fld_q_1_datain_0 (w_sub02_q_datain),
			.o_fld_q_1_dataout_0 (w_sub02_q_dataout),
			.i_fld_q_1_r_w_0 (w_sub02_q_r_w),
			.i_fld_result_2_addr_0 (w_sub02_result_addr),
			.i_fld_result_2_datain_0 (w_sub02_result_datain),
			.o_fld_result_2_dataout_0 (w_sub02_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub02_result_r_w),
			.i_fld_u_0_addr_0 (w_sub02_u_addr),
			.i_fld_u_0_datain_0 (w_sub02_u_datain),
			.o_fld_u_0_dataout_0 (w_sub02_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub02_u_r_w),
			.o_run_busy (w_sub02_run_busy),
			.i_run_req (r_sub02_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub01
		sub01_inst(
			.i_fld_q_1_addr_0 (w_sub01_q_addr),
			.i_fld_q_1_datain_0 (w_sub01_q_datain),
			.o_fld_q_1_dataout_0 (w_sub01_q_dataout),
			.i_fld_q_1_r_w_0 (w_sub01_q_r_w),
			.i_fld_result_2_addr_0 (w_sub01_result_addr),
			.i_fld_result_2_datain_0 (w_sub01_result_datain),
			.o_fld_result_2_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub01_result_r_w),
			.i_fld_u_0_addr_0 (w_sub01_u_addr),
			.i_fld_u_0_datain_0 (w_sub01_u_datain),
			.o_fld_u_0_dataout_0 (w_sub01_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub01_u_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub00
		sub00_inst(
			.i_fld_q_1_addr_0 (w_sub00_q_addr),
			.i_fld_q_1_datain_0 (w_sub00_q_datain),
			.o_fld_q_1_dataout_0 (w_sub00_q_dataout),
			.i_fld_q_1_r_w_0 (w_sub00_q_r_w),
			.i_fld_result_2_addr_0 (w_sub00_result_addr),
			.i_fld_result_2_datain_0 (w_sub00_result_datain),
			.o_fld_result_2_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_2_r_w_0 (w_sub00_result_r_w),
			.i_fld_u_0_addr_0 (w_sub00_u_addr),
			.i_fld_u_0_datain_0 (w_sub00_u_datain),
			.o_fld_u_0_dataout_0 (w_sub00_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub00_u_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_u_0(
			.clk (clock),
			.ce_0 (w_fld_u_0_ce_0),
			.addr_0 (w_fld_u_0_addr_0),
			.datain_0 (w_fld_u_0_datain_0),
			.dataout_0 (w_fld_u_0_dataout_0),
			.r_w_0 (w_fld_u_0_r_w_0),
			.ce_1 (w_fld_u_0_ce_1),
			.addr_1 (r_fld_u_0_addr_1),
			.datain_1 (r_fld_u_0_datain_1),
			.dataout_1 (w_fld_u_0_dataout_1),
			.r_w_1 (r_fld_u_0_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_uu_1(
			.clk (clock),
			.ce_0 (w_fld_uu_1_ce_0),
			.addr_0 (w_fld_uu_1_addr_0),
			.datain_0 (w_fld_uu_1_datain_0),
			.dataout_0 (w_fld_uu_1_dataout_0),
			.r_w_0 (w_fld_uu_1_r_w_0),
			.ce_1 (w_fld_uu_1_ce_1),
			.addr_1 (r_fld_uu_1_addr_1),
			.datain_1 (r_fld_uu_1_datain_1),
			.dataout_1 (w_fld_uu_1_dataout_1),
			.r_w_1 (r_fld_uu_1_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_q_2(
			.clk (clock),
			.ce_0 (w_fld_q_2_ce_0),
			.addr_0 (w_fld_q_2_addr_0),
			.datain_0 (w_fld_q_2_datain_0),
			.dataout_0 (w_fld_q_2_dataout_0),
			.r_w_0 (w_fld_q_2_r_w_0),
			.ce_1 (w_fld_q_2_ce_1),
			.addr_1 (r_fld_q_2_addr_1),
			.datain_1 (r_fld_q_2_datain_1),
			.dataout_1 (w_fld_q_2_dataout_1),
			.r_w_1 (r_fld_q_2_r_w_1)
		);

	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						7'h61: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 7'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h0: begin
							r_sys_run_phase <= 7'h2;
						end

						7'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h4;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h5;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp8) ? 7'h9 : 7'hf);

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h5;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'ha;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp11) ? 7'hd : 7'h6);

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h6)) begin
										r_sys_run_phase <= 7'ha;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h10;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp98) ? 7'h14 : 7'h61);

									end
								end

							endcase
						end

						7'h11: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h10;

									end
								end

							endcase
						end

						7'h14: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h15;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp101) ? 7'h18 : 7'h1a);

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1b)) begin
										r_sys_run_phase <= 7'h15;

									end
								end

							endcase
						end

						7'h1a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h1b;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp265) ? 7'h1f : 7'h2b);

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h1b;

									end
								end

							endcase
						end

						7'h1f: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h20;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp269) ? 7'h23 : 7'h25);

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 7'h20;

									end
								end

							endcase
						end

						7'h25: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h26;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp344) ? 7'h29 : 7'h1c);

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 7'h26;

									end
								end

							endcase
						end

						7'h2b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h2c;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp419) ? 7'h30 : 7'h3b);

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h2c;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h31;

									end
								end

							endcase
						end

						7'h31: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp423) ? 7'h34 : 7'h36);

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 7'h31;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h37;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp498) ? 7'h3a : 7'h2d);

									end
								end

							endcase
						end

						7'h3a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 7'h37;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								3'h3: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_phase <= 7'h3d;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								3'h3: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_phase <= 7'h3f;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h40;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp573) ? 7'h44 : 7'h50);

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h40;

									end
								end

							endcase
						end

						7'h44: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h45;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp578) ? 7'h48 : 7'h4a);

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 7'h45;

									end
								end

							endcase
						end

						7'h4a: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h4b;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp653) ? 7'h4e : 7'h41);

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 7'h4b;

									end
								end

							endcase
						end

						7'h50: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h51;

									end
								end

							endcase
						end

						7'h51: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp728) ? 7'h55 : 7'h11);

									end
								end

							endcase
						end

						7'h52: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h51;

									end
								end

							endcase
						end

						7'h55: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h56;

									end
								end

							endcase
						end

						7'h56: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp733) ? 7'h59 : 7'h5b);

									end
								end

							endcase
						end

						7'h59: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 7'h56;

									end
								end

							endcase
						end

						7'h5b: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 7'h5c;

									end
								end

							endcase
						end

						7'h5c: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp808) ? 7'h5f : 7'h52);

									end
								end

							endcase
						end

						7'h5f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_phase <= 7'h5c;

									end
								end

							endcase
						end

						7'h61: begin
							r_sys_run_phase <= 7'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 3'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h6)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h11: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h14: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1b)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h1a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h2b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h31: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h3a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h44: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h4a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h50: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h51: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h52: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h55: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h56: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h59: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h5b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h5c: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						7'h5f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 5'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h6)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h5)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h11: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h14: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1b)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h1a)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h1a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h2b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h31: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h3a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub00_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub01_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub02_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub03_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h44: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h4a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h50: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h51: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h52: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h55: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h56: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h59: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h5b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h5c: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						7'h5f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						7'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						7'h61: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp15[14:0] );

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0) || (r_sys_run_step==5'h4) || (r_sys_run_step==5'h8) || (r_sys_run_step==5'hc) || (r_sys_run_step==5'h10) || (r_sys_run_step==5'h14) || (r_sys_run_step==5'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp105[14:0] );

									end
									else
									if((r_sys_run_step==5'h1) || (r_sys_run_step==5'h5) || (r_sys_run_step==5'h9) || (r_sys_run_step==5'hd) || (r_sys_run_step==5'h11) || (r_sys_run_step==5'h15) || (r_sys_run_step==5'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp109[14:0] );

									end
									else
									if((r_sys_run_step==5'h2) || (r_sys_run_step==5'h6) || (r_sys_run_step==5'ha) || (r_sys_run_step==5'he) || (r_sys_run_step==5'h12) || (r_sys_run_step==5'h16) || (r_sys_run_step==5'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp114[14:0] );

									end
									else
									if((r_sys_run_step==5'h3) || (r_sys_run_step==5'h7) || (r_sys_run_step==5'hb) || (r_sys_run_step==5'hf) || (r_sys_run_step==5'h13) || (r_sys_run_step==5'h17) || (r_sys_run_step==5'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp119[14:0] );

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp278[14:0] );

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp353[14:0] );

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp432[14:0] );

									end
								end

							endcase
						end

						7'h3a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp507[14:0] );

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp583[14:0] );

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp658[14:0] );

									end
								end

							endcase
						end

						7'h59: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp738[14:0] );

									end
								end

							endcase
						end

						7'h5f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp813[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp18;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h2) || (r_sys_run_step==5'h6) || (r_sys_run_step==5'ha) || (r_sys_run_step==5'he) || (r_sys_run_step==5'h12) || (r_sys_run_step==5'h16) || (r_sys_run_step==5'h1a)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp117;

									end
									else
									if((r_sys_run_step==5'h0) || (r_sys_run_step==5'h4) || (r_sys_run_step==5'h8) || (r_sys_run_step==5'hc) || (r_sys_run_step==5'h10) || (r_sys_run_step==5'h14) || (r_sys_run_step==5'h18)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp107;

									end
									else
									if((r_sys_run_step==5'h1) || (r_sys_run_step==5'h3) || (r_sys_run_step==5'h5) || (r_sys_run_step==5'h7) || (r_sys_run_step==5'h9) || (r_sys_run_step==5'hb) || (r_sys_run_step==5'hd) || (r_sys_run_step==5'hf) || (r_sys_run_step==5'h11) || (r_sys_run_step==5'h13) || (r_sys_run_step==5'h15) || (r_sys_run_step==5'h17) || (r_sys_run_step==5'h19) || (r_sys_run_step==5'h1b)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp112;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp586;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp661;

									end
								end

							endcase
						end

						7'h59: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp741;

									end
								end

							endcase
						end

						7'h5f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp816;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h1b)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h59: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h5f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h61: begin
							r_fld_u_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_uu_1_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_uu_1_addr_1 <= $signed( w_sys_tmp20[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_uu_1_datain_1 <= w_sys_tmp18;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_uu_1_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_uu_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h61: begin
							r_fld_uu_1_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_q_2_addr_1 <= 15'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_q_2_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h61: begin
							r_fld_q_2_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_7 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_7 <= w_sys_tmp10;

									end
								end

							endcase
						end

						7'h1a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_7 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_7 <= w_sys_tmp268;

									end
								end

							endcase
						end

						7'h2b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_7 <= w_sys_tmp418;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_7 <= w_sys_tmp422;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_7 <= w_sys_tmp572;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_7 <= w_sys_tmp576;

									end
								end

							endcase
						end

						7'h50: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_7 <= w_sys_tmp727;

									end
								end

							endcase
						end

						7'h52: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_7 <= w_sys_tmp731;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_8 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_j_8 <= w_sys_tmp25;

									end
								end

							endcase
						end

						7'h14: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_8 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0) || (r_sys_run_step==5'h4) || (r_sys_run_step==5'h8) || (r_sys_run_step==5'hc) || (r_sys_run_step==5'h10) || (r_sys_run_step==5'h14) || (r_sys_run_step==5'h18)) begin
										r_run_j_8 <= w_sys_tmp126;

									end
								end

							endcase
						end

						7'h1f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_8 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_8 <= w_sys_tmp282;

									end
								end

							endcase
						end

						7'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_8 <= w_sys_tmp343;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_8 <= w_sys_tmp357;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_8 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_8 <= w_sys_tmp436;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_8 <= w_sys_tmp497;

									end
								end

							endcase
						end

						7'h3a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_8 <= w_sys_tmp511;

									end
								end

							endcase
						end

						7'h44: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_8 <= w_sys_tmp577;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_8 <= w_sys_tmp591;

									end
								end

							endcase
						end

						7'h4a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_8 <= w_sys_tmp652;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_8 <= w_sys_tmp666;

									end
								end

							endcase
						end

						7'h55: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_8 <= w_sys_tmp732;

									end
								end

							endcase
						end

						7'h59: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_8 <= w_sys_tmp746;

									end
								end

							endcase
						end

						7'h5b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_8 <= w_sys_tmp807;

									end
								end

							endcase
						end

						7'h5f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_run_j_8 <= w_sys_tmp821;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hf: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_n_9 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h11: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_n_9 <= w_sys_tmp100;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_mx_10 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_my_11 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_nlast_12 <= w_sys_intOne;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_dx_13 <= w_sys_tmp4;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_dy_14 <= w_sys_tmp4;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_r1_15 <= w_sys_tmp6;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_r2_16 <= w_sys_tmp6;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_dt_17 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_18 <= r_run_j_8;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_18 <= w_sys_tmp24;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h14: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_19 <= r_run_j_8;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h3) || (r_sys_run_step==5'h7) || (r_sys_run_step==5'hb) || (r_sys_run_step==5'hf) || (r_sys_run_step==5'h13) || (r_sys_run_step==5'h17) || (r_sys_run_step==5'h1b)) begin
										r_run_copy0_j_19 <= w_sys_tmp123;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h14: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy1_j_20 <= r_run_j_8;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h2) || (r_sys_run_step==5'h6) || (r_sys_run_step==5'ha) || (r_sys_run_step==5'he) || (r_sys_run_step==5'h12) || (r_sys_run_step==5'h16) || (r_sys_run_step==5'h1a)) begin
										r_run_copy1_j_20 <= w_sys_tmp124;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h14: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy2_j_21 <= r_run_j_8;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1) || (r_sys_run_step==5'h5) || (r_sys_run_step==5'h9) || (r_sys_run_step==5'hd) || (r_sys_run_step==5'h11) || (r_sys_run_step==5'h15) || (r_sys_run_step==5'h19)) begin
										r_run_copy2_j_21 <= w_sys_tmp125;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h1f: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_22 <= r_run_j_8;

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_22 <= w_sys_tmp281;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h25: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_23 <= r_run_j_8;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_23 <= w_sys_tmp356;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h30: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_24 <= r_run_j_8;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_24 <= w_sys_tmp435;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_25 <= r_run_j_8;

									end
								end

							endcase
						end

						7'h3a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_25 <= w_sys_tmp510;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h44: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_26 <= r_run_j_8;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_26 <= w_sys_tmp590;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4a: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_27 <= r_run_j_8;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_27 <= w_sys_tmp665;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h55: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_28 <= r_run_j_8;

									end
								end

							endcase
						end

						7'h59: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_28 <= w_sys_tmp745;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h5b: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_29 <= r_run_j_8;

									end
								end

							endcase
						end

						7'h5f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_copy0_j_29 <= w_sys_tmp820;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp503[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub03_u_datain <= w_sys_tmp506;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub03_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h61: begin
							r_sub03_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_q_addr <= 15'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_q_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_q_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_q_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_q_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_q_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h61: begin
							r_sub03_q_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h5f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp817[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h5f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h61: begin
							r_sub03_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp428[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub02_u_datain <= w_sys_tmp431;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h34: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub02_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h61: begin
							r_sub02_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_q_addr <= 15'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_q_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_q_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_q_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_q_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_q_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h61: begin
							r_sub02_q_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h59: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp742[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h59: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h61: begin
							r_sub02_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								3'h2: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h29: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp349[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h29: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub01_u_datain <= w_sys_tmp352;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h29: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub01_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h61: begin
							r_sub01_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_q_addr <= 15'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_q_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_q_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_q_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_q_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_q_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h61: begin
							r_sub01_q_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp662[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h61: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								3'h3: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h23: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp274[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h23: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub00_u_datain <= w_sys_tmp277;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h23: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub00_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h61: begin
							r_sub00_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_q_addr <= 15'sh0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_q_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_q_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_q_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_q_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_q_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h61: begin
							r_sub00_q_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h48: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp587[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h61: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


endmodule
